magic
tech sky130B
magscale 1 2
timestamp 1667928660
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 137830 700680 137836 700732
rect 137888 700720 137894 700732
rect 157334 700720 157340 700732
rect 137888 700692 157340 700720
rect 137888 700680 137894 700692
rect 157334 700680 157340 700692
rect 157392 700680 157398 700732
rect 155954 700612 155960 700664
rect 156012 700652 156018 700664
rect 202782 700652 202788 700664
rect 156012 700624 202788 700652
rect 156012 700612 156018 700624
rect 202782 700612 202788 700624
rect 202840 700612 202846 700664
rect 157242 700544 157248 700596
rect 157300 700584 157306 700596
rect 218974 700584 218980 700596
rect 157300 700556 218980 700584
rect 157300 700544 157306 700556
rect 218974 700544 218980 700556
rect 219032 700544 219038 700596
rect 89162 700476 89168 700528
rect 89220 700516 89226 700528
rect 160738 700516 160744 700528
rect 89220 700488 160744 700516
rect 89220 700476 89226 700488
rect 160738 700476 160744 700488
rect 160796 700476 160802 700528
rect 24302 700408 24308 700460
rect 24360 700448 24366 700460
rect 162210 700448 162216 700460
rect 24360 700420 162216 700448
rect 24360 700408 24366 700420
rect 162210 700408 162216 700420
rect 162268 700408 162274 700460
rect 8110 700340 8116 700392
rect 8168 700380 8174 700392
rect 162118 700380 162124 700392
rect 8168 700352 162124 700380
rect 8168 700340 8174 700352
rect 162118 700340 162124 700352
rect 162176 700340 162182 700392
rect 148318 700272 148324 700324
rect 148376 700312 148382 700324
rect 543458 700312 543464 700324
rect 148376 700284 543464 700312
rect 148376 700272 148382 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 559650 700312 559656 700324
rect 547846 700284 559656 700312
rect 542998 700204 543004 700256
rect 543056 700244 543062 700256
rect 547846 700244 547874 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 543056 700216 547874 700244
rect 543056 700204 543062 700216
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106918 699700 106924 699712
rect 105504 699672 106924 699700
rect 105504 699660 105510 699672
rect 106918 699660 106924 699672
rect 106976 699660 106982 699712
rect 265618 699660 265624 699712
rect 265676 699700 265682 699712
rect 267642 699700 267648 699712
rect 265676 699672 267648 699700
rect 265676 699660 265682 699672
rect 267642 699660 267648 699672
rect 267700 699660 267706 699712
rect 347038 699660 347044 699712
rect 347096 699700 347102 699712
rect 348786 699700 348792 699712
rect 347096 699672 348792 699700
rect 347096 699660 347102 699672
rect 348786 699660 348792 699672
rect 348844 699660 348850 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 428458 699660 428464 699712
rect 428516 699700 428522 699712
rect 429838 699700 429844 699712
rect 428516 699672 429844 699700
rect 428516 699660 428522 699672
rect 429838 699660 429844 699672
rect 429896 699660 429902 699712
rect 146294 696940 146300 696992
rect 146352 696980 146358 696992
rect 580166 696980 580172 696992
rect 146352 696952 580172 696980
rect 146352 696940 146358 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 161474 683244 161480 683256
rect 3476 683216 161480 683244
rect 3476 683204 3482 683216
rect 161474 683204 161480 683216
rect 161532 683204 161538 683256
rect 146938 683136 146944 683188
rect 146996 683176 147002 683188
rect 580166 683176 580172 683188
rect 146996 683148 580172 683176
rect 146996 683136 147002 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 163498 670732 163504 670744
rect 3568 670704 163504 670732
rect 3568 670692 3574 670704
rect 163498 670692 163504 670704
rect 163556 670692 163562 670744
rect 185578 670692 185584 670744
rect 185636 670732 185642 670744
rect 580166 670732 580172 670744
rect 185636 670704 580172 670732
rect 185636 670692 185642 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 149698 660288 149704 660340
rect 149756 660328 149762 660340
rect 462314 660328 462320 660340
rect 149756 660300 462320 660328
rect 149756 660288 149762 660300
rect 462314 660288 462320 660300
rect 462372 660288 462378 660340
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 163590 656928 163596 656940
rect 3476 656900 163596 656928
rect 3476 656888 3482 656900
rect 163590 656888 163596 656900
rect 163648 656888 163654 656940
rect 182818 643084 182824 643136
rect 182876 643124 182882 643136
rect 580166 643124 580172 643136
rect 182876 643096 580172 643124
rect 182876 643084 182882 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 164234 632108 164240 632120
rect 3476 632080 164240 632108
rect 3476 632068 3482 632080
rect 164234 632068 164240 632080
rect 164292 632068 164298 632120
rect 197998 630640 198004 630692
rect 198056 630680 198062 630692
rect 580166 630680 580172 630692
rect 198056 630652 580172 630680
rect 198056 630640 198062 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 164878 618304 164884 618316
rect 3200 618276 164884 618304
rect 3200 618264 3206 618276
rect 164878 618264 164884 618276
rect 164936 618264 164942 618316
rect 143534 616836 143540 616888
rect 143592 616876 143598 616888
rect 580166 616876 580172 616888
rect 143592 616848 580172 616876
rect 143592 616836 143598 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 164970 605860 164976 605872
rect 3292 605832 164976 605860
rect 3292 605820 3298 605832
rect 164970 605820 164976 605832
rect 165028 605820 165034 605872
rect 142154 590656 142160 590708
rect 142212 590696 142218 590708
rect 579798 590696 579804 590708
rect 142212 590668 579804 590696
rect 142212 590656 142218 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 165614 579680 165620 579692
rect 3384 579652 165620 579680
rect 3384 579640 3390 579652
rect 165614 579640 165620 579652
rect 165672 579640 165678 579692
rect 144178 576852 144184 576904
rect 144236 576892 144242 576904
rect 580166 576892 580172 576904
rect 144236 576864 580172 576892
rect 144236 576852 144242 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 167638 565876 167644 565888
rect 3476 565848 167644 565876
rect 3476 565836 3482 565848
rect 167638 565836 167644 565848
rect 167696 565836 167702 565888
rect 142430 563048 142436 563100
rect 142488 563088 142494 563100
rect 579798 563088 579804 563100
rect 142488 563060 579804 563088
rect 142488 563048 142494 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 165706 553432 165712 553444
rect 3476 553404 165712 553432
rect 3476 553392 3482 553404
rect 165706 553392 165712 553404
rect 165764 553392 165770 553444
rect 188338 536800 188344 536852
rect 188396 536840 188402 536852
rect 580166 536840 580172 536852
rect 188396 536812 580172 536840
rect 188396 536800 188402 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 166994 527184 167000 527196
rect 3476 527156 167000 527184
rect 3476 527144 3482 527156
rect 166994 527144 167000 527156
rect 167052 527144 167058 527196
rect 142798 524424 142804 524476
rect 142856 524464 142862 524476
rect 580166 524464 580172 524476
rect 142856 524436 580172 524464
rect 142856 524424 142862 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 2774 514768 2780 514820
rect 2832 514808 2838 514820
rect 4798 514808 4804 514820
rect 2832 514780 4804 514808
rect 2832 514768 2838 514780
rect 4798 514768 4804 514780
rect 4856 514768 4862 514820
rect 181438 510620 181444 510672
rect 181496 510660 181502 510672
rect 580166 510660 580172 510672
rect 181496 510632 580172 510660
rect 181496 510620 181502 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 167270 501004 167276 501016
rect 3108 500976 167276 501004
rect 3108 500964 3114 500976
rect 167270 500964 167276 500976
rect 167328 500964 167334 501016
rect 139394 484372 139400 484424
rect 139452 484412 139458 484424
rect 580166 484412 580172 484424
rect 139452 484384 580172 484412
rect 139452 484372 139458 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 140038 470568 140044 470620
rect 140096 470608 140102 470620
rect 579982 470608 579988 470620
rect 140096 470580 579988 470608
rect 140096 470568 140102 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 170398 462380 170404 462392
rect 3568 462352 170404 462380
rect 3568 462340 3574 462352
rect 170398 462340 170404 462352
rect 170456 462340 170462 462392
rect 180058 456764 180064 456816
rect 180116 456804 180122 456816
rect 580166 456804 580172 456816
rect 180116 456776 580172 456804
rect 180116 456764 180122 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 170490 448576 170496 448588
rect 3200 448548 170496 448576
rect 3200 448536 3206 448548
rect 170490 448536 170496 448548
rect 170548 448536 170554 448588
rect 157426 447788 157432 447840
rect 157484 447828 157490 447840
rect 169754 447828 169760 447840
rect 157484 447800 169760 447828
rect 157484 447788 157490 447800
rect 169754 447788 169760 447800
rect 169812 447788 169818 447840
rect 138658 430584 138664 430636
rect 138716 430624 138722 430636
rect 580166 430624 580172 430636
rect 138716 430596 580172 430624
rect 138716 430584 138722 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 169754 422328 169760 422340
rect 3568 422300 169760 422328
rect 3568 422288 3574 422300
rect 169754 422288 169760 422300
rect 169812 422288 169818 422340
rect 138750 418140 138756 418192
rect 138808 418180 138814 418192
rect 580166 418180 580172 418192
rect 138808 418152 580172 418180
rect 138808 418140 138814 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 2866 409844 2872 409896
rect 2924 409884 2930 409896
rect 171778 409884 171784 409896
rect 2924 409856 171784 409884
rect 2924 409844 2930 409856
rect 171778 409844 171784 409856
rect 171836 409844 171842 409896
rect 184198 404336 184204 404388
rect 184256 404376 184262 404388
rect 580166 404376 580172 404388
rect 184256 404348 580172 404376
rect 184256 404336 184262 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3510 397468 3516 397520
rect 3568 397508 3574 397520
rect 171870 397508 171876 397520
rect 3568 397480 171876 397508
rect 3568 397468 3574 397480
rect 171870 397468 171876 397480
rect 171928 397468 171934 397520
rect 178678 378156 178684 378208
rect 178736 378196 178742 378208
rect 580166 378196 580172 378208
rect 178736 378168 580172 378196
rect 178736 378156 178742 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 3510 371220 3516 371272
rect 3568 371260 3574 371272
rect 152458 371260 152464 371272
rect 3568 371232 152464 371260
rect 3568 371220 3574 371232
rect 152458 371220 152464 371232
rect 152516 371220 152522 371272
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 113818 357456 113824 357468
rect 3200 357428 113824 357456
rect 3200 357416 3206 357428
rect 113818 357416 113824 357428
rect 113876 357416 113882 357468
rect 135254 351908 135260 351960
rect 135312 351948 135318 351960
rect 580166 351948 580172 351960
rect 135312 351920 580172 351948
rect 135312 351908 135318 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3510 345176 3516 345228
rect 3568 345216 3574 345228
rect 7558 345216 7564 345228
rect 3568 345188 7564 345216
rect 3568 345176 3574 345188
rect 7558 345176 7564 345188
rect 7616 345176 7622 345228
rect 134518 324300 134524 324352
rect 134576 324340 134582 324352
rect 580166 324340 580172 324352
rect 134576 324312 580172 324340
rect 134576 324300 134582 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 173894 318832 173900 318844
rect 3384 318804 173900 318832
rect 3384 318792 3390 318804
rect 173894 318792 173900 318804
rect 173952 318792 173958 318844
rect 135898 311856 135904 311908
rect 135956 311896 135962 311908
rect 579982 311896 579988 311908
rect 135956 311868 579988 311896
rect 135956 311856 135962 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 3510 304988 3516 305040
rect 3568 305028 3574 305040
rect 175918 305028 175924 305040
rect 3568 305000 175924 305028
rect 3568 304988 3574 305000
rect 175918 304988 175924 305000
rect 175976 304988 175982 305040
rect 134610 298120 134616 298172
rect 134668 298160 134674 298172
rect 580166 298160 580172 298172
rect 134668 298132 580172 298160
rect 134668 298120 134674 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 3510 292544 3516 292596
rect 3568 292584 3574 292596
rect 174538 292584 174544 292596
rect 3568 292556 174544 292584
rect 3568 292544 3574 292556
rect 174538 292544 174544 292556
rect 174596 292544 174602 292596
rect 113818 291796 113824 291848
rect 113876 291836 113882 291848
rect 173158 291836 173164 291848
rect 113876 291808 173164 291836
rect 113876 291796 113882 291808
rect 173158 291796 173164 291808
rect 173216 291796 173222 291848
rect 4798 289076 4804 289128
rect 4856 289116 4862 289128
rect 169018 289116 169024 289128
rect 4856 289088 169024 289116
rect 4856 289076 4862 289088
rect 169018 289076 169024 289088
rect 169076 289076 169082 289128
rect 151078 287648 151084 287700
rect 151136 287688 151142 287700
rect 477494 287688 477500 287700
rect 151136 287660 477500 287688
rect 151136 287648 151142 287660
rect 477494 287648 477500 287660
rect 477552 287648 477558 287700
rect 145558 286288 145564 286340
rect 145616 286328 145622 286340
rect 197998 286328 198004 286340
rect 145616 286300 198004 286328
rect 145616 286288 145622 286300
rect 197998 286288 198004 286300
rect 198056 286288 198062 286340
rect 189074 284928 189080 284980
rect 189132 284968 189138 284980
rect 265618 284968 265624 284980
rect 189132 284940 265624 284968
rect 189132 284928 189138 284940
rect 265618 284928 265624 284940
rect 265676 284928 265682 284980
rect 154574 284316 154580 284368
rect 154632 284356 154638 284368
rect 189074 284356 189080 284368
rect 154632 284328 189080 284356
rect 154632 284316 154638 284328
rect 189074 284316 189080 284328
rect 189132 284316 189138 284368
rect 207014 283568 207020 283620
rect 207072 283608 207078 283620
rect 364334 283608 364340 283620
rect 207072 283580 364340 283608
rect 207072 283568 207078 283580
rect 364334 283568 364340 283580
rect 364392 283568 364398 283620
rect 151814 282888 151820 282940
rect 151872 282928 151878 282940
rect 207014 282928 207020 282940
rect 151872 282900 207020 282928
rect 151872 282888 151878 282900
rect 207014 282888 207020 282900
rect 207072 282888 207078 282940
rect 147950 280780 147956 280832
rect 148008 280820 148014 280832
rect 527174 280820 527180 280832
rect 148008 280792 527180 280820
rect 148008 280780 148014 280792
rect 527174 280780 527180 280792
rect 527232 280780 527238 280832
rect 144914 279420 144920 279472
rect 144972 279460 144978 279472
rect 182818 279460 182824 279472
rect 144972 279432 182824 279460
rect 144972 279420 144978 279432
rect 182818 279420 182824 279432
rect 182876 279420 182882 279472
rect 141418 277992 141424 278044
rect 141476 278032 141482 278044
rect 188338 278032 188344 278044
rect 141476 278004 188344 278032
rect 141476 277992 141482 278004
rect 188338 277992 188344 278004
rect 188396 277992 188402 278044
rect 137278 276632 137284 276684
rect 137336 276672 137342 276684
rect 184198 276672 184204 276684
rect 137336 276644 184204 276672
rect 137336 276632 137342 276644
rect 184198 276632 184204 276644
rect 184256 276632 184262 276684
rect 40034 275272 40040 275324
rect 40092 275312 40098 275324
rect 160094 275312 160100 275324
rect 40092 275284 160100 275312
rect 40092 275272 40098 275284
rect 160094 275272 160100 275284
rect 160152 275272 160158 275324
rect 187694 275272 187700 275324
rect 187752 275312 187758 275324
rect 331214 275312 331220 275324
rect 187752 275284 331220 275312
rect 187752 275272 187758 275284
rect 331214 275272 331220 275284
rect 331272 275272 331278 275324
rect 153378 274660 153384 274712
rect 153436 274700 153442 274712
rect 187694 274700 187700 274712
rect 153436 274672 187700 274700
rect 153436 274660 153442 274672
rect 187694 274660 187700 274672
rect 187752 274660 187758 274712
rect 71774 273912 71780 273964
rect 71832 273952 71838 273964
rect 159358 273952 159364 273964
rect 71832 273924 159364 273952
rect 71832 273912 71838 273924
rect 159358 273912 159364 273924
rect 159416 273912 159422 273964
rect 189166 273912 189172 273964
rect 189224 273952 189230 273964
rect 234614 273952 234620 273964
rect 189224 273924 234620 273952
rect 189224 273912 189230 273924
rect 234614 273912 234620 273924
rect 234672 273912 234678 273964
rect 156046 273232 156052 273284
rect 156104 273272 156110 273284
rect 189166 273272 189172 273284
rect 156104 273244 189172 273272
rect 156104 273232 156110 273244
rect 189166 273232 189172 273244
rect 189224 273232 189230 273284
rect 132494 271872 132500 271924
rect 132552 271912 132558 271924
rect 580166 271912 580172 271924
rect 132552 271884 580172 271912
rect 132552 271872 132558 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 137370 271192 137376 271244
rect 137428 271232 137434 271244
rect 178678 271232 178684 271244
rect 137428 271204 178684 271232
rect 137428 271192 137434 271204
rect 178678 271192 178684 271204
rect 178736 271192 178742 271244
rect 149054 271124 149060 271176
rect 149112 271164 149118 271176
rect 494054 271164 494060 271176
rect 149112 271136 494060 271164
rect 149112 271124 149118 271136
rect 494054 271124 494060 271136
rect 494112 271124 494118 271176
rect 7558 269832 7564 269884
rect 7616 269872 7622 269884
rect 172698 269872 172704 269884
rect 7616 269844 172704 269872
rect 7616 269832 7622 269844
rect 172698 269832 172704 269844
rect 172756 269832 172762 269884
rect 147766 269764 147772 269816
rect 147824 269804 147830 269816
rect 542998 269804 543004 269816
rect 147824 269776 543004 269804
rect 147824 269764 147830 269776
rect 542998 269764 543004 269776
rect 543056 269764 543062 269816
rect 3418 268336 3424 268388
rect 3476 268376 3482 268388
rect 120810 268376 120816 268388
rect 3476 268348 120816 268376
rect 3476 268336 3482 268348
rect 120810 268336 120816 268348
rect 120868 268336 120874 268388
rect 146202 268336 146208 268388
rect 146260 268376 146266 268388
rect 185578 268376 185584 268388
rect 146260 268348 185584 268376
rect 146260 268336 146266 268348
rect 185578 268336 185584 268348
rect 185636 268336 185642 268388
rect 120810 267724 120816 267776
rect 120868 267764 120874 267776
rect 168374 267764 168380 267776
rect 120868 267736 168380 267764
rect 120868 267724 120874 267736
rect 168374 267724 168380 267736
rect 168432 267724 168438 267776
rect 207566 266976 207572 267028
rect 207624 267016 207630 267028
rect 299474 267016 299480 267028
rect 207624 266988 299480 267016
rect 207624 266976 207630 266988
rect 299474 266976 299480 266988
rect 299532 266976 299538 267028
rect 154390 266432 154396 266484
rect 154448 266472 154454 266484
rect 207566 266472 207572 266484
rect 154448 266444 207572 266472
rect 154448 266432 154454 266444
rect 207566 266432 207572 266444
rect 207624 266432 207630 266484
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 175918 266404 175924 266416
rect 3108 266376 175924 266404
rect 3108 266364 3114 266376
rect 175918 266364 175924 266376
rect 175976 266364 175982 266416
rect 152458 265752 152464 265804
rect 152516 265792 152522 265804
rect 173342 265792 173348 265804
rect 152516 265764 173348 265792
rect 152516 265752 152522 265764
rect 173342 265752 173348 265764
rect 173400 265752 173406 265804
rect 141326 265684 141332 265736
rect 141384 265724 141390 265736
rect 181438 265724 181444 265736
rect 141384 265696 181444 265724
rect 141384 265684 141390 265696
rect 181438 265684 181444 265696
rect 181496 265684 181502 265736
rect 106918 265616 106924 265668
rect 106976 265656 106982 265668
rect 158714 265656 158720 265668
rect 106976 265628 158720 265656
rect 106976 265616 106982 265628
rect 158714 265616 158720 265628
rect 158772 265616 158778 265668
rect 174538 265616 174544 265668
rect 174596 265656 174602 265668
rect 194870 265656 194876 265668
rect 174596 265628 194876 265656
rect 174596 265616 174602 265628
rect 194870 265616 194876 265628
rect 194928 265616 194934 265668
rect 172790 265548 172796 265600
rect 172848 265588 172854 265600
rect 196250 265588 196256 265600
rect 172848 265560 196256 265588
rect 172848 265548 172854 265560
rect 196250 265548 196256 265560
rect 196308 265548 196314 265600
rect 173434 265480 173440 265532
rect 173492 265520 173498 265532
rect 197354 265520 197360 265532
rect 173492 265492 197360 265520
rect 173492 265480 173498 265492
rect 197354 265480 197360 265492
rect 197412 265480 197418 265532
rect 164878 265412 164884 265464
rect 164936 265452 164942 265464
rect 165430 265452 165436 265464
rect 164936 265424 165436 265452
rect 164936 265412 164942 265424
rect 165430 265412 165436 265424
rect 165488 265412 165494 265464
rect 170214 265412 170220 265464
rect 170272 265452 170278 265464
rect 170490 265452 170496 265464
rect 170272 265424 170496 265452
rect 170272 265412 170278 265424
rect 170490 265412 170496 265424
rect 170548 265452 170554 265464
rect 196158 265452 196164 265464
rect 170548 265424 196164 265452
rect 170548 265412 170554 265424
rect 196158 265412 196164 265424
rect 196216 265412 196222 265464
rect 171778 265344 171784 265396
rect 171836 265384 171842 265396
rect 199010 265384 199016 265396
rect 171836 265356 199016 265384
rect 171836 265344 171842 265356
rect 199010 265344 199016 265356
rect 199068 265344 199074 265396
rect 170398 265276 170404 265328
rect 170456 265316 170462 265328
rect 170674 265316 170680 265328
rect 170456 265288 170680 265316
rect 170456 265276 170462 265288
rect 170674 265276 170680 265288
rect 170732 265316 170738 265328
rect 199194 265316 199200 265328
rect 170732 265288 199200 265316
rect 170732 265276 170738 265288
rect 199194 265276 199200 265288
rect 199252 265276 199258 265328
rect 118326 265208 118332 265260
rect 118384 265248 118390 265260
rect 138750 265248 138756 265260
rect 118384 265220 138756 265248
rect 118384 265208 118390 265220
rect 138750 265208 138756 265220
rect 138808 265208 138814 265260
rect 168742 265208 168748 265260
rect 168800 265248 168806 265260
rect 169018 265248 169024 265260
rect 168800 265220 169024 265248
rect 168800 265208 168806 265220
rect 169018 265208 169024 265220
rect 169076 265248 169082 265260
rect 197998 265248 198004 265260
rect 169076 265220 198004 265248
rect 169076 265208 169082 265220
rect 197998 265208 198004 265220
rect 198056 265208 198062 265260
rect 114186 265140 114192 265192
rect 114244 265180 114250 265192
rect 135898 265180 135904 265192
rect 114244 265152 135904 265180
rect 114244 265140 114250 265152
rect 135898 265140 135904 265152
rect 135956 265140 135962 265192
rect 160830 265140 160836 265192
rect 160888 265180 160894 265192
rect 194778 265180 194784 265192
rect 160888 265152 194784 265180
rect 160888 265140 160894 265152
rect 194778 265140 194784 265152
rect 194836 265140 194842 265192
rect 119982 265072 119988 265124
rect 120040 265112 120046 265124
rect 146938 265112 146944 265124
rect 120040 265084 146944 265112
rect 120040 265072 120046 265084
rect 146938 265072 146944 265084
rect 146996 265072 147002 265124
rect 163498 265072 163504 265124
rect 163556 265112 163562 265124
rect 197906 265112 197912 265124
rect 163556 265084 197912 265112
rect 163556 265072 163562 265084
rect 197906 265072 197912 265084
rect 197964 265072 197970 265124
rect 119890 265004 119896 265056
rect 119948 265044 119954 265056
rect 148502 265044 148508 265056
rect 119948 265016 148508 265044
rect 119948 265004 119954 265016
rect 148502 265004 148508 265016
rect 148560 265004 148566 265056
rect 157242 265004 157248 265056
rect 157300 265044 157306 265056
rect 192202 265044 192208 265056
rect 157300 265016 192208 265044
rect 157300 265004 157306 265016
rect 192202 265004 192208 265016
rect 192260 265004 192266 265056
rect 120718 264936 120724 264988
rect 120776 264976 120782 264988
rect 150710 264976 150716 264988
rect 120776 264948 150716 264976
rect 120776 264936 120782 264948
rect 150710 264936 150716 264948
rect 150768 264976 150774 264988
rect 151078 264976 151084 264988
rect 150768 264948 151084 264976
rect 150768 264936 150774 264948
rect 151078 264936 151084 264948
rect 151136 264936 151142 264988
rect 165430 264936 165436 264988
rect 165488 264976 165494 264988
rect 203242 264976 203248 264988
rect 165488 264948 203248 264976
rect 165488 264936 165494 264948
rect 203242 264936 203248 264948
rect 203300 264936 203306 264988
rect 139486 264188 139492 264240
rect 139544 264228 139550 264240
rect 180058 264228 180064 264240
rect 139544 264200 180064 264228
rect 139544 264188 139550 264200
rect 180058 264188 180064 264200
rect 180116 264188 180122 264240
rect 204806 264188 204812 264240
rect 204864 264228 204870 264240
rect 428458 264228 428464 264240
rect 204864 264200 428464 264228
rect 204864 264188 204870 264200
rect 428458 264188 428464 264200
rect 428516 264188 428522 264240
rect 172606 263848 172612 263900
rect 172664 263888 172670 263900
rect 173342 263888 173348 263900
rect 172664 263860 173348 263888
rect 172664 263848 172670 263860
rect 173342 263848 173348 263860
rect 173400 263888 173406 263900
rect 190638 263888 190644 263900
rect 173400 263860 190644 263888
rect 173400 263848 173406 263860
rect 190638 263848 190644 263860
rect 190696 263848 190702 263900
rect 175734 263780 175740 263832
rect 175792 263820 175798 263832
rect 199286 263820 199292 263832
rect 175792 263792 199292 263820
rect 175792 263780 175798 263792
rect 199286 263780 199292 263792
rect 199344 263780 199350 263832
rect 115474 263712 115480 263764
rect 115532 263752 115538 263764
rect 134426 263752 134432 263764
rect 115532 263724 134432 263752
rect 115532 263712 115538 263724
rect 134426 263712 134432 263724
rect 134484 263752 134490 263764
rect 134610 263752 134616 263764
rect 134484 263724 134616 263752
rect 134484 263712 134490 263724
rect 134610 263712 134616 263724
rect 134668 263712 134674 263764
rect 158714 263712 158720 263764
rect 158772 263752 158778 263764
rect 159266 263752 159272 263764
rect 158772 263724 159272 263752
rect 158772 263712 158778 263724
rect 159266 263712 159272 263724
rect 159324 263752 159330 263764
rect 190730 263752 190736 263764
rect 159324 263724 190736 263752
rect 159324 263712 159330 263724
rect 190730 263712 190736 263724
rect 190788 263712 190794 263764
rect 115566 263644 115572 263696
rect 115624 263684 115630 263696
rect 137278 263684 137284 263696
rect 115624 263656 137284 263684
rect 115624 263644 115630 263656
rect 137278 263644 137284 263656
rect 137336 263684 137342 263696
rect 137554 263684 137560 263696
rect 137336 263656 137560 263684
rect 137336 263644 137342 263656
rect 137554 263644 137560 263656
rect 137612 263644 137618 263696
rect 153194 263644 153200 263696
rect 153252 263684 153258 263696
rect 158806 263684 158812 263696
rect 153252 263656 158812 263684
rect 153252 263644 153258 263656
rect 158806 263644 158812 263656
rect 158864 263684 158870 263696
rect 193766 263684 193772 263696
rect 158864 263656 193772 263684
rect 158864 263644 158870 263656
rect 193766 263644 193772 263656
rect 193824 263644 193830 263696
rect 111518 263576 111524 263628
rect 111576 263616 111582 263628
rect 137370 263616 137376 263628
rect 111576 263588 137376 263616
rect 111576 263576 111582 263588
rect 137370 263576 137376 263588
rect 137428 263576 137434 263628
rect 150894 263576 150900 263628
rect 150952 263616 150958 263628
rect 204806 263616 204812 263628
rect 150952 263588 204812 263616
rect 150952 263576 150958 263588
rect 204806 263576 204812 263588
rect 204864 263576 204870 263628
rect 580258 263548 580264 263560
rect 142126 263520 580264 263548
rect 137462 263440 137468 263492
rect 137520 263480 137526 263492
rect 142126 263480 142154 263520
rect 580258 263508 580264 263520
rect 580316 263508 580322 263560
rect 137520 263452 142154 263480
rect 137520 263440 137526 263452
rect 153194 263440 153200 263492
rect 153252 263480 153258 263492
rect 153378 263480 153384 263492
rect 153252 263452 153384 263480
rect 153252 263440 153258 263452
rect 153378 263440 153384 263452
rect 153436 263440 153442 263492
rect 171686 263236 171692 263288
rect 171744 263276 171750 263288
rect 171870 263276 171876 263288
rect 171744 263248 171876 263276
rect 171744 263236 171750 263248
rect 171870 263236 171876 263248
rect 171928 263236 171934 263288
rect 177758 263168 177764 263220
rect 177816 263208 177822 263220
rect 193950 263208 193956 263220
rect 177816 263180 193956 263208
rect 177816 263168 177822 263180
rect 193950 263168 193956 263180
rect 194008 263168 194014 263220
rect 3418 263100 3424 263152
rect 3476 263140 3482 263152
rect 178034 263140 178040 263152
rect 3476 263112 178040 263140
rect 3476 263100 3482 263112
rect 178034 263100 178040 263112
rect 178092 263100 178098 263152
rect 118142 263032 118148 263084
rect 118200 263072 118206 263084
rect 125962 263072 125968 263084
rect 118200 263044 125968 263072
rect 118200 263032 118206 263044
rect 125962 263032 125968 263044
rect 126020 263032 126026 263084
rect 131114 263032 131120 263084
rect 131172 263072 131178 263084
rect 131758 263072 131764 263084
rect 131172 263044 131764 263072
rect 131172 263032 131178 263044
rect 131758 263032 131764 263044
rect 131816 263072 131822 263084
rect 580534 263072 580540 263084
rect 131816 263044 580540 263072
rect 131816 263032 131822 263044
rect 580534 263032 580540 263044
rect 580592 263032 580598 263084
rect 113818 262964 113824 263016
rect 113876 263004 113882 263016
rect 130102 263004 130108 263016
rect 113876 262976 130108 263004
rect 113876 262964 113882 262976
rect 130102 262964 130108 262976
rect 130160 263004 130166 263016
rect 580350 263004 580356 263016
rect 130160 262976 580356 263004
rect 130160 262964 130166 262976
rect 580350 262964 580356 262976
rect 580408 262964 580414 263016
rect 112346 262896 112352 262948
rect 112404 262936 112410 262948
rect 128354 262936 128360 262948
rect 112404 262908 128360 262936
rect 112404 262896 112410 262908
rect 128354 262896 128360 262908
rect 128412 262896 128418 262948
rect 164970 262896 164976 262948
rect 165028 262936 165034 262948
rect 192386 262936 192392 262948
rect 165028 262908 192392 262936
rect 165028 262896 165034 262908
rect 192386 262896 192392 262908
rect 192444 262896 192450 262948
rect 114094 262828 114100 262880
rect 114152 262868 114158 262880
rect 134518 262868 134524 262880
rect 114152 262840 134524 262868
rect 114152 262828 114158 262840
rect 134518 262828 134524 262840
rect 134576 262868 134582 262880
rect 134794 262868 134800 262880
rect 134576 262840 134800 262868
rect 134576 262828 134582 262840
rect 134794 262828 134800 262840
rect 134852 262828 134858 262880
rect 155862 262828 155868 262880
rect 155920 262868 155926 262880
rect 189350 262868 189356 262880
rect 155920 262840 189356 262868
rect 155920 262828 155926 262840
rect 189350 262828 189356 262840
rect 189408 262868 189414 262880
rect 282914 262868 282920 262880
rect 189408 262840 282920 262868
rect 189408 262828 189414 262840
rect 282914 262828 282920 262840
rect 282972 262828 282978 262880
rect 112622 262760 112628 262812
rect 112680 262800 112686 262812
rect 131114 262800 131120 262812
rect 112680 262772 131120 262800
rect 112680 262760 112686 262772
rect 131114 262760 131120 262772
rect 131172 262760 131178 262812
rect 159358 262760 159364 262812
rect 159416 262800 159422 262812
rect 159910 262800 159916 262812
rect 159416 262772 159916 262800
rect 159416 262760 159422 262772
rect 159910 262760 159916 262772
rect 159968 262800 159974 262812
rect 194042 262800 194048 262812
rect 159968 262772 194048 262800
rect 159968 262760 159974 262772
rect 194042 262760 194048 262772
rect 194100 262760 194106 262812
rect 113910 262692 113916 262744
rect 113968 262732 113974 262744
rect 133046 262732 133052 262744
rect 113968 262704 133052 262732
rect 113968 262692 113974 262704
rect 133046 262692 133052 262704
rect 133104 262692 133110 262744
rect 171686 262692 171692 262744
rect 171744 262732 171750 262744
rect 206002 262732 206008 262744
rect 171744 262704 206008 262732
rect 171744 262692 171750 262704
rect 206002 262692 206008 262704
rect 206060 262692 206066 262744
rect 109770 262624 109776 262676
rect 109828 262664 109834 262676
rect 138658 262664 138664 262676
rect 109828 262636 138664 262664
rect 109828 262624 109834 262636
rect 138658 262624 138664 262636
rect 138716 262624 138722 262676
rect 162210 262624 162216 262676
rect 162268 262664 162274 262676
rect 204622 262664 204628 262676
rect 162268 262636 204628 262664
rect 162268 262624 162274 262636
rect 204622 262624 204628 262636
rect 204680 262624 204686 262676
rect 3602 262556 3608 262608
rect 3660 262596 3666 262608
rect 176746 262596 176752 262608
rect 3660 262568 176752 262596
rect 3660 262556 3666 262568
rect 176746 262556 176752 262568
rect 176804 262556 176810 262608
rect 182910 262556 182916 262608
rect 182968 262596 182974 262608
rect 190454 262596 190460 262608
rect 182968 262568 190460 262596
rect 182968 262556 182974 262568
rect 190454 262556 190460 262568
rect 190512 262556 190518 262608
rect 3510 262488 3516 262540
rect 3568 262528 3574 262540
rect 178402 262528 178408 262540
rect 3568 262500 178408 262528
rect 3568 262488 3574 262500
rect 178402 262488 178408 262500
rect 178460 262488 178466 262540
rect 115382 262420 115388 262472
rect 115440 262460 115446 262472
rect 123202 262460 123208 262472
rect 115440 262432 123208 262460
rect 115440 262420 115446 262432
rect 123202 262420 123208 262432
rect 123260 262420 123266 262472
rect 178034 262420 178040 262472
rect 178092 262460 178098 262472
rect 194962 262460 194968 262472
rect 178092 262432 194968 262460
rect 178092 262420 178098 262432
rect 194962 262420 194968 262432
rect 195020 262420 195026 262472
rect 116854 262352 116860 262404
rect 116912 262392 116918 262404
rect 127618 262392 127624 262404
rect 116912 262364 127624 262392
rect 116912 262352 116918 262364
rect 127618 262352 127624 262364
rect 127676 262352 127682 262404
rect 132034 262352 132040 262404
rect 132092 262392 132098 262404
rect 580442 262392 580448 262404
rect 132092 262364 580448 262392
rect 132092 262352 132098 262364
rect 580442 262352 580448 262364
rect 580500 262352 580506 262404
rect 121362 262284 121368 262336
rect 121420 262324 121426 262336
rect 128722 262324 128728 262336
rect 121420 262296 128728 262324
rect 121420 262284 121426 262296
rect 128722 262284 128728 262296
rect 128780 262284 128786 262336
rect 183462 262284 183468 262336
rect 183520 262324 183526 262336
rect 190822 262324 190828 262336
rect 183520 262296 190828 262324
rect 183520 262284 183526 262296
rect 190822 262284 190828 262296
rect 190880 262284 190886 262336
rect 181254 262216 181260 262268
rect 181312 262256 181318 262268
rect 190546 262256 190552 262268
rect 181312 262228 190552 262256
rect 181312 262216 181318 262228
rect 190546 262216 190552 262228
rect 190604 262216 190610 262268
rect 4798 261400 4804 261452
rect 4856 261440 4862 261452
rect 177758 261440 177764 261452
rect 4856 261412 177764 261440
rect 4856 261400 4862 261412
rect 177758 261400 177764 261412
rect 177816 261400 177822 261452
rect 115290 261332 115296 261384
rect 115348 261372 115354 261384
rect 137462 261372 137468 261384
rect 115348 261344 137468 261372
rect 115348 261332 115354 261344
rect 137462 261332 137468 261344
rect 137520 261332 137526 261384
rect 176746 261332 176752 261384
rect 176804 261372 176810 261384
rect 197814 261372 197820 261384
rect 176804 261344 197820 261372
rect 176804 261332 176810 261344
rect 197814 261332 197820 261344
rect 197872 261332 197878 261384
rect 133046 261264 133052 261316
rect 133104 261304 133110 261316
rect 472618 261304 472624 261316
rect 133104 261276 472624 261304
rect 133104 261264 133110 261276
rect 472618 261264 472624 261276
rect 472676 261264 472682 261316
rect 116486 261196 116492 261248
rect 116544 261236 116550 261248
rect 134334 261236 134340 261248
rect 116544 261208 134340 261236
rect 116544 261196 116550 261208
rect 134334 261196 134340 261208
rect 134392 261196 134398 261248
rect 180150 261196 180156 261248
rect 180208 261236 180214 261248
rect 193674 261236 193680 261248
rect 180208 261208 193680 261236
rect 180208 261196 180214 261208
rect 193674 261196 193680 261208
rect 193732 261196 193738 261248
rect 121270 261128 121276 261180
rect 121328 261168 121334 261180
rect 132034 261168 132040 261180
rect 121328 261140 132040 261168
rect 121328 261128 121334 261140
rect 132034 261128 132040 261140
rect 132092 261128 132098 261180
rect 180518 261128 180524 261180
rect 180576 261168 180582 261180
rect 195054 261168 195060 261180
rect 180576 261140 195060 261168
rect 180576 261128 180582 261140
rect 195054 261128 195060 261140
rect 195112 261128 195118 261180
rect 118050 261060 118056 261112
rect 118108 261100 118114 261112
rect 131114 261100 131120 261112
rect 118108 261072 131120 261100
rect 118108 261060 118114 261072
rect 131114 261060 131120 261072
rect 131172 261060 131178 261112
rect 181990 261060 181996 261112
rect 182048 261100 182054 261112
rect 199102 261100 199108 261112
rect 182048 261072 199108 261100
rect 182048 261060 182054 261072
rect 199102 261060 199108 261072
rect 199160 261060 199166 261112
rect 119522 260992 119528 261044
rect 119580 261032 119586 261044
rect 125594 261032 125600 261044
rect 119580 261004 125600 261032
rect 119580 260992 119586 261004
rect 125594 260992 125600 261004
rect 125652 260992 125658 261044
rect 178402 260992 178408 261044
rect 178460 261032 178466 261044
rect 196434 261032 196440 261044
rect 178460 261004 196440 261032
rect 178460 260992 178466 261004
rect 196434 260992 196440 261004
rect 196492 260992 196498 261044
rect 119614 260924 119620 260976
rect 119672 260964 119678 260976
rect 127066 260964 127072 260976
rect 119672 260936 127072 260964
rect 119672 260924 119678 260936
rect 127066 260924 127072 260936
rect 127124 260924 127130 260976
rect 181806 260924 181812 260976
rect 181864 260964 181870 260976
rect 192110 260964 192116 260976
rect 181864 260936 192116 260964
rect 181864 260924 181870 260936
rect 192110 260924 192116 260936
rect 192168 260924 192174 260976
rect 119246 260856 119252 260908
rect 119304 260896 119310 260908
rect 130378 260896 130384 260908
rect 119304 260868 130384 260896
rect 119304 260856 119310 260868
rect 130378 260856 130384 260868
rect 130436 260856 130442 260908
rect 184750 260856 184756 260908
rect 184808 260896 184814 260908
rect 196342 260896 196348 260908
rect 184808 260868 196348 260896
rect 184808 260856 184814 260868
rect 196342 260856 196348 260868
rect 196400 260856 196406 260908
rect 119430 260788 119436 260840
rect 119488 260828 119494 260840
rect 124306 260828 124312 260840
rect 119488 260800 124312 260828
rect 119488 260788 119494 260800
rect 124306 260788 124312 260800
rect 124364 260788 124370 260840
rect 167270 260788 167276 260840
rect 167328 260828 167334 260840
rect 168190 260828 168196 260840
rect 167328 260800 168196 260828
rect 167328 260788 167334 260800
rect 168190 260788 168196 260800
rect 168248 260788 168254 260840
rect 117866 260720 117872 260772
rect 117924 260760 117930 260772
rect 122834 260760 122840 260772
rect 117924 260732 122840 260760
rect 117924 260720 117930 260732
rect 122834 260720 122840 260732
rect 122892 260720 122898 260772
rect 173894 260380 173900 260432
rect 173952 260420 173958 260432
rect 181898 260420 181904 260432
rect 173952 260392 181904 260420
rect 173952 260380 173958 260392
rect 181898 260380 181904 260392
rect 181956 260380 181962 260432
rect 134334 260312 134340 260364
rect 134392 260352 134398 260364
rect 187786 260352 187792 260364
rect 134392 260324 187792 260352
rect 134392 260312 134398 260324
rect 187786 260312 187792 260324
rect 187844 260312 187850 260364
rect 166626 260244 166632 260296
rect 166684 260284 166690 260296
rect 206094 260284 206100 260296
rect 166684 260256 206100 260284
rect 166684 260244 166690 260256
rect 206094 260244 206100 260256
rect 206152 260244 206158 260296
rect 7558 260176 7564 260228
rect 7616 260216 7622 260228
rect 176194 260216 176200 260228
rect 7616 260188 176200 260216
rect 7616 260176 7622 260188
rect 176194 260176 176200 260188
rect 176252 260176 176258 260228
rect 184106 260176 184112 260228
rect 184164 260216 184170 260228
rect 192478 260216 192484 260228
rect 184164 260188 192484 260216
rect 184164 260176 184170 260188
rect 192478 260176 192484 260188
rect 192536 260176 192542 260228
rect 157334 260108 157340 260160
rect 157392 260148 157398 260160
rect 158300 260148 158306 260160
rect 157392 260120 158306 260148
rect 157392 260108 157398 260120
rect 158300 260108 158306 260120
rect 158358 260108 158364 260160
rect 165706 260108 165712 260160
rect 165764 260148 165770 260160
rect 166580 260148 166586 260160
rect 165764 260120 166586 260148
rect 165764 260108 165770 260120
rect 166580 260108 166586 260120
rect 166638 260108 166644 260160
rect 169754 260108 169760 260160
rect 169812 260148 169818 260160
rect 170996 260148 171002 260160
rect 169812 260120 171002 260148
rect 169812 260108 169818 260120
rect 170996 260108 171002 260120
rect 171054 260148 171060 260160
rect 200574 260148 200580 260160
rect 171054 260120 200580 260148
rect 171054 260108 171060 260120
rect 200574 260108 200580 260120
rect 200632 260108 200638 260160
rect 116394 260040 116400 260092
rect 116452 260080 116458 260092
rect 147950 260080 147956 260092
rect 116452 260052 147956 260080
rect 116452 260040 116458 260052
rect 147950 260040 147956 260052
rect 148008 260040 148014 260092
rect 166994 260040 167000 260092
rect 167052 260080 167058 260092
rect 167684 260080 167690 260092
rect 167052 260052 167690 260080
rect 167052 260040 167058 260052
rect 167684 260040 167690 260052
rect 167742 260080 167748 260092
rect 167742 260052 171134 260080
rect 167742 260040 167748 260052
rect 116670 259972 116676 260024
rect 116728 260012 116734 260024
rect 139394 260012 139400 260024
rect 116728 259984 139400 260012
rect 116728 259972 116734 259984
rect 139394 259972 139400 259984
rect 139452 259972 139458 260024
rect 171106 260012 171134 260052
rect 181898 260040 181904 260092
rect 181956 260080 181962 260092
rect 193858 260080 193864 260092
rect 181956 260052 193864 260080
rect 181956 260040 181962 260052
rect 193858 260040 193864 260052
rect 193916 260040 193922 260092
rect 189258 260012 189264 260024
rect 171106 259984 189264 260012
rect 189258 259972 189264 259984
rect 189316 259972 189322 260024
rect 119338 259904 119344 259956
rect 119396 259944 119402 259956
rect 132494 259944 132500 259956
rect 119396 259916 132500 259944
rect 119396 259904 119402 259916
rect 132494 259904 132500 259916
rect 132552 259944 132558 259956
rect 133138 259944 133144 259956
rect 132552 259916 133144 259944
rect 132552 259904 132558 259916
rect 133138 259904 133144 259916
rect 133196 259904 133202 259956
rect 166350 259904 166356 259956
rect 166408 259944 166414 259956
rect 190914 259944 190920 259956
rect 166408 259916 190920 259944
rect 166408 259904 166414 259916
rect 190914 259904 190920 259916
rect 190972 259904 190978 259956
rect 117958 259836 117964 259888
rect 118016 259876 118022 259888
rect 140866 259876 140872 259888
rect 118016 259848 140872 259876
rect 118016 259836 118022 259848
rect 140866 259836 140872 259848
rect 140924 259836 140930 259888
rect 176102 259836 176108 259888
rect 176160 259876 176166 259888
rect 203334 259876 203340 259888
rect 176160 259848 203340 259876
rect 176160 259836 176166 259848
rect 203334 259836 203340 259848
rect 203392 259836 203398 259888
rect 115198 259768 115204 259820
rect 115256 259808 115262 259820
rect 139670 259808 139676 259820
rect 115256 259780 139676 259808
rect 115256 259768 115262 259780
rect 139670 259768 139676 259780
rect 139728 259768 139734 259820
rect 168098 259768 168104 259820
rect 168156 259808 168162 259820
rect 196618 259808 196624 259820
rect 168156 259780 196624 259808
rect 168156 259768 168162 259780
rect 196618 259768 196624 259780
rect 196676 259768 196682 259820
rect 116578 259700 116584 259752
rect 116636 259740 116642 259752
rect 142430 259740 142436 259752
rect 116636 259712 142436 259740
rect 116636 259700 116642 259712
rect 142430 259700 142436 259712
rect 142488 259700 142494 259752
rect 158070 259700 158076 259752
rect 158128 259740 158134 259752
rect 189718 259740 189724 259752
rect 158128 259712 189724 259740
rect 158128 259700 158134 259712
rect 189718 259700 189724 259712
rect 189776 259700 189782 259752
rect 112530 259632 112536 259684
rect 112588 259672 112594 259684
rect 142154 259672 142160 259684
rect 112588 259644 142160 259672
rect 112588 259632 112594 259644
rect 142154 259632 142160 259644
rect 142212 259672 142218 259684
rect 143074 259672 143080 259684
rect 142212 259644 143080 259672
rect 142212 259632 142218 259644
rect 143074 259632 143080 259644
rect 143132 259632 143138 259684
rect 158622 259632 158628 259684
rect 158680 259672 158686 259684
rect 184106 259672 184112 259684
rect 158680 259644 184112 259672
rect 158680 259632 158686 259644
rect 184106 259632 184112 259644
rect 184164 259632 184170 259684
rect 184566 259632 184572 259684
rect 184624 259672 184630 259684
rect 192570 259672 192576 259684
rect 184624 259644 192576 259672
rect 184624 259632 184630 259644
rect 192570 259632 192576 259644
rect 192628 259632 192634 259684
rect 112806 259564 112812 259616
rect 112864 259604 112870 259616
rect 124858 259604 124864 259616
rect 112864 259576 124864 259604
rect 112864 259564 112870 259576
rect 124858 259564 124864 259576
rect 124916 259564 124922 259616
rect 179414 259564 179420 259616
rect 179472 259604 179478 259616
rect 189626 259604 189632 259616
rect 179472 259576 189632 259604
rect 179472 259564 179478 259576
rect 189626 259564 189632 259576
rect 189684 259564 189690 259616
rect 113726 259496 113732 259548
rect 113784 259536 113790 259548
rect 129274 259536 129280 259548
rect 113784 259508 129280 259536
rect 113784 259496 113790 259508
rect 129274 259496 129280 259508
rect 129332 259496 129338 259548
rect 184014 259496 184020 259548
rect 184072 259536 184078 259548
rect 207658 259536 207664 259548
rect 184072 259508 207664 259536
rect 184072 259496 184078 259508
rect 207658 259496 207664 259508
rect 207716 259496 207722 259548
rect 112898 259428 112904 259480
rect 112956 259468 112962 259480
rect 126514 259468 126520 259480
rect 112956 259440 126520 259468
rect 112956 259428 112962 259440
rect 126514 259428 126520 259440
rect 126572 259428 126578 259480
rect 176378 259428 176384 259480
rect 176436 259468 176442 259480
rect 196526 259468 196532 259480
rect 176436 259440 196532 259468
rect 176436 259428 176442 259440
rect 196526 259428 196532 259440
rect 196584 259428 196590 259480
rect 187786 259360 187792 259412
rect 187844 259400 187850 259412
rect 580166 259400 580172 259412
rect 187844 259372 580172 259400
rect 187844 259360 187850 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 472618 245556 472624 245608
rect 472676 245596 472682 245608
rect 579706 245596 579712 245608
rect 472676 245568 579712 245596
rect 472676 245556 472682 245568
rect 579706 245556 579712 245568
rect 579764 245556 579770 245608
rect 3326 241068 3332 241120
rect 3384 241108 3390 241120
rect 7558 241108 7564 241120
rect 3384 241080 7564 241108
rect 3384 241068 3390 241080
rect 7558 241068 7564 241080
rect 7616 241068 7622 241120
rect 2774 215228 2780 215280
rect 2832 215268 2838 215280
rect 4798 215268 4804 215280
rect 2832 215240 4804 215268
rect 2832 215228 2838 215240
rect 4798 215228 4804 215240
rect 4856 215228 4862 215280
rect 471238 206932 471244 206984
rect 471296 206972 471302 206984
rect 580166 206972 580172 206984
rect 471296 206944 580172 206972
rect 471296 206932 471302 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 187142 200852 187148 200864
rect 131868 200824 144914 200852
rect 131868 200728 131896 200824
rect 132052 200756 137048 200784
rect 132052 200728 132080 200756
rect 123938 200676 123944 200728
rect 123996 200716 124002 200728
rect 123996 200688 129734 200716
rect 123996 200676 124002 200688
rect 120626 200608 120632 200660
rect 120684 200648 120690 200660
rect 129706 200648 129734 200688
rect 131850 200676 131856 200728
rect 131908 200676 131914 200728
rect 132034 200676 132040 200728
rect 132092 200676 132098 200728
rect 137020 200648 137048 200756
rect 144886 200648 144914 200824
rect 183526 200824 187148 200852
rect 162826 200756 177390 200784
rect 120684 200620 122834 200648
rect 129706 200620 135944 200648
rect 137020 200620 142154 200648
rect 144886 200620 150526 200648
rect 120684 200608 120690 200620
rect 108942 200540 108948 200592
rect 109000 200580 109006 200592
rect 122806 200580 122834 200620
rect 132218 200580 132224 200592
rect 109000 200552 115934 200580
rect 122806 200552 132224 200580
rect 109000 200540 109006 200552
rect 115906 200512 115934 200552
rect 132218 200540 132224 200552
rect 132276 200540 132282 200592
rect 123938 200512 123944 200524
rect 115906 200484 123944 200512
rect 123938 200472 123944 200484
rect 123996 200472 124002 200524
rect 128998 200472 129004 200524
rect 129056 200512 129062 200524
rect 132034 200512 132040 200524
rect 129056 200484 132040 200512
rect 129056 200472 129062 200484
rect 132034 200472 132040 200484
rect 132092 200472 132098 200524
rect 135916 200512 135944 200620
rect 142126 200580 142154 200620
rect 142126 200552 150434 200580
rect 135916 200484 140774 200512
rect 107562 200404 107568 200456
rect 107620 200444 107626 200456
rect 120626 200444 120632 200456
rect 107620 200416 120632 200444
rect 107620 200404 107626 200416
rect 120626 200404 120632 200416
rect 120684 200404 120690 200456
rect 118602 200336 118608 200388
rect 118660 200376 118666 200388
rect 131850 200376 131856 200388
rect 118660 200348 131856 200376
rect 118660 200336 118666 200348
rect 131850 200336 131856 200348
rect 131908 200336 131914 200388
rect 140746 200376 140774 200484
rect 140746 200348 142798 200376
rect 118510 200268 118516 200320
rect 118568 200308 118574 200320
rect 118568 200280 140452 200308
rect 118568 200268 118574 200280
rect 117222 200200 117228 200252
rect 117280 200240 117286 200252
rect 117280 200212 134794 200240
rect 117280 200200 117286 200212
rect 129642 200132 129648 200184
rect 129700 200172 129706 200184
rect 129700 200144 134702 200172
rect 129700 200132 129706 200144
rect 119430 200064 119436 200116
rect 119488 200104 119494 200116
rect 125042 200104 125048 200116
rect 119488 200076 125048 200104
rect 119488 200064 119494 200076
rect 125042 200064 125048 200076
rect 125100 200064 125106 200116
rect 133202 200076 133874 200104
rect 126606 199996 126612 200048
rect 126664 200036 126670 200048
rect 133202 200036 133230 200076
rect 126664 200008 133230 200036
rect 126664 199996 126670 200008
rect 130654 199928 130660 199980
rect 130712 199968 130718 199980
rect 133846 199968 133874 200076
rect 130712 199940 133138 199968
rect 133846 199940 134150 199968
rect 130712 199928 130718 199940
rect 133110 199912 133138 199940
rect 134122 199912 134150 199940
rect 134674 199912 134702 200144
rect 134766 200036 134794 200212
rect 135134 200212 136634 200240
rect 135134 200036 135162 200212
rect 136606 200172 136634 200212
rect 140424 200172 140452 200280
rect 136606 200144 138934 200172
rect 140424 200144 140544 200172
rect 134766 200008 135162 200036
rect 135226 200076 138842 200104
rect 129274 199860 129280 199912
rect 129332 199900 129338 199912
rect 132908 199900 132914 199912
rect 129332 199872 132914 199900
rect 129332 199860 129338 199872
rect 132908 199860 132914 199872
rect 132966 199860 132972 199912
rect 133000 199860 133006 199912
rect 133058 199860 133064 199912
rect 133092 199860 133098 199912
rect 133150 199860 133156 199912
rect 133736 199860 133742 199912
rect 133794 199860 133800 199912
rect 133920 199860 133926 199912
rect 133978 199860 133984 199912
rect 134104 199860 134110 199912
rect 134162 199860 134168 199912
rect 134380 199860 134386 199912
rect 134438 199860 134444 199912
rect 134472 199860 134478 199912
rect 134530 199860 134536 199912
rect 134656 199860 134662 199912
rect 134714 199860 134720 199912
rect 134840 199860 134846 199912
rect 134898 199860 134904 199912
rect 127158 199792 127164 199844
rect 127216 199832 127222 199844
rect 132540 199832 132546 199844
rect 127216 199804 132546 199832
rect 127216 199792 127222 199804
rect 132540 199792 132546 199804
rect 132598 199792 132604 199844
rect 126974 199724 126980 199776
rect 127032 199764 127038 199776
rect 133018 199764 133046 199860
rect 133754 199776 133782 199860
rect 127032 199736 133046 199764
rect 127032 199724 127038 199736
rect 133690 199724 133696 199776
rect 133748 199736 133782 199776
rect 133938 199776 133966 199860
rect 134398 199776 134426 199860
rect 133938 199736 133972 199776
rect 133748 199724 133754 199736
rect 133966 199724 133972 199736
rect 134024 199724 134030 199776
rect 134058 199724 134064 199776
rect 134116 199764 134122 199776
rect 134288 199764 134294 199776
rect 134116 199736 134294 199764
rect 134116 199724 134122 199736
rect 134288 199724 134294 199736
rect 134346 199724 134352 199776
rect 134380 199724 134386 199776
rect 134438 199724 134444 199776
rect 134490 199764 134518 199860
rect 134610 199764 134616 199776
rect 134490 199736 134616 199764
rect 134610 199724 134616 199736
rect 134668 199724 134674 199776
rect 134702 199724 134708 199776
rect 134760 199764 134766 199776
rect 134858 199764 134886 199860
rect 134760 199736 134886 199764
rect 134760 199724 134766 199736
rect 132310 199656 132316 199708
rect 132368 199696 132374 199708
rect 135024 199696 135030 199708
rect 132368 199668 135030 199696
rect 132368 199656 132374 199668
rect 135024 199656 135030 199668
rect 135082 199656 135088 199708
rect 104526 199588 104532 199640
rect 104584 199628 104590 199640
rect 135226 199628 135254 200076
rect 135410 199940 135852 199968
rect 135410 199912 135438 199940
rect 135300 199860 135306 199912
rect 135358 199860 135364 199912
rect 135392 199860 135398 199912
rect 135450 199860 135456 199912
rect 135576 199860 135582 199912
rect 135634 199860 135640 199912
rect 135668 199860 135674 199912
rect 135726 199860 135732 199912
rect 104584 199600 135254 199628
rect 135318 199628 135346 199860
rect 135594 199640 135622 199860
rect 135686 199708 135714 199860
rect 135686 199668 135720 199708
rect 135714 199656 135720 199668
rect 135772 199656 135778 199708
rect 135824 199640 135852 199940
rect 135962 199940 136864 199968
rect 135962 199912 135990 199940
rect 135944 199860 135950 199912
rect 136002 199860 136008 199912
rect 136036 199860 136042 199912
rect 136094 199860 136100 199912
rect 136128 199860 136134 199912
rect 136186 199860 136192 199912
rect 136312 199860 136318 199912
rect 136370 199860 136376 199912
rect 136496 199860 136502 199912
rect 136554 199860 136560 199912
rect 136680 199860 136686 199912
rect 136738 199860 136744 199912
rect 136054 199776 136082 199860
rect 135990 199724 135996 199776
rect 136048 199736 136082 199776
rect 136048 199724 136054 199736
rect 136146 199708 136174 199860
rect 136330 199776 136358 199860
rect 136330 199736 136364 199776
rect 136358 199724 136364 199736
rect 136416 199724 136422 199776
rect 136514 199764 136542 199860
rect 136698 199776 136726 199860
rect 136514 199736 136588 199764
rect 136698 199736 136732 199776
rect 136082 199656 136088 199708
rect 136140 199668 136174 199708
rect 136140 199656 136146 199668
rect 136560 199640 136588 199736
rect 136726 199724 136732 199736
rect 136784 199724 136790 199776
rect 135438 199628 135444 199640
rect 135318 199600 135444 199628
rect 104584 199588 104590 199600
rect 135438 199588 135444 199600
rect 135496 199588 135502 199640
rect 135594 199600 135628 199640
rect 135622 199588 135628 199600
rect 135680 199588 135686 199640
rect 135806 199588 135812 199640
rect 135864 199588 135870 199640
rect 136542 199588 136548 199640
rect 136600 199588 136606 199640
rect 136726 199588 136732 199640
rect 136784 199628 136790 199640
rect 136836 199628 136864 199940
rect 138170 199940 138290 199968
rect 137048 199860 137054 199912
rect 137106 199860 137112 199912
rect 137324 199860 137330 199912
rect 137382 199860 137388 199912
rect 137876 199860 137882 199912
rect 137934 199860 137940 199912
rect 137968 199860 137974 199912
rect 138026 199860 138032 199912
rect 138170 199900 138198 199940
rect 138262 199912 138290 199940
rect 138814 199912 138842 200076
rect 138078 199872 138198 199900
rect 137066 199708 137094 199860
rect 137140 199792 137146 199844
rect 137198 199832 137204 199844
rect 137198 199792 137232 199832
rect 137066 199668 137100 199708
rect 137094 199656 137100 199668
rect 137152 199656 137158 199708
rect 136784 199600 136864 199628
rect 136784 199588 136790 199600
rect 136910 199588 136916 199640
rect 136968 199628 136974 199640
rect 137204 199628 137232 199792
rect 137342 199776 137370 199860
rect 137342 199736 137376 199776
rect 137370 199724 137376 199736
rect 137428 199724 137434 199776
rect 137894 199764 137922 199860
rect 137848 199736 137922 199764
rect 137848 199640 137876 199736
rect 137986 199708 138014 199860
rect 137922 199656 137928 199708
rect 137980 199668 138014 199708
rect 137980 199656 137986 199668
rect 138078 199640 138106 199872
rect 138244 199860 138250 199912
rect 138302 199860 138308 199912
rect 138336 199860 138342 199912
rect 138394 199860 138400 199912
rect 138520 199860 138526 199912
rect 138578 199860 138584 199912
rect 138796 199860 138802 199912
rect 138854 199860 138860 199912
rect 138354 199640 138382 199860
rect 138538 199832 138566 199860
rect 136968 199600 137232 199628
rect 136968 199588 136974 199600
rect 137830 199588 137836 199640
rect 137888 199588 137894 199640
rect 138078 199600 138112 199640
rect 138106 199588 138112 199600
rect 138164 199588 138170 199640
rect 138290 199588 138296 199640
rect 138348 199600 138382 199640
rect 138492 199804 138566 199832
rect 138492 199628 138520 199804
rect 138566 199724 138572 199776
rect 138624 199764 138630 199776
rect 138906 199764 138934 200144
rect 139256 199900 139262 199912
rect 139228 199860 139262 199900
rect 139314 199860 139320 199912
rect 139348 199860 139354 199912
rect 139406 199860 139412 199912
rect 139440 199860 139446 199912
rect 139498 199860 139504 199912
rect 139532 199860 139538 199912
rect 139590 199860 139596 199912
rect 139716 199860 139722 199912
rect 139774 199900 139780 199912
rect 139774 199860 139808 199900
rect 139900 199860 139906 199912
rect 139958 199860 139964 199912
rect 139992 199860 139998 199912
rect 140050 199860 140056 199912
rect 140268 199860 140274 199912
rect 140326 199860 140332 199912
rect 139228 199776 139256 199860
rect 139366 199832 139394 199860
rect 139320 199804 139394 199832
rect 138624 199736 138934 199764
rect 138624 199724 138630 199736
rect 139210 199724 139216 199776
rect 139268 199724 139274 199776
rect 139320 199708 139348 199804
rect 139458 199776 139486 199860
rect 139550 199832 139578 199860
rect 139550 199804 139624 199832
rect 139458 199736 139492 199776
rect 139486 199724 139492 199736
rect 139544 199724 139550 199776
rect 139302 199656 139308 199708
rect 139360 199656 139366 199708
rect 139394 199656 139400 199708
rect 139452 199696 139458 199708
rect 139596 199696 139624 199804
rect 139780 199776 139808 199860
rect 139918 199832 139946 199860
rect 139872 199804 139946 199832
rect 139872 199776 139900 199804
rect 140010 199776 140038 199860
rect 139762 199724 139768 199776
rect 139820 199724 139826 199776
rect 139854 199724 139860 199776
rect 139912 199724 139918 199776
rect 139946 199724 139952 199776
rect 140004 199736 140038 199776
rect 140004 199724 140010 199736
rect 139452 199668 139624 199696
rect 139452 199656 139458 199668
rect 138658 199628 138664 199640
rect 138492 199600 138664 199628
rect 138348 199588 138354 199600
rect 138658 199588 138664 199600
rect 138716 199588 138722 199640
rect 138750 199588 138756 199640
rect 138808 199628 138814 199640
rect 140286 199628 140314 199860
rect 140360 199792 140366 199844
rect 140418 199792 140424 199844
rect 138808 199600 140314 199628
rect 140378 199640 140406 199792
rect 140378 199600 140412 199640
rect 138808 199588 138814 199600
rect 140406 199588 140412 199600
rect 140464 199588 140470 199640
rect 140516 199628 140544 200144
rect 140608 199940 141050 199968
rect 140608 199696 140636 199940
rect 141022 199912 141050 199940
rect 142770 199912 142798 200348
rect 144564 200212 149882 200240
rect 142862 199940 143442 199968
rect 140728 199860 140734 199912
rect 140786 199860 140792 199912
rect 140820 199860 140826 199912
rect 140878 199860 140884 199912
rect 141004 199860 141010 199912
rect 141062 199860 141068 199912
rect 141740 199900 141746 199912
rect 141114 199872 141746 199900
rect 140746 199776 140774 199860
rect 140682 199724 140688 199776
rect 140740 199736 140774 199776
rect 140838 199764 140866 199860
rect 140958 199764 140964 199776
rect 140838 199736 140964 199764
rect 140740 199724 140746 199736
rect 140958 199724 140964 199736
rect 141016 199724 141022 199776
rect 140774 199696 140780 199708
rect 140608 199668 140780 199696
rect 140774 199656 140780 199668
rect 140832 199656 140838 199708
rect 140866 199656 140872 199708
rect 140924 199696 140930 199708
rect 141114 199696 141142 199872
rect 141740 199860 141746 199872
rect 141798 199860 141804 199912
rect 141832 199860 141838 199912
rect 141890 199860 141896 199912
rect 142016 199860 142022 199912
rect 142074 199860 142080 199912
rect 142108 199860 142114 199912
rect 142166 199860 142172 199912
rect 142200 199860 142206 199912
rect 142258 199860 142264 199912
rect 142292 199860 142298 199912
rect 142350 199860 142356 199912
rect 142384 199860 142390 199912
rect 142442 199900 142448 199912
rect 142442 199872 142614 199900
rect 142442 199860 142448 199872
rect 141556 199832 141562 199844
rect 141528 199792 141562 199832
rect 141614 199792 141620 199844
rect 141528 199708 141556 199792
rect 140924 199668 141142 199696
rect 140924 199656 140930 199668
rect 141510 199656 141516 199708
rect 141568 199656 141574 199708
rect 141850 199640 141878 199860
rect 142034 199640 142062 199860
rect 141602 199628 141608 199640
rect 140516 199600 141608 199628
rect 141602 199588 141608 199600
rect 141660 199588 141666 199640
rect 141786 199588 141792 199640
rect 141844 199600 141878 199640
rect 141844 199588 141850 199600
rect 141970 199588 141976 199640
rect 142028 199600 142062 199640
rect 142028 199588 142034 199600
rect 97626 199520 97632 199572
rect 97684 199560 97690 199572
rect 142126 199560 142154 199860
rect 142218 199776 142246 199860
rect 142310 199832 142338 199860
rect 142586 199832 142614 199872
rect 142752 199860 142758 199912
rect 142810 199860 142816 199912
rect 142310 199804 142384 199832
rect 142586 199804 142752 199832
rect 142218 199736 142252 199776
rect 142246 199724 142252 199736
rect 142304 199724 142310 199776
rect 142246 199588 142252 199640
rect 142304 199628 142310 199640
rect 142356 199628 142384 199804
rect 142724 199776 142752 199804
rect 142706 199724 142712 199776
rect 142764 199724 142770 199776
rect 142304 199600 142384 199628
rect 142304 199588 142310 199600
rect 97684 199532 142154 199560
rect 97684 199520 97690 199532
rect 142338 199520 142344 199572
rect 142396 199560 142402 199572
rect 142862 199560 142890 199940
rect 143414 199912 143442 199940
rect 143598 199940 143810 199968
rect 143120 199860 143126 199912
rect 143178 199860 143184 199912
rect 143212 199860 143218 199912
rect 143270 199860 143276 199912
rect 143396 199860 143402 199912
rect 143454 199860 143460 199912
rect 143488 199860 143494 199912
rect 143546 199860 143552 199912
rect 143138 199696 143166 199860
rect 142396 199532 142890 199560
rect 143000 199668 143166 199696
rect 143000 199560 143028 199668
rect 143074 199588 143080 199640
rect 143132 199628 143138 199640
rect 143230 199628 143258 199860
rect 143304 199792 143310 199844
rect 143362 199792 143368 199844
rect 143132 199600 143258 199628
rect 143132 199588 143138 199600
rect 143322 199572 143350 199792
rect 143506 199776 143534 199860
rect 143442 199724 143448 199776
rect 143500 199736 143534 199776
rect 143500 199724 143506 199736
rect 143598 199696 143626 199940
rect 143782 199912 143810 199940
rect 143672 199860 143678 199912
rect 143730 199860 143736 199912
rect 143764 199860 143770 199912
rect 143822 199860 143828 199912
rect 143948 199860 143954 199912
rect 144006 199860 144012 199912
rect 144040 199860 144046 199912
rect 144098 199860 144104 199912
rect 144132 199860 144138 199912
rect 144190 199860 144196 199912
rect 144224 199860 144230 199912
rect 144282 199860 144288 199912
rect 144316 199860 144322 199912
rect 144374 199860 144380 199912
rect 143690 199764 143718 199860
rect 143966 199776 143994 199860
rect 143810 199764 143816 199776
rect 143690 199736 143816 199764
rect 143810 199724 143816 199736
rect 143868 199724 143874 199776
rect 143902 199724 143908 199776
rect 143960 199736 143994 199776
rect 143960 199724 143966 199736
rect 144058 199708 144086 199860
rect 143598 199668 143672 199696
rect 143644 199640 143672 199668
rect 143994 199656 144000 199708
rect 144052 199668 144086 199708
rect 144052 199656 144058 199668
rect 143626 199588 143632 199640
rect 143684 199588 143690 199640
rect 143166 199560 143172 199572
rect 143000 199532 143172 199560
rect 142396 199520 142402 199532
rect 143166 199520 143172 199532
rect 143224 199520 143230 199572
rect 143258 199520 143264 199572
rect 143316 199532 143350 199572
rect 143316 199520 143322 199532
rect 97902 199452 97908 199504
rect 97960 199492 97966 199504
rect 144150 199492 144178 199860
rect 144242 199776 144270 199860
rect 144334 199832 144362 199860
rect 144334 199804 144408 199832
rect 144380 199776 144408 199804
rect 144242 199736 144276 199776
rect 144270 199724 144276 199736
rect 144328 199724 144334 199776
rect 144362 199724 144368 199776
rect 144420 199724 144426 199776
rect 144564 199628 144592 200212
rect 145392 199940 146294 199968
rect 144776 199860 144782 199912
rect 144834 199860 144840 199912
rect 144960 199860 144966 199912
rect 145018 199860 145024 199912
rect 144794 199776 144822 199860
rect 144730 199724 144736 199776
rect 144788 199736 144822 199776
rect 144788 199724 144794 199736
rect 97960 199464 144178 199492
rect 144242 199600 144592 199628
rect 97960 199452 97966 199464
rect 116946 199384 116952 199436
rect 117004 199424 117010 199436
rect 123570 199424 123576 199436
rect 117004 199396 123576 199424
rect 117004 199384 117010 199396
rect 123570 199384 123576 199396
rect 123628 199384 123634 199436
rect 127894 199384 127900 199436
rect 127952 199424 127958 199436
rect 127952 199396 143304 199424
rect 127952 199384 127958 199396
rect 115658 199316 115664 199368
rect 115716 199356 115722 199368
rect 143276 199356 143304 199396
rect 143718 199384 143724 199436
rect 143776 199424 143782 199436
rect 144242 199424 144270 199600
rect 144978 199572 145006 199860
rect 145144 199724 145150 199776
rect 145202 199724 145208 199776
rect 145162 199640 145190 199724
rect 145098 199588 145104 199640
rect 145156 199600 145190 199640
rect 145156 199588 145162 199600
rect 144546 199520 144552 199572
rect 144604 199560 144610 199572
rect 144604 199532 144914 199560
rect 144978 199532 145012 199572
rect 144604 199520 144610 199532
rect 144886 199504 144914 199532
rect 145006 199520 145012 199532
rect 145064 199520 145070 199572
rect 145392 199560 145420 199940
rect 146266 199912 146294 199940
rect 147554 199940 147858 199968
rect 145512 199900 145518 199912
rect 145484 199860 145518 199900
rect 145570 199860 145576 199912
rect 145604 199860 145610 199912
rect 145662 199860 145668 199912
rect 145696 199860 145702 199912
rect 145754 199860 145760 199912
rect 145788 199860 145794 199912
rect 145846 199860 145852 199912
rect 146248 199860 146254 199912
rect 146306 199860 146312 199912
rect 146340 199860 146346 199912
rect 146398 199860 146404 199912
rect 146708 199860 146714 199912
rect 146766 199860 146772 199912
rect 146984 199860 146990 199912
rect 147042 199860 147048 199912
rect 145484 199776 145512 199860
rect 145466 199724 145472 199776
rect 145524 199724 145530 199776
rect 145622 199764 145650 199860
rect 145576 199736 145650 199764
rect 145576 199708 145604 199736
rect 145714 199708 145742 199860
rect 145558 199656 145564 199708
rect 145616 199656 145622 199708
rect 145650 199656 145656 199708
rect 145708 199668 145742 199708
rect 145806 199708 145834 199860
rect 146358 199832 146386 199860
rect 146312 199804 146386 199832
rect 145972 199724 145978 199776
rect 146030 199724 146036 199776
rect 146156 199724 146162 199776
rect 146214 199764 146220 199776
rect 146214 199724 146248 199764
rect 145806 199668 145840 199708
rect 145708 199656 145714 199668
rect 145834 199656 145840 199668
rect 145892 199656 145898 199708
rect 145990 199696 146018 199724
rect 145990 199668 146064 199696
rect 146036 199640 146064 199668
rect 146220 199640 146248 199724
rect 145742 199588 145748 199640
rect 145800 199628 145806 199640
rect 145926 199628 145932 199640
rect 145800 199600 145932 199628
rect 145800 199588 145806 199600
rect 145926 199588 145932 199600
rect 145984 199588 145990 199640
rect 146018 199588 146024 199640
rect 146076 199588 146082 199640
rect 146202 199588 146208 199640
rect 146260 199588 146266 199640
rect 145392 199532 145788 199560
rect 145760 199504 145788 199532
rect 144886 199464 144920 199504
rect 144914 199452 144920 199464
rect 144972 199452 144978 199504
rect 145742 199452 145748 199504
rect 145800 199452 145806 199504
rect 146312 199492 146340 199804
rect 146478 199696 146484 199708
rect 146404 199668 146484 199696
rect 146404 199640 146432 199668
rect 146478 199656 146484 199668
rect 146536 199656 146542 199708
rect 146726 199640 146754 199860
rect 146386 199588 146392 199640
rect 146444 199588 146450 199640
rect 146662 199588 146668 199640
rect 146720 199600 146754 199640
rect 147002 199628 147030 199860
rect 147352 199724 147358 199776
rect 147410 199724 147416 199776
rect 147370 199696 147398 199724
rect 147324 199668 147398 199696
rect 147324 199640 147352 199668
rect 147002 199600 147260 199628
rect 146720 199588 146726 199600
rect 146570 199520 146576 199572
rect 146628 199560 146634 199572
rect 147122 199560 147128 199572
rect 146628 199532 147128 199560
rect 146628 199520 146634 199532
rect 147122 199520 147128 199532
rect 147180 199520 147186 199572
rect 146386 199492 146392 199504
rect 146312 199464 146392 199492
rect 146386 199452 146392 199464
rect 146444 199452 146450 199504
rect 143776 199396 144270 199424
rect 143776 199384 143782 199396
rect 146938 199384 146944 199436
rect 146996 199424 147002 199436
rect 147232 199424 147260 199600
rect 147306 199588 147312 199640
rect 147364 199588 147370 199640
rect 147554 199572 147582 199940
rect 147830 199912 147858 199940
rect 148934 199940 149514 199968
rect 147628 199860 147634 199912
rect 147686 199860 147692 199912
rect 147720 199860 147726 199912
rect 147778 199860 147784 199912
rect 147812 199860 147818 199912
rect 147870 199860 147876 199912
rect 147904 199860 147910 199912
rect 147962 199860 147968 199912
rect 148088 199860 148094 199912
rect 148146 199860 148152 199912
rect 148180 199860 148186 199912
rect 148238 199860 148244 199912
rect 148272 199860 148278 199912
rect 148330 199900 148336 199912
rect 148330 199872 148502 199900
rect 148330 199860 148336 199872
rect 147646 199696 147674 199860
rect 147738 199832 147766 199860
rect 147738 199804 147812 199832
rect 147784 199708 147812 199804
rect 147922 199708 147950 199860
rect 148106 199776 148134 199860
rect 148198 199832 148226 199860
rect 148198 199804 148272 199832
rect 148244 199776 148272 199804
rect 148364 199792 148370 199844
rect 148422 199792 148428 199844
rect 148106 199736 148140 199776
rect 148134 199724 148140 199736
rect 148192 199724 148198 199776
rect 148226 199724 148232 199776
rect 148284 199724 148290 199776
rect 147646 199668 147720 199696
rect 147692 199640 147720 199668
rect 147766 199656 147772 199708
rect 147824 199656 147830 199708
rect 147858 199656 147864 199708
rect 147916 199668 147950 199708
rect 147916 199656 147922 199668
rect 147674 199588 147680 199640
rect 147732 199588 147738 199640
rect 147950 199588 147956 199640
rect 148008 199628 148014 199640
rect 148382 199628 148410 199792
rect 148474 199696 148502 199872
rect 148548 199860 148554 199912
rect 148606 199860 148612 199912
rect 148824 199900 148830 199912
rect 148704 199872 148830 199900
rect 148566 199832 148594 199860
rect 148566 199804 148640 199832
rect 148474 199668 148548 199696
rect 148008 199600 148410 199628
rect 148008 199588 148014 199600
rect 147554 199532 147588 199572
rect 147582 199520 147588 199532
rect 147640 199520 147646 199572
rect 148318 199520 148324 199572
rect 148376 199560 148382 199572
rect 148520 199560 148548 199668
rect 148612 199640 148640 199804
rect 148704 199640 148732 199872
rect 148824 199860 148830 199872
rect 148882 199860 148888 199912
rect 148594 199588 148600 199640
rect 148652 199588 148658 199640
rect 148686 199588 148692 199640
rect 148744 199588 148750 199640
rect 148376 199532 148548 199560
rect 148376 199520 148382 199532
rect 148934 199504 148962 199940
rect 149486 199912 149514 199940
rect 149854 199912 149882 200212
rect 150406 199912 150434 200552
rect 150498 199968 150526 200620
rect 162826 200580 162854 200756
rect 177362 200716 177390 200756
rect 180058 200716 180064 200728
rect 176626 200688 177298 200716
rect 177362 200688 180064 200716
rect 176626 200648 176654 200688
rect 156754 200552 158714 200580
rect 150498 199940 150618 199968
rect 149192 199860 149198 199912
rect 149250 199860 149256 199912
rect 149376 199860 149382 199912
rect 149434 199860 149440 199912
rect 149468 199860 149474 199912
rect 149526 199860 149532 199912
rect 149560 199860 149566 199912
rect 149618 199860 149624 199912
rect 149652 199860 149658 199912
rect 149710 199860 149716 199912
rect 149836 199860 149842 199912
rect 149894 199860 149900 199912
rect 150020 199860 150026 199912
rect 150078 199860 150084 199912
rect 150112 199860 150118 199912
rect 150170 199860 150176 199912
rect 150388 199860 150394 199912
rect 150446 199860 150452 199912
rect 150480 199860 150486 199912
rect 150538 199860 150544 199912
rect 149210 199560 149238 199860
rect 149284 199724 149290 199776
rect 149342 199724 149348 199776
rect 148870 199452 148876 199504
rect 148928 199464 148962 199504
rect 149072 199532 149238 199560
rect 149302 199572 149330 199724
rect 149394 199628 149422 199860
rect 149578 199708 149606 199860
rect 149670 199764 149698 199860
rect 149744 199792 149750 199844
rect 149802 199832 149808 199844
rect 149928 199832 149934 199844
rect 149802 199792 149836 199832
rect 149670 199736 149744 199764
rect 149716 199708 149744 199736
rect 149808 199708 149836 199792
rect 149900 199792 149934 199832
rect 149986 199792 149992 199844
rect 149900 199708 149928 199792
rect 149578 199668 149612 199708
rect 149606 199656 149612 199668
rect 149664 199656 149670 199708
rect 149698 199656 149704 199708
rect 149756 199656 149762 199708
rect 149790 199656 149796 199708
rect 149848 199656 149854 199708
rect 149882 199656 149888 199708
rect 149940 199656 149946 199708
rect 149394 199600 149560 199628
rect 149532 199572 149560 199600
rect 149302 199532 149336 199572
rect 148928 199452 148934 199464
rect 146996 199396 147260 199424
rect 149072 199424 149100 199532
rect 149330 199520 149336 199532
rect 149388 199520 149394 199572
rect 149514 199520 149520 199572
rect 149572 199520 149578 199572
rect 150038 199504 150066 199860
rect 149974 199452 149980 199504
rect 150032 199464 150066 199504
rect 150032 199452 150038 199464
rect 149422 199424 149428 199436
rect 149072 199396 149428 199424
rect 146996 199384 147002 199396
rect 149422 199384 149428 199396
rect 149480 199384 149486 199436
rect 150130 199356 150158 199860
rect 150498 199696 150526 199860
rect 150590 199776 150618 199940
rect 150728 199940 150986 199968
rect 150572 199724 150578 199776
rect 150630 199724 150636 199776
rect 150452 199668 150526 199696
rect 150452 199640 150480 199668
rect 150434 199588 150440 199640
rect 150492 199588 150498 199640
rect 150526 199588 150532 199640
rect 150584 199628 150590 199640
rect 150728 199628 150756 199940
rect 150958 199912 150986 199940
rect 154270 199940 155632 199968
rect 154270 199912 154298 199940
rect 150848 199900 150854 199912
rect 150584 199600 150756 199628
rect 150820 199860 150854 199900
rect 150906 199860 150912 199912
rect 150940 199860 150946 199912
rect 150998 199860 151004 199912
rect 151032 199860 151038 199912
rect 151090 199860 151096 199912
rect 151124 199860 151130 199912
rect 151182 199860 151188 199912
rect 151308 199860 151314 199912
rect 151366 199860 151372 199912
rect 151400 199860 151406 199912
rect 151458 199900 151464 199912
rect 151584 199900 151590 199912
rect 151458 199860 151492 199900
rect 150584 199588 150590 199600
rect 150820 199492 150848 199860
rect 151050 199776 151078 199860
rect 150986 199724 150992 199776
rect 151044 199736 151078 199776
rect 151044 199724 151050 199736
rect 151142 199708 151170 199860
rect 151326 199776 151354 199860
rect 151326 199736 151360 199776
rect 151354 199724 151360 199736
rect 151412 199724 151418 199776
rect 151078 199656 151084 199708
rect 151136 199668 151170 199708
rect 151136 199656 151142 199668
rect 150894 199520 150900 199572
rect 150952 199560 150958 199572
rect 151464 199560 151492 199860
rect 151556 199860 151590 199900
rect 151642 199860 151648 199912
rect 151676 199860 151682 199912
rect 151734 199860 151740 199912
rect 151860 199860 151866 199912
rect 151918 199860 151924 199912
rect 152044 199860 152050 199912
rect 152102 199860 152108 199912
rect 152136 199860 152142 199912
rect 152194 199860 152200 199912
rect 152228 199860 152234 199912
rect 152286 199900 152292 199912
rect 152286 199872 152366 199900
rect 152286 199860 152292 199872
rect 151556 199776 151584 199860
rect 151538 199724 151544 199776
rect 151596 199724 151602 199776
rect 151694 199708 151722 199860
rect 151630 199656 151636 199708
rect 151688 199668 151722 199708
rect 151688 199656 151694 199668
rect 150952 199532 151492 199560
rect 151878 199572 151906 199860
rect 152062 199708 152090 199860
rect 152154 199764 152182 199860
rect 152154 199736 152228 199764
rect 152200 199708 152228 199736
rect 152062 199668 152096 199708
rect 152090 199656 152096 199668
rect 152148 199656 152154 199708
rect 152182 199656 152188 199708
rect 152240 199656 152246 199708
rect 151878 199532 151912 199572
rect 150952 199520 150958 199532
rect 151906 199520 151912 199532
rect 151964 199520 151970 199572
rect 152338 199560 152366 199872
rect 152412 199860 152418 199912
rect 152470 199860 152476 199912
rect 152504 199860 152510 199912
rect 152562 199860 152568 199912
rect 152688 199900 152694 199912
rect 152660 199860 152694 199900
rect 152746 199860 152752 199912
rect 152780 199860 152786 199912
rect 152838 199860 152844 199912
rect 152872 199860 152878 199912
rect 152930 199860 152936 199912
rect 153148 199860 153154 199912
rect 153206 199860 153212 199912
rect 153240 199860 153246 199912
rect 153298 199860 153304 199912
rect 153516 199860 153522 199912
rect 153574 199860 153580 199912
rect 154068 199860 154074 199912
rect 154126 199860 154132 199912
rect 154160 199860 154166 199912
rect 154218 199860 154224 199912
rect 154252 199860 154258 199912
rect 154310 199860 154316 199912
rect 154436 199900 154442 199912
rect 154408 199860 154442 199900
rect 154494 199860 154500 199912
rect 154528 199860 154534 199912
rect 154586 199860 154592 199912
rect 154712 199860 154718 199912
rect 154770 199900 154776 199912
rect 154770 199860 154804 199900
rect 154896 199860 154902 199912
rect 154954 199860 154960 199912
rect 154988 199860 154994 199912
rect 155046 199860 155052 199912
rect 155172 199860 155178 199912
rect 155230 199860 155236 199912
rect 155356 199860 155362 199912
rect 155414 199860 155420 199912
rect 152430 199776 152458 199860
rect 152522 199832 152550 199860
rect 152522 199804 152596 199832
rect 152568 199776 152596 199804
rect 152660 199776 152688 199860
rect 152798 199776 152826 199860
rect 152430 199736 152464 199776
rect 152458 199724 152464 199736
rect 152516 199724 152522 199776
rect 152550 199724 152556 199776
rect 152608 199724 152614 199776
rect 152642 199724 152648 199776
rect 152700 199724 152706 199776
rect 152734 199724 152740 199776
rect 152792 199736 152826 199776
rect 152792 199724 152798 199736
rect 152890 199708 152918 199860
rect 152826 199656 152832 199708
rect 152884 199668 152918 199708
rect 153166 199696 153194 199860
rect 153120 199668 153194 199696
rect 152884 199656 152890 199668
rect 153120 199640 153148 199668
rect 153258 199640 153286 199860
rect 153534 199640 153562 199860
rect 154086 199696 154114 199860
rect 154178 199776 154206 199860
rect 154408 199776 154436 199860
rect 154546 199832 154574 199860
rect 154500 199804 154574 199832
rect 154500 199776 154528 199804
rect 154178 199736 154212 199776
rect 154206 199724 154212 199736
rect 154264 199724 154270 199776
rect 154390 199724 154396 199776
rect 154448 199724 154454 199776
rect 154482 199724 154488 199776
rect 154540 199724 154546 199776
rect 154776 199696 154804 199860
rect 154914 199832 154942 199860
rect 154868 199804 154942 199832
rect 154868 199776 154896 199804
rect 155006 199776 155034 199860
rect 155190 199776 155218 199860
rect 154850 199724 154856 199776
rect 154908 199724 154914 199776
rect 154942 199724 154948 199776
rect 155000 199736 155034 199776
rect 155000 199724 155006 199736
rect 155126 199724 155132 199776
rect 155184 199736 155218 199776
rect 155184 199724 155190 199736
rect 155034 199696 155040 199708
rect 154086 199668 154712 199696
rect 154776 199668 155040 199696
rect 154684 199640 154712 199668
rect 155034 199656 155040 199668
rect 155092 199656 155098 199708
rect 155374 199640 155402 199860
rect 153102 199588 153108 199640
rect 153160 199588 153166 199640
rect 153258 199600 153292 199640
rect 153286 199588 153292 199600
rect 153344 199588 153350 199640
rect 153470 199588 153476 199640
rect 153528 199600 153562 199640
rect 153528 199588 153534 199600
rect 154022 199588 154028 199640
rect 154080 199628 154086 199640
rect 154574 199628 154580 199640
rect 154080 199600 154580 199628
rect 154080 199588 154086 199600
rect 154574 199588 154580 199600
rect 154632 199588 154638 199640
rect 154666 199588 154672 199640
rect 154724 199588 154730 199640
rect 155310 199588 155316 199640
rect 155368 199600 155402 199640
rect 155368 199588 155374 199600
rect 153194 199560 153200 199572
rect 152338 199532 153200 199560
rect 153194 199520 153200 199532
rect 153252 199520 153258 199572
rect 153930 199560 153936 199572
rect 153304 199532 153936 199560
rect 153304 199492 153332 199532
rect 153930 199520 153936 199532
rect 153988 199520 153994 199572
rect 155604 199504 155632 199940
rect 156018 199940 156690 199968
rect 156018 199912 156046 199940
rect 155908 199860 155914 199912
rect 155966 199860 155972 199912
rect 156000 199860 156006 199912
rect 156058 199860 156064 199912
rect 156184 199860 156190 199912
rect 156242 199860 156248 199912
rect 156460 199860 156466 199912
rect 156518 199860 156524 199912
rect 155926 199776 155954 199860
rect 155926 199736 155960 199776
rect 155954 199724 155960 199736
rect 156012 199724 156018 199776
rect 150820 199464 151216 199492
rect 150618 199384 150624 199436
rect 150676 199424 150682 199436
rect 151078 199424 151084 199436
rect 150676 199396 151084 199424
rect 150676 199384 150682 199396
rect 151078 199384 151084 199396
rect 151136 199384 151142 199436
rect 115716 199328 143212 199356
rect 143276 199328 150158 199356
rect 151188 199356 151216 199464
rect 151280 199464 153332 199492
rect 151280 199436 151308 199464
rect 153654 199452 153660 199504
rect 153712 199492 153718 199504
rect 154206 199492 154212 199504
rect 153712 199464 154212 199492
rect 153712 199452 153718 199464
rect 154206 199452 154212 199464
rect 154264 199452 154270 199504
rect 155586 199452 155592 199504
rect 155644 199452 155650 199504
rect 156202 199492 156230 199860
rect 156478 199628 156506 199860
rect 156662 199696 156690 199940
rect 156754 199912 156782 200552
rect 158686 200376 158714 200552
rect 160066 200552 162854 200580
rect 162918 200620 176654 200648
rect 177270 200648 177298 200688
rect 180058 200676 180064 200688
rect 180116 200676 180122 200728
rect 180518 200676 180524 200728
rect 180576 200716 180582 200728
rect 183526 200716 183554 200824
rect 187142 200812 187148 200824
rect 187200 200812 187206 200864
rect 180576 200688 183554 200716
rect 180576 200676 180582 200688
rect 180150 200648 180156 200660
rect 177270 200620 180156 200648
rect 160066 200376 160094 200552
rect 162918 200512 162946 200620
rect 180150 200608 180156 200620
rect 180208 200608 180214 200660
rect 182818 200580 182824 200592
rect 158686 200348 160094 200376
rect 161170 200484 162946 200512
rect 164206 200552 176654 200580
rect 158962 200008 160922 200036
rect 157122 199940 157334 199968
rect 156736 199860 156742 199912
rect 156794 199860 156800 199912
rect 156828 199860 156834 199912
rect 156886 199860 156892 199912
rect 156920 199860 156926 199912
rect 156978 199860 156984 199912
rect 157012 199860 157018 199912
rect 157070 199860 157076 199912
rect 156846 199832 156874 199860
rect 156800 199804 156874 199832
rect 156800 199776 156828 199804
rect 156938 199776 156966 199860
rect 156782 199724 156788 199776
rect 156840 199724 156846 199776
rect 156874 199724 156880 199776
rect 156932 199736 156966 199776
rect 156932 199724 156938 199736
rect 156662 199668 156920 199696
rect 156892 199640 156920 199668
rect 157030 199640 157058 199860
rect 156598 199628 156604 199640
rect 156478 199600 156604 199628
rect 156598 199588 156604 199600
rect 156656 199588 156662 199640
rect 156874 199588 156880 199640
rect 156932 199588 156938 199640
rect 156966 199588 156972 199640
rect 157024 199600 157058 199640
rect 157024 199588 157030 199600
rect 157122 199572 157150 199940
rect 157306 199912 157334 199940
rect 157398 199940 157702 199968
rect 157196 199860 157202 199912
rect 157254 199860 157260 199912
rect 157288 199860 157294 199912
rect 157346 199860 157352 199912
rect 157214 199640 157242 199860
rect 157214 199600 157248 199640
rect 157242 199588 157248 199600
rect 157300 199588 157306 199640
rect 157398 199628 157426 199940
rect 157674 199912 157702 199940
rect 157858 199940 158898 199968
rect 157858 199912 157886 199940
rect 157472 199860 157478 199912
rect 157530 199860 157536 199912
rect 157564 199860 157570 199912
rect 157622 199860 157628 199912
rect 157656 199860 157662 199912
rect 157714 199860 157720 199912
rect 157840 199860 157846 199912
rect 157898 199860 157904 199912
rect 157932 199860 157938 199912
rect 157990 199900 157996 199912
rect 157990 199860 158024 199900
rect 158208 199860 158214 199912
rect 158266 199860 158272 199912
rect 158484 199860 158490 199912
rect 158542 199860 158548 199912
rect 158576 199860 158582 199912
rect 158634 199860 158640 199912
rect 157490 199708 157518 199860
rect 157582 199764 157610 199860
rect 157886 199764 157892 199776
rect 157582 199736 157892 199764
rect 157886 199724 157892 199736
rect 157944 199724 157950 199776
rect 157490 199668 157524 199708
rect 157518 199656 157524 199668
rect 157576 199656 157582 199708
rect 157610 199656 157616 199708
rect 157668 199696 157674 199708
rect 157996 199696 158024 199860
rect 158226 199776 158254 199860
rect 158226 199736 158260 199776
rect 158254 199724 158260 199736
rect 158312 199724 158318 199776
rect 157668 199668 158024 199696
rect 157668 199656 157674 199668
rect 158502 199640 158530 199860
rect 158594 199776 158622 199860
rect 158594 199736 158628 199776
rect 158622 199724 158628 199736
rect 158680 199724 158686 199776
rect 157702 199628 157708 199640
rect 157398 199600 157708 199628
rect 157702 199588 157708 199600
rect 157760 199588 157766 199640
rect 158438 199588 158444 199640
rect 158496 199600 158530 199640
rect 158870 199628 158898 199940
rect 158962 199912 158990 200008
rect 159514 199940 160324 199968
rect 159514 199912 159542 199940
rect 158944 199860 158950 199912
rect 159002 199860 159008 199912
rect 159036 199860 159042 199912
rect 159094 199860 159100 199912
rect 159128 199860 159134 199912
rect 159186 199860 159192 199912
rect 159220 199860 159226 199912
rect 159278 199860 159284 199912
rect 159496 199860 159502 199912
rect 159554 199860 159560 199912
rect 159588 199860 159594 199912
rect 159646 199860 159652 199912
rect 159772 199860 159778 199912
rect 159830 199860 159836 199912
rect 159864 199860 159870 199912
rect 159922 199860 159928 199912
rect 160140 199860 160146 199912
rect 160198 199860 160204 199912
rect 159054 199776 159082 199860
rect 158990 199724 158996 199776
rect 159048 199736 159082 199776
rect 159048 199724 159054 199736
rect 159146 199708 159174 199860
rect 159238 199776 159266 199860
rect 159606 199776 159634 199860
rect 159790 199832 159818 199860
rect 159238 199736 159272 199776
rect 159266 199724 159272 199736
rect 159324 199724 159330 199776
rect 159542 199724 159548 199776
rect 159600 199736 159634 199776
rect 159744 199804 159818 199832
rect 159600 199724 159606 199736
rect 159146 199668 159180 199708
rect 159174 199656 159180 199668
rect 159232 199656 159238 199708
rect 159358 199628 159364 199640
rect 158870 199600 159364 199628
rect 158496 199588 158502 199600
rect 159358 199588 159364 199600
rect 159416 199588 159422 199640
rect 159744 199572 159772 199804
rect 159882 199708 159910 199860
rect 159956 199792 159962 199844
rect 160014 199792 160020 199844
rect 159818 199656 159824 199708
rect 159876 199668 159910 199708
rect 159876 199656 159882 199668
rect 159974 199640 160002 199792
rect 159910 199588 159916 199640
rect 159968 199600 160002 199640
rect 159968 199588 159974 199600
rect 157122 199532 157156 199572
rect 157150 199520 157156 199532
rect 157208 199520 157214 199572
rect 159726 199520 159732 199572
rect 159784 199520 159790 199572
rect 160002 199520 160008 199572
rect 160060 199560 160066 199572
rect 160158 199560 160186 199860
rect 160296 199640 160324 199940
rect 160480 199940 160830 199968
rect 160278 199588 160284 199640
rect 160336 199588 160342 199640
rect 160480 199572 160508 199940
rect 160802 199912 160830 199940
rect 160600 199900 160606 199912
rect 160572 199860 160606 199900
rect 160658 199860 160664 199912
rect 160692 199860 160698 199912
rect 160750 199860 160756 199912
rect 160784 199860 160790 199912
rect 160842 199860 160848 199912
rect 160572 199696 160600 199860
rect 160710 199832 160738 199860
rect 160710 199804 160784 199832
rect 160756 199776 160784 199804
rect 160738 199724 160744 199776
rect 160796 199724 160802 199776
rect 160894 199764 160922 200008
rect 161170 199912 161198 200484
rect 161538 199940 162302 199968
rect 160968 199860 160974 199912
rect 161026 199860 161032 199912
rect 161152 199860 161158 199912
rect 161210 199860 161216 199912
rect 161428 199860 161434 199912
rect 161486 199860 161492 199912
rect 160986 199832 161014 199860
rect 161446 199832 161474 199860
rect 160986 199804 161152 199832
rect 161124 199776 161152 199804
rect 161308 199804 161474 199832
rect 161014 199764 161020 199776
rect 160894 199736 161020 199764
rect 161014 199724 161020 199736
rect 161072 199724 161078 199776
rect 161106 199724 161112 199776
rect 161164 199724 161170 199776
rect 160572 199668 160692 199696
rect 160664 199628 160692 199668
rect 161198 199628 161204 199640
rect 160664 199600 161204 199628
rect 161198 199588 161204 199600
rect 161256 199588 161262 199640
rect 160060 199532 160186 199560
rect 160060 199520 160066 199532
rect 160462 199520 160468 199572
rect 160520 199520 160526 199572
rect 160922 199520 160928 199572
rect 160980 199560 160986 199572
rect 161308 199560 161336 199804
rect 161538 199764 161566 199940
rect 162274 199912 162302 199940
rect 162550 199940 163268 199968
rect 162550 199912 162578 199940
rect 161612 199860 161618 199912
rect 161670 199860 161676 199912
rect 161704 199860 161710 199912
rect 161762 199860 161768 199912
rect 162072 199860 162078 199912
rect 162130 199860 162136 199912
rect 162256 199860 162262 199912
rect 162314 199860 162320 199912
rect 162532 199860 162538 199912
rect 162590 199860 162596 199912
rect 162624 199860 162630 199912
rect 162682 199860 162688 199912
rect 162808 199860 162814 199912
rect 162866 199860 162872 199912
rect 162992 199860 162998 199912
rect 163050 199860 163056 199912
rect 163084 199860 163090 199912
rect 163142 199860 163148 199912
rect 161400 199736 161566 199764
rect 161630 199776 161658 199860
rect 161722 199832 161750 199860
rect 161722 199804 161796 199832
rect 161630 199736 161664 199776
rect 161400 199572 161428 199736
rect 161658 199724 161664 199736
rect 161716 199724 161722 199776
rect 161474 199588 161480 199640
rect 161532 199628 161538 199640
rect 161768 199628 161796 199804
rect 161532 199600 161796 199628
rect 161532 199588 161538 199600
rect 160980 199532 161336 199560
rect 160980 199520 160986 199532
rect 161382 199520 161388 199572
rect 161440 199520 161446 199572
rect 161566 199520 161572 199572
rect 161624 199560 161630 199572
rect 162090 199560 162118 199860
rect 162642 199708 162670 199860
rect 162642 199668 162676 199708
rect 162670 199656 162676 199668
rect 162728 199656 162734 199708
rect 162826 199640 162854 199860
rect 163010 199764 163038 199860
rect 162964 199736 163038 199764
rect 162964 199640 162992 199736
rect 163102 199708 163130 199860
rect 163038 199656 163044 199708
rect 163096 199668 163130 199708
rect 163096 199656 163102 199668
rect 162826 199600 162860 199640
rect 162854 199588 162860 199600
rect 162912 199588 162918 199640
rect 162946 199588 162952 199640
rect 163004 199588 163010 199640
rect 161624 199532 162118 199560
rect 163240 199560 163268 199940
rect 163562 199940 163958 199968
rect 163360 199860 163366 199912
rect 163418 199860 163424 199912
rect 163378 199628 163406 199860
rect 163562 199696 163590 199940
rect 163930 199912 163958 199940
rect 164206 199912 164234 200552
rect 176626 200512 176654 200552
rect 176718 200552 182824 200580
rect 176718 200512 176746 200552
rect 182818 200540 182824 200552
rect 182876 200540 182882 200592
rect 164298 200484 172974 200512
rect 176626 200484 176746 200512
rect 163636 199860 163642 199912
rect 163694 199900 163700 199912
rect 163694 199872 163774 199900
rect 163694 199860 163700 199872
rect 163746 199696 163774 199872
rect 163820 199860 163826 199912
rect 163878 199860 163884 199912
rect 163912 199860 163918 199912
rect 163970 199860 163976 199912
rect 164096 199860 164102 199912
rect 164154 199860 164160 199912
rect 164188 199860 164194 199912
rect 164246 199860 164252 199912
rect 163838 199776 163866 199860
rect 163838 199736 163872 199776
rect 163866 199724 163872 199736
rect 163924 199724 163930 199776
rect 163958 199724 163964 199776
rect 164016 199764 164022 199776
rect 164114 199764 164142 199860
rect 164016 199736 164142 199764
rect 164016 199724 164022 199736
rect 164050 199696 164056 199708
rect 163562 199668 163636 199696
rect 163746 199668 164056 199696
rect 163608 199628 163636 199668
rect 164050 199656 164056 199668
rect 164108 199656 164114 199708
rect 163682 199628 163688 199640
rect 163378 199600 163544 199628
rect 163608 199600 163688 199628
rect 163516 199572 163544 199600
rect 163682 199588 163688 199600
rect 163740 199588 163746 199640
rect 163240 199532 163452 199560
rect 161624 199520 161630 199532
rect 160094 199492 160100 199504
rect 156202 199464 160100 199492
rect 160094 199452 160100 199464
rect 160152 199452 160158 199504
rect 163314 199492 163320 199504
rect 160388 199464 163320 199492
rect 151262 199384 151268 199436
rect 151320 199384 151326 199436
rect 151446 199384 151452 199436
rect 151504 199424 151510 199436
rect 160388 199424 160416 199464
rect 163314 199452 163320 199464
rect 163372 199452 163378 199504
rect 163424 199492 163452 199532
rect 163498 199520 163504 199572
rect 163556 199520 163562 199572
rect 163774 199492 163780 199504
rect 163424 199464 163780 199492
rect 163774 199452 163780 199464
rect 163832 199452 163838 199504
rect 151504 199396 160416 199424
rect 151504 199384 151510 199396
rect 161014 199384 161020 199436
rect 161072 199424 161078 199436
rect 164298 199424 164326 200484
rect 172946 200376 172974 200484
rect 172946 200348 177712 200376
rect 177684 200240 177712 200348
rect 177850 200336 177856 200388
rect 177908 200376 177914 200388
rect 202874 200376 202880 200388
rect 177908 200348 202880 200376
rect 177908 200336 177914 200348
rect 202874 200336 202880 200348
rect 202932 200336 202938 200388
rect 181438 200268 181444 200320
rect 181496 200308 181502 200320
rect 191558 200308 191564 200320
rect 181496 200280 191564 200308
rect 181496 200268 181502 200280
rect 191558 200268 191564 200280
rect 191616 200268 191622 200320
rect 193398 200240 193404 200252
rect 177684 200212 193404 200240
rect 193398 200200 193404 200212
rect 193456 200200 193462 200252
rect 216950 200172 216956 200184
rect 168346 200144 178034 200172
rect 164390 199940 165292 199968
rect 164390 199912 164418 199940
rect 164372 199860 164378 199912
rect 164430 199860 164436 199912
rect 164464 199860 164470 199912
rect 164522 199860 164528 199912
rect 164648 199860 164654 199912
rect 164706 199860 164712 199912
rect 164924 199860 164930 199912
rect 164982 199860 164988 199912
rect 165108 199860 165114 199912
rect 165166 199860 165172 199912
rect 164482 199832 164510 199860
rect 164436 199804 164510 199832
rect 164436 199776 164464 199804
rect 164418 199724 164424 199776
rect 164476 199724 164482 199776
rect 164666 199640 164694 199860
rect 164942 199640 164970 199860
rect 164666 199600 164700 199640
rect 164694 199588 164700 199600
rect 164752 199588 164758 199640
rect 164942 199600 164976 199640
rect 164970 199588 164976 199600
rect 165028 199588 165034 199640
rect 164786 199520 164792 199572
rect 164844 199560 164850 199572
rect 165126 199560 165154 199860
rect 164844 199532 165154 199560
rect 165264 199560 165292 199940
rect 165356 199940 165706 199968
rect 165356 199640 165384 199940
rect 165678 199912 165706 199940
rect 166828 199940 167914 199968
rect 165568 199900 165574 199912
rect 165494 199872 165574 199900
rect 165494 199764 165522 199872
rect 165568 199860 165574 199872
rect 165626 199860 165632 199912
rect 165660 199860 165666 199912
rect 165718 199860 165724 199912
rect 165752 199860 165758 199912
rect 165810 199860 165816 199912
rect 166028 199860 166034 199912
rect 166086 199860 166092 199912
rect 166120 199860 166126 199912
rect 166178 199860 166184 199912
rect 166212 199860 166218 199912
rect 166270 199860 166276 199912
rect 166396 199860 166402 199912
rect 166454 199860 166460 199912
rect 166488 199860 166494 199912
rect 166546 199860 166552 199912
rect 166672 199860 166678 199912
rect 166730 199860 166736 199912
rect 165770 199832 165798 199860
rect 165770 199804 165936 199832
rect 165798 199764 165804 199776
rect 165494 199736 165804 199764
rect 165798 199724 165804 199736
rect 165856 199724 165862 199776
rect 165706 199656 165712 199708
rect 165764 199696 165770 199708
rect 165908 199696 165936 199804
rect 165764 199668 165936 199696
rect 165764 199656 165770 199668
rect 165338 199588 165344 199640
rect 165396 199588 165402 199640
rect 165614 199560 165620 199572
rect 165264 199532 165620 199560
rect 164844 199520 164850 199532
rect 165614 199520 165620 199532
rect 165672 199520 165678 199572
rect 166046 199560 166074 199860
rect 166000 199532 166074 199560
rect 161072 199396 164326 199424
rect 161072 199384 161078 199396
rect 164418 199384 164424 199436
rect 164476 199424 164482 199436
rect 164476 199396 165108 199424
rect 164476 199384 164482 199396
rect 151722 199356 151728 199368
rect 151188 199328 151728 199356
rect 115716 199316 115722 199328
rect 114462 199248 114468 199300
rect 114520 199288 114526 199300
rect 142154 199288 142160 199300
rect 114520 199260 142160 199288
rect 114520 199248 114526 199260
rect 142154 199248 142160 199260
rect 142212 199248 142218 199300
rect 143184 199288 143212 199328
rect 151722 199316 151728 199328
rect 151780 199316 151786 199368
rect 153194 199316 153200 199368
rect 153252 199356 153258 199368
rect 153930 199356 153936 199368
rect 153252 199328 153936 199356
rect 153252 199316 153258 199328
rect 153930 199316 153936 199328
rect 153988 199316 153994 199368
rect 154546 199328 165016 199356
rect 146846 199288 146852 199300
rect 143184 199260 146852 199288
rect 146846 199248 146852 199260
rect 146904 199248 146910 199300
rect 115842 199180 115848 199232
rect 115900 199220 115906 199232
rect 148226 199220 148232 199232
rect 115900 199192 148232 199220
rect 115900 199180 115906 199192
rect 148226 199180 148232 199192
rect 148284 199180 148290 199232
rect 151814 199180 151820 199232
rect 151872 199220 151878 199232
rect 154546 199220 154574 199328
rect 159358 199248 159364 199300
rect 159416 199288 159422 199300
rect 164602 199288 164608 199300
rect 159416 199260 164608 199288
rect 159416 199248 159422 199260
rect 164602 199248 164608 199260
rect 164660 199248 164666 199300
rect 151872 199192 154574 199220
rect 151872 199180 151878 199192
rect 156598 199180 156604 199232
rect 156656 199220 156662 199232
rect 164418 199220 164424 199232
rect 156656 199192 164424 199220
rect 156656 199180 156662 199192
rect 164418 199180 164424 199192
rect 164476 199180 164482 199232
rect 164988 199220 165016 199328
rect 165080 199288 165108 199396
rect 165522 199384 165528 199436
rect 165580 199424 165586 199436
rect 166000 199424 166028 199532
rect 166138 199504 166166 199860
rect 166230 199776 166258 199860
rect 166212 199724 166218 199776
rect 166270 199724 166276 199776
rect 166414 199696 166442 199860
rect 166276 199668 166442 199696
rect 166506 199696 166534 199860
rect 166506 199668 166580 199696
rect 166276 199560 166304 199668
rect 166442 199560 166448 199572
rect 166276 199532 166448 199560
rect 166442 199520 166448 199532
rect 166500 199520 166506 199572
rect 166074 199452 166080 199504
rect 166132 199464 166166 199504
rect 166132 199452 166138 199464
rect 166350 199452 166356 199504
rect 166408 199492 166414 199504
rect 166552 199492 166580 199668
rect 166690 199640 166718 199860
rect 166828 199640 166856 199940
rect 167886 199912 167914 199940
rect 167040 199860 167046 199912
rect 167098 199860 167104 199912
rect 167132 199860 167138 199912
rect 167190 199860 167196 199912
rect 167316 199860 167322 199912
rect 167374 199860 167380 199912
rect 167776 199860 167782 199912
rect 167834 199860 167840 199912
rect 167868 199860 167874 199912
rect 167926 199860 167932 199912
rect 168052 199860 168058 199912
rect 168110 199860 168116 199912
rect 167058 199640 167086 199860
rect 166626 199588 166632 199640
rect 166684 199600 166718 199640
rect 166684 199588 166690 199600
rect 166810 199588 166816 199640
rect 166868 199588 166874 199640
rect 166994 199588 167000 199640
rect 167052 199600 167086 199640
rect 167052 199588 167058 199600
rect 167150 199572 167178 199860
rect 167086 199520 167092 199572
rect 167144 199532 167178 199572
rect 167144 199520 167150 199532
rect 167334 199504 167362 199860
rect 167794 199708 167822 199860
rect 168070 199708 168098 199860
rect 167794 199668 167828 199708
rect 167822 199656 167828 199668
rect 167880 199656 167886 199708
rect 168006 199656 168012 199708
rect 168064 199668 168098 199708
rect 168064 199656 168070 199668
rect 167546 199520 167552 199572
rect 167604 199560 167610 199572
rect 168346 199560 168374 200144
rect 178006 200104 178034 200144
rect 182146 200144 216956 200172
rect 181438 200104 181444 200116
rect 171198 200076 176976 200104
rect 178006 200076 181444 200104
rect 169266 199940 169616 199968
rect 169266 199912 169294 199940
rect 168512 199860 168518 199912
rect 168570 199860 168576 199912
rect 168696 199860 168702 199912
rect 168754 199860 168760 199912
rect 168972 199860 168978 199912
rect 169030 199860 169036 199912
rect 169248 199860 169254 199912
rect 169306 199860 169312 199912
rect 169340 199860 169346 199912
rect 169398 199860 169404 199912
rect 168530 199776 168558 199860
rect 168714 199776 168742 199860
rect 168990 199832 169018 199860
rect 168530 199736 168564 199776
rect 168558 199724 168564 199736
rect 168616 199724 168622 199776
rect 168650 199724 168656 199776
rect 168708 199736 168742 199776
rect 168944 199804 169018 199832
rect 168708 199724 168714 199736
rect 167604 199532 168374 199560
rect 167604 199520 167610 199532
rect 166408 199464 166580 199492
rect 166408 199452 166414 199464
rect 167270 199452 167276 199504
rect 167328 199464 167362 199504
rect 167328 199452 167334 199464
rect 168006 199452 168012 199504
rect 168064 199492 168070 199504
rect 168558 199492 168564 199504
rect 168064 199464 168564 199492
rect 168064 199452 168070 199464
rect 168558 199452 168564 199464
rect 168616 199452 168622 199504
rect 168944 199492 168972 199804
rect 169358 199696 169386 199860
rect 169036 199668 169386 199696
rect 169588 199696 169616 199940
rect 169708 199860 169714 199912
rect 169766 199900 169772 199912
rect 169766 199872 169938 199900
rect 169766 199860 169772 199872
rect 169588 199668 169708 199696
rect 169036 199560 169064 199668
rect 169110 199588 169116 199640
rect 169168 199628 169174 199640
rect 169570 199628 169576 199640
rect 169168 199600 169576 199628
rect 169168 199588 169174 199600
rect 169570 199588 169576 199600
rect 169628 199588 169634 199640
rect 169294 199560 169300 199572
rect 169036 199532 169300 199560
rect 169294 199520 169300 199532
rect 169352 199520 169358 199572
rect 169386 199520 169392 199572
rect 169444 199560 169450 199572
rect 169680 199560 169708 199668
rect 169444 199532 169708 199560
rect 169910 199560 169938 199872
rect 169984 199860 169990 199912
rect 170042 199860 170048 199912
rect 170444 199860 170450 199912
rect 170502 199860 170508 199912
rect 170628 199860 170634 199912
rect 170686 199860 170692 199912
rect 170812 199860 170818 199912
rect 170870 199860 170876 199912
rect 170002 199640 170030 199860
rect 170462 199776 170490 199860
rect 170646 199776 170674 199860
rect 170462 199736 170496 199776
rect 170490 199724 170496 199736
rect 170548 199724 170554 199776
rect 170582 199724 170588 199776
rect 170640 199736 170674 199776
rect 170640 199724 170646 199736
rect 170830 199640 170858 199860
rect 171198 199832 171226 200076
rect 176948 200036 176976 200076
rect 181438 200064 181444 200076
rect 181496 200064 181502 200116
rect 178494 200036 178500 200048
rect 174096 200008 176884 200036
rect 176948 200008 178500 200036
rect 174096 199968 174124 200008
rect 176856 199968 176884 200008
rect 178494 199996 178500 200008
rect 178552 199996 178558 200048
rect 171290 199940 171594 199968
rect 171290 199912 171318 199940
rect 171272 199860 171278 199912
rect 171330 199860 171336 199912
rect 171364 199860 171370 199912
rect 171422 199860 171428 199912
rect 171456 199860 171462 199912
rect 171514 199860 171520 199912
rect 171382 199832 171410 199860
rect 171198 199804 171410 199832
rect 171474 199640 171502 199860
rect 170002 199600 170036 199640
rect 170030 199588 170036 199600
rect 170088 199588 170094 199640
rect 170766 199588 170772 199640
rect 170824 199600 170858 199640
rect 170824 199588 170830 199600
rect 171410 199588 171416 199640
rect 171468 199600 171502 199640
rect 171468 199588 171474 199600
rect 171042 199560 171048 199572
rect 169910 199532 171048 199560
rect 169444 199520 169450 199532
rect 171042 199520 171048 199532
rect 171100 199520 171106 199572
rect 171318 199520 171324 199572
rect 171376 199560 171382 199572
rect 171566 199560 171594 199940
rect 172670 199940 174124 199968
rect 174188 199940 174538 199968
rect 176856 199940 176930 199968
rect 171916 199860 171922 199912
rect 171974 199860 171980 199912
rect 172008 199860 172014 199912
rect 172066 199860 172072 199912
rect 172284 199860 172290 199912
rect 172342 199860 172348 199912
rect 172468 199860 172474 199912
rect 172526 199900 172532 199912
rect 172670 199900 172698 199940
rect 172526 199872 172698 199900
rect 172526 199860 172532 199872
rect 172744 199860 172750 199912
rect 172802 199860 172808 199912
rect 172836 199860 172842 199912
rect 172894 199860 172900 199912
rect 173020 199860 173026 199912
rect 173078 199860 173084 199912
rect 173112 199860 173118 199912
rect 173170 199860 173176 199912
rect 173664 199860 173670 199912
rect 173722 199860 173728 199912
rect 173848 199860 173854 199912
rect 173906 199860 173912 199912
rect 174032 199860 174038 199912
rect 174090 199900 174096 199912
rect 174090 199860 174124 199900
rect 171934 199696 171962 199860
rect 171888 199668 171962 199696
rect 172026 199696 172054 199860
rect 172302 199764 172330 199860
rect 172762 199832 172790 199860
rect 172440 199804 172790 199832
rect 172302 199736 172376 199764
rect 172026 199668 172284 199696
rect 171888 199640 171916 199668
rect 172256 199640 172284 199668
rect 172348 199640 172376 199736
rect 171870 199588 171876 199640
rect 171928 199588 171934 199640
rect 172238 199588 172244 199640
rect 172296 199588 172302 199640
rect 172330 199588 172336 199640
rect 172388 199588 172394 199640
rect 171376 199532 171594 199560
rect 171376 199520 171382 199532
rect 172054 199520 172060 199572
rect 172112 199560 172118 199572
rect 172440 199560 172468 199804
rect 172854 199764 172882 199860
rect 173038 199776 173066 199860
rect 172716 199736 172882 199764
rect 172716 199628 172744 199736
rect 172974 199724 172980 199776
rect 173032 199736 173066 199776
rect 173032 199724 173038 199736
rect 172790 199656 172796 199708
rect 172848 199696 172854 199708
rect 173130 199696 173158 199860
rect 173204 199792 173210 199844
rect 173262 199792 173268 199844
rect 173480 199792 173486 199844
rect 173538 199792 173544 199844
rect 173222 199764 173250 199792
rect 173222 199736 173296 199764
rect 172848 199668 173158 199696
rect 172848 199656 172854 199668
rect 172882 199628 172888 199640
rect 172716 199600 172888 199628
rect 172882 199588 172888 199600
rect 172940 199588 172946 199640
rect 173158 199588 173164 199640
rect 173216 199628 173222 199640
rect 173268 199628 173296 199736
rect 173388 199724 173394 199776
rect 173446 199724 173452 199776
rect 173406 199640 173434 199724
rect 173216 199600 173296 199628
rect 173216 199588 173222 199600
rect 173342 199588 173348 199640
rect 173400 199600 173434 199640
rect 173498 199640 173526 199792
rect 173682 199708 173710 199860
rect 173618 199656 173624 199708
rect 173676 199668 173710 199708
rect 173866 199696 173894 199860
rect 174096 199776 174124 199860
rect 174078 199724 174084 199776
rect 174136 199724 174142 199776
rect 173866 199668 173940 199696
rect 173676 199656 173682 199668
rect 173912 199640 173940 199668
rect 173498 199600 173532 199640
rect 173400 199588 173406 199600
rect 173526 199588 173532 199600
rect 173584 199588 173590 199640
rect 173894 199588 173900 199640
rect 173952 199588 173958 199640
rect 172112 199532 172468 199560
rect 172112 199520 172118 199532
rect 173066 199520 173072 199572
rect 173124 199560 173130 199572
rect 173986 199560 173992 199572
rect 173124 199532 173992 199560
rect 173124 199520 173130 199532
rect 173986 199520 173992 199532
rect 174044 199520 174050 199572
rect 174188 199560 174216 199940
rect 174510 199912 174538 199940
rect 174492 199860 174498 199912
rect 174550 199860 174556 199912
rect 174768 199860 174774 199912
rect 174826 199860 174832 199912
rect 175044 199860 175050 199912
rect 175102 199900 175108 199912
rect 175102 199872 175366 199900
rect 175102 199860 175108 199872
rect 174786 199708 174814 199860
rect 174722 199656 174728 199708
rect 174780 199668 174814 199708
rect 174780 199656 174786 199668
rect 175338 199572 175366 199872
rect 175412 199860 175418 199912
rect 175470 199860 175476 199912
rect 175504 199860 175510 199912
rect 175562 199860 175568 199912
rect 175688 199860 175694 199912
rect 175746 199860 175752 199912
rect 175780 199860 175786 199912
rect 175838 199860 175844 199912
rect 175872 199860 175878 199912
rect 175930 199860 175936 199912
rect 176056 199860 176062 199912
rect 176114 199860 176120 199912
rect 176148 199860 176154 199912
rect 176206 199860 176212 199912
rect 176608 199900 176614 199912
rect 176534 199872 176614 199900
rect 175430 199640 175458 199860
rect 175522 199696 175550 199860
rect 175706 199708 175734 199860
rect 175798 199776 175826 199860
rect 175890 199832 175918 199860
rect 175890 199804 175964 199832
rect 175936 199776 175964 199804
rect 176074 199776 176102 199860
rect 175798 199736 175832 199776
rect 175826 199724 175832 199736
rect 175884 199724 175890 199776
rect 175918 199724 175924 199776
rect 175976 199724 175982 199776
rect 176010 199724 176016 199776
rect 176068 199736 176102 199776
rect 176068 199724 176074 199736
rect 176166 199708 176194 199860
rect 176332 199792 176338 199844
rect 176390 199792 176396 199844
rect 176424 199792 176430 199844
rect 176482 199792 176488 199844
rect 176350 199708 176378 199792
rect 175522 199668 175596 199696
rect 175706 199668 175740 199708
rect 175568 199640 175596 199668
rect 175734 199656 175740 199668
rect 175792 199656 175798 199708
rect 176102 199656 176108 199708
rect 176160 199668 176194 199708
rect 176160 199656 176166 199668
rect 176286 199656 176292 199708
rect 176344 199668 176378 199708
rect 176344 199656 176350 199668
rect 176442 199640 176470 199792
rect 175430 199600 175464 199640
rect 175458 199588 175464 199600
rect 175516 199588 175522 199640
rect 175550 199588 175556 199640
rect 175608 199588 175614 199640
rect 176378 199588 176384 199640
rect 176436 199600 176470 199640
rect 176436 199588 176442 199600
rect 174262 199560 174268 199572
rect 174188 199532 174268 199560
rect 174262 199520 174268 199532
rect 174320 199520 174326 199572
rect 174446 199520 174452 199572
rect 174504 199560 174510 199572
rect 175090 199560 175096 199572
rect 174504 199532 175096 199560
rect 174504 199520 174510 199532
rect 175090 199520 175096 199532
rect 175148 199520 175154 199572
rect 175338 199532 175372 199572
rect 175366 199520 175372 199532
rect 175424 199520 175430 199572
rect 176194 199520 176200 199572
rect 176252 199560 176258 199572
rect 176534 199560 176562 199872
rect 176608 199860 176614 199872
rect 176666 199860 176672 199912
rect 176792 199860 176798 199912
rect 176850 199860 176856 199912
rect 176810 199764 176838 199860
rect 176764 199736 176838 199764
rect 176764 199640 176792 199736
rect 176902 199708 176930 199940
rect 177160 199860 177166 199912
rect 177218 199900 177224 199912
rect 181346 199900 181352 199912
rect 177218 199872 181352 199900
rect 177218 199860 177224 199872
rect 181346 199860 181352 199872
rect 181404 199860 181410 199912
rect 177666 199792 177672 199844
rect 177724 199832 177730 199844
rect 182146 199832 182174 200144
rect 216950 200132 216956 200144
rect 217008 200132 217014 200184
rect 177724 199804 182174 199832
rect 177724 199792 177730 199804
rect 179598 199724 179604 199776
rect 179656 199764 179662 199776
rect 215386 199764 215392 199776
rect 179656 199736 215392 199764
rect 179656 199724 179662 199736
rect 215386 199724 215392 199736
rect 215444 199724 215450 199776
rect 176838 199656 176844 199708
rect 176896 199668 176930 199708
rect 176896 199656 176902 199668
rect 177942 199656 177948 199708
rect 178000 199696 178006 199708
rect 215846 199696 215852 199708
rect 178000 199668 215852 199696
rect 178000 199656 178006 199668
rect 215846 199656 215852 199668
rect 215904 199656 215910 199708
rect 176746 199588 176752 199640
rect 176804 199588 176810 199640
rect 217594 199628 217600 199640
rect 177868 199600 217600 199628
rect 176252 199532 176562 199560
rect 176252 199520 176258 199532
rect 169018 199492 169024 199504
rect 168944 199464 169024 199492
rect 169018 199452 169024 199464
rect 169076 199452 169082 199504
rect 169110 199452 169116 199504
rect 169168 199492 169174 199504
rect 177868 199492 177896 199600
rect 217594 199588 217600 199600
rect 217652 199588 217658 199640
rect 217042 199560 217048 199572
rect 169168 199464 177896 199492
rect 178006 199532 217048 199560
rect 169168 199452 169174 199464
rect 165580 199396 166028 199424
rect 165580 199384 165586 199396
rect 168374 199384 168380 199436
rect 168432 199424 168438 199436
rect 178006 199424 178034 199532
rect 217042 199520 217048 199532
rect 217100 199520 217106 199572
rect 182910 199452 182916 199504
rect 182968 199492 182974 199504
rect 190454 199492 190460 199504
rect 182968 199464 190460 199492
rect 182968 199452 182974 199464
rect 190454 199452 190460 199464
rect 190512 199452 190518 199504
rect 168432 199396 178034 199424
rect 168432 199384 168438 199396
rect 180794 199384 180800 199436
rect 180852 199424 180858 199436
rect 190546 199424 190552 199436
rect 180852 199396 190552 199424
rect 180852 199384 180858 199396
rect 190546 199384 190552 199396
rect 190604 199384 190610 199436
rect 165154 199316 165160 199368
rect 165212 199356 165218 199368
rect 165430 199356 165436 199368
rect 165212 199328 165436 199356
rect 165212 199316 165218 199328
rect 165430 199316 165436 199328
rect 165488 199316 165494 199368
rect 166810 199316 166816 199368
rect 166868 199356 166874 199368
rect 192754 199356 192760 199368
rect 166868 199328 192760 199356
rect 166868 199316 166874 199328
rect 192754 199316 192760 199328
rect 192812 199316 192818 199368
rect 190454 199288 190460 199300
rect 165080 199260 190460 199288
rect 190454 199248 190460 199260
rect 190512 199248 190518 199300
rect 165154 199220 165160 199232
rect 164988 199192 165160 199220
rect 165154 199180 165160 199192
rect 165212 199180 165218 199232
rect 165430 199180 165436 199232
rect 165488 199220 165494 199232
rect 219526 199220 219532 199232
rect 165488 199192 219532 199220
rect 165488 199180 165494 199192
rect 219526 199180 219532 199192
rect 219584 199180 219590 199232
rect 112990 199112 112996 199164
rect 113048 199152 113054 199164
rect 145374 199152 145380 199164
rect 113048 199124 145380 199152
rect 113048 199112 113054 199124
rect 145374 199112 145380 199124
rect 145432 199112 145438 199164
rect 156322 199112 156328 199164
rect 156380 199152 156386 199164
rect 215478 199152 215484 199164
rect 156380 199124 215484 199152
rect 156380 199112 156386 199124
rect 215478 199112 215484 199124
rect 215536 199112 215542 199164
rect 114278 199044 114284 199096
rect 114336 199084 114342 199096
rect 146110 199084 146116 199096
rect 114336 199056 146116 199084
rect 114336 199044 114342 199056
rect 146110 199044 146116 199056
rect 146168 199044 146174 199096
rect 154758 199044 154764 199096
rect 154816 199084 154822 199096
rect 215938 199084 215944 199096
rect 154816 199056 215944 199084
rect 154816 199044 154822 199056
rect 215938 199044 215944 199056
rect 215996 199044 216002 199096
rect 113082 198976 113088 199028
rect 113140 199016 113146 199028
rect 146754 199016 146760 199028
rect 113140 198988 146760 199016
rect 113140 198976 113146 198988
rect 146754 198976 146760 198988
rect 146812 198976 146818 199028
rect 154482 198976 154488 199028
rect 154540 199016 154546 199028
rect 215294 199016 215300 199028
rect 154540 198988 215300 199016
rect 154540 198976 154546 198988
rect 215294 198976 215300 198988
rect 215352 198976 215358 199028
rect 115750 198908 115756 198960
rect 115808 198948 115814 198960
rect 149606 198948 149612 198960
rect 115808 198920 149612 198948
rect 115808 198908 115814 198920
rect 149606 198908 149612 198920
rect 149664 198908 149670 198960
rect 165614 198908 165620 198960
rect 165672 198948 165678 198960
rect 177390 198948 177396 198960
rect 165672 198920 177396 198948
rect 165672 198908 165678 198920
rect 177390 198908 177396 198920
rect 177448 198908 177454 198960
rect 117130 198840 117136 198892
rect 117188 198880 117194 198892
rect 117188 198852 123524 198880
rect 117188 198840 117194 198852
rect 118418 198772 118424 198824
rect 118476 198812 118482 198824
rect 123496 198812 123524 198852
rect 123570 198840 123576 198892
rect 123628 198880 123634 198892
rect 147306 198880 147312 198892
rect 123628 198852 147312 198880
rect 123628 198840 123634 198852
rect 147306 198840 147312 198852
rect 147364 198840 147370 198892
rect 165798 198840 165804 198892
rect 165856 198880 165862 198892
rect 183002 198880 183008 198892
rect 165856 198852 183008 198880
rect 165856 198840 165862 198852
rect 183002 198840 183008 198852
rect 183060 198840 183066 198892
rect 146018 198812 146024 198824
rect 118476 198784 118694 198812
rect 123496 198784 146024 198812
rect 118476 198772 118482 198784
rect 118666 198744 118694 198784
rect 146018 198772 146024 198784
rect 146076 198772 146082 198824
rect 157150 198772 157156 198824
rect 157208 198812 157214 198824
rect 157334 198812 157340 198824
rect 157208 198784 157340 198812
rect 157208 198772 157214 198784
rect 157334 198772 157340 198784
rect 157392 198772 157398 198824
rect 162302 198772 162308 198824
rect 162360 198812 162366 198824
rect 180334 198812 180340 198824
rect 162360 198784 180340 198812
rect 162360 198772 162366 198784
rect 180334 198772 180340 198784
rect 180392 198772 180398 198824
rect 145742 198744 145748 198756
rect 118666 198716 145748 198744
rect 145742 198704 145748 198716
rect 145800 198704 145806 198756
rect 155034 198704 155040 198756
rect 155092 198744 155098 198756
rect 181530 198744 181536 198756
rect 155092 198716 181536 198744
rect 155092 198704 155098 198716
rect 181530 198704 181536 198716
rect 181588 198704 181594 198756
rect 142154 198636 142160 198688
rect 142212 198676 142218 198688
rect 153838 198676 153844 198688
rect 142212 198648 153844 198676
rect 142212 198636 142218 198648
rect 153838 198636 153844 198648
rect 153896 198636 153902 198688
rect 155678 198636 155684 198688
rect 155736 198676 155742 198688
rect 177022 198676 177028 198688
rect 155736 198648 177028 198676
rect 155736 198636 155742 198648
rect 177022 198636 177028 198648
rect 177080 198636 177086 198688
rect 177114 198636 177120 198688
rect 177172 198676 177178 198688
rect 181622 198676 181628 198688
rect 177172 198648 181628 198676
rect 177172 198636 177178 198648
rect 181622 198636 181628 198648
rect 181680 198636 181686 198688
rect 132126 198568 132132 198620
rect 132184 198608 132190 198620
rect 135990 198608 135996 198620
rect 132184 198580 135996 198608
rect 132184 198568 132190 198580
rect 135990 198568 135996 198580
rect 136048 198568 136054 198620
rect 136818 198568 136824 198620
rect 136876 198608 136882 198620
rect 138658 198608 138664 198620
rect 136876 198580 138664 198608
rect 136876 198568 136882 198580
rect 138658 198568 138664 198580
rect 138716 198568 138722 198620
rect 143626 198568 143632 198620
rect 143684 198608 143690 198620
rect 150802 198608 150808 198620
rect 143684 198580 150808 198608
rect 143684 198568 143690 198580
rect 150802 198568 150808 198580
rect 150860 198568 150866 198620
rect 165154 198568 165160 198620
rect 165212 198608 165218 198620
rect 168374 198608 168380 198620
rect 165212 198580 168380 198608
rect 165212 198568 165218 198580
rect 168374 198568 168380 198580
rect 168432 198568 168438 198620
rect 169726 198580 173158 198608
rect 121178 198500 121184 198552
rect 121236 198540 121242 198552
rect 144638 198540 144644 198552
rect 121236 198512 144644 198540
rect 121236 198500 121242 198512
rect 144638 198500 144644 198512
rect 144696 198500 144702 198552
rect 154850 198500 154856 198552
rect 154908 198540 154914 198552
rect 169726 198540 169754 198580
rect 154908 198512 169754 198540
rect 173130 198540 173158 198580
rect 173986 198568 173992 198620
rect 174044 198608 174050 198620
rect 200114 198608 200120 198620
rect 174044 198580 200120 198608
rect 174044 198568 174050 198580
rect 200114 198568 200120 198580
rect 200172 198568 200178 198620
rect 186958 198540 186964 198552
rect 173130 198512 186964 198540
rect 154908 198500 154914 198512
rect 186958 198500 186964 198512
rect 187016 198500 187022 198552
rect 123570 198432 123576 198484
rect 123628 198472 123634 198484
rect 139394 198472 139400 198484
rect 123628 198444 139400 198472
rect 123628 198432 123634 198444
rect 139394 198432 139400 198444
rect 139452 198432 139458 198484
rect 170030 198432 170036 198484
rect 170088 198472 170094 198484
rect 181438 198472 181444 198484
rect 170088 198444 181444 198472
rect 170088 198432 170094 198444
rect 181438 198432 181444 198444
rect 181496 198432 181502 198484
rect 181622 198432 181628 198484
rect 181680 198472 181686 198484
rect 211430 198472 211436 198484
rect 181680 198444 211436 198472
rect 181680 198432 181686 198444
rect 211430 198432 211436 198444
rect 211488 198432 211494 198484
rect 121086 198364 121092 198416
rect 121144 198404 121150 198416
rect 144362 198404 144368 198416
rect 121144 198376 144368 198404
rect 121144 198364 121150 198376
rect 144362 198364 144368 198376
rect 144420 198364 144426 198416
rect 169386 198364 169392 198416
rect 169444 198404 169450 198416
rect 171042 198404 171048 198416
rect 169444 198376 171048 198404
rect 169444 198364 169450 198376
rect 171042 198364 171048 198376
rect 171100 198364 171106 198416
rect 173250 198364 173256 198416
rect 173308 198404 173314 198416
rect 212810 198404 212816 198416
rect 173308 198376 212816 198404
rect 173308 198364 173314 198376
rect 212810 198364 212816 198376
rect 212868 198364 212874 198416
rect 118694 198296 118700 198348
rect 118752 198336 118758 198348
rect 143350 198336 143356 198348
rect 118752 198308 143356 198336
rect 118752 198296 118758 198308
rect 143350 198296 143356 198308
rect 143408 198296 143414 198348
rect 151078 198296 151084 198348
rect 151136 198336 151142 198348
rect 154942 198336 154948 198348
rect 151136 198308 154948 198336
rect 151136 198296 151142 198308
rect 154942 198296 154948 198308
rect 155000 198296 155006 198348
rect 211246 198336 211252 198348
rect 174924 198308 211252 198336
rect 119798 198228 119804 198280
rect 119856 198268 119862 198280
rect 138566 198268 138572 198280
rect 119856 198240 138572 198268
rect 119856 198228 119862 198240
rect 138566 198228 138572 198240
rect 138624 198228 138630 198280
rect 170214 198228 170220 198280
rect 170272 198268 170278 198280
rect 174924 198268 174952 198308
rect 211246 198296 211252 198308
rect 211304 198296 211310 198348
rect 170272 198240 174952 198268
rect 170272 198228 170278 198240
rect 177022 198228 177028 198280
rect 177080 198268 177086 198280
rect 180242 198268 180248 198280
rect 177080 198240 180248 198268
rect 177080 198228 177086 198240
rect 180242 198228 180248 198240
rect 180300 198228 180306 198280
rect 181438 198228 181444 198280
rect 181496 198268 181502 198280
rect 211522 198268 211528 198280
rect 181496 198240 211528 198268
rect 181496 198228 181502 198240
rect 211522 198228 211528 198240
rect 211580 198228 211586 198280
rect 105722 198160 105728 198212
rect 105780 198200 105786 198212
rect 132126 198200 132132 198212
rect 105780 198172 132132 198200
rect 105780 198160 105786 198172
rect 132126 198160 132132 198172
rect 132184 198160 132190 198212
rect 176194 198160 176200 198212
rect 176252 198200 176258 198212
rect 178402 198200 178408 198212
rect 176252 198172 178408 198200
rect 176252 198160 176258 198172
rect 178402 198160 178408 198172
rect 178460 198160 178466 198212
rect 178494 198160 178500 198212
rect 178552 198200 178558 198212
rect 212902 198200 212908 198212
rect 178552 198172 212908 198200
rect 178552 198160 178558 198172
rect 212902 198160 212908 198172
rect 212960 198160 212966 198212
rect 110322 198092 110328 198144
rect 110380 198132 110386 198144
rect 142338 198132 142344 198144
rect 110380 198104 142344 198132
rect 110380 198092 110386 198104
rect 142338 198092 142344 198104
rect 142396 198092 142402 198144
rect 158714 198092 158720 198144
rect 158772 198132 158778 198144
rect 158772 198104 167178 198132
rect 158772 198092 158778 198104
rect 105630 198024 105636 198076
rect 105688 198064 105694 198076
rect 136910 198064 136916 198076
rect 105688 198036 136916 198064
rect 105688 198024 105694 198036
rect 136910 198024 136916 198036
rect 136968 198024 136974 198076
rect 143350 198024 143356 198076
rect 143408 198064 143414 198076
rect 145006 198064 145012 198076
rect 143408 198036 145012 198064
rect 143408 198024 143414 198036
rect 145006 198024 145012 198036
rect 145064 198024 145070 198076
rect 108390 197956 108396 198008
rect 108448 197996 108454 198008
rect 142246 197996 142252 198008
rect 108448 197968 142252 197996
rect 108448 197956 108454 197968
rect 142246 197956 142252 197968
rect 142304 197956 142310 198008
rect 167150 197996 167178 198104
rect 167822 198092 167828 198144
rect 167880 198132 167886 198144
rect 170490 198132 170496 198144
rect 167880 198104 170496 198132
rect 167880 198092 167886 198104
rect 170490 198092 170496 198104
rect 170548 198092 170554 198144
rect 171870 198092 171876 198144
rect 171928 198132 171934 198144
rect 214282 198132 214288 198144
rect 171928 198104 214288 198132
rect 171928 198092 171934 198104
rect 214282 198092 214288 198104
rect 214340 198092 214346 198144
rect 174998 198024 175004 198076
rect 175056 198064 175062 198076
rect 214466 198064 214472 198076
rect 175056 198036 214472 198064
rect 175056 198024 175062 198036
rect 214466 198024 214472 198036
rect 214524 198024 214530 198076
rect 167730 197996 167736 198008
rect 167150 197968 167736 197996
rect 167730 197956 167736 197968
rect 167788 197956 167794 198008
rect 168834 197956 168840 198008
rect 168892 197996 168898 198008
rect 176194 197996 176200 198008
rect 168892 197968 176200 197996
rect 168892 197956 168898 197968
rect 176194 197956 176200 197968
rect 176252 197956 176258 198008
rect 214650 197996 214656 198008
rect 179386 197968 214656 197996
rect 120534 197888 120540 197940
rect 120592 197928 120598 197940
rect 120592 197900 135254 197928
rect 120592 197888 120598 197900
rect 135226 197860 135254 197900
rect 167656 197900 174216 197928
rect 143994 197860 144000 197872
rect 135226 197832 144000 197860
rect 143994 197820 144000 197832
rect 144052 197820 144058 197872
rect 158806 197820 158812 197872
rect 158864 197860 158870 197872
rect 167656 197860 167684 197900
rect 158864 197832 167684 197860
rect 158864 197820 158870 197832
rect 170766 197820 170772 197872
rect 170824 197860 170830 197872
rect 174188 197860 174216 197900
rect 178678 197860 178684 197872
rect 170824 197832 174124 197860
rect 174188 197832 178684 197860
rect 170824 197820 170830 197832
rect 138566 197752 138572 197804
rect 138624 197792 138630 197804
rect 144178 197792 144184 197804
rect 138624 197764 144184 197792
rect 138624 197752 138630 197764
rect 144178 197752 144184 197764
rect 144236 197752 144242 197804
rect 162578 197752 162584 197804
rect 162636 197792 162642 197804
rect 171042 197792 171048 197804
rect 162636 197764 171048 197792
rect 162636 197752 162642 197764
rect 171042 197752 171048 197764
rect 171100 197752 171106 197804
rect 174096 197792 174124 197832
rect 178678 197820 178684 197832
rect 178736 197820 178742 197872
rect 179386 197792 179414 197968
rect 214650 197956 214656 197968
rect 214708 197956 214714 198008
rect 174096 197764 179414 197792
rect 176746 197684 176752 197736
rect 176804 197724 176810 197736
rect 179414 197724 179420 197736
rect 176804 197696 179420 197724
rect 176804 197684 176810 197696
rect 179414 197684 179420 197696
rect 179472 197684 179478 197736
rect 166442 197616 166448 197668
rect 166500 197656 166506 197668
rect 178770 197656 178776 197668
rect 166500 197628 178776 197656
rect 166500 197616 166506 197628
rect 178770 197616 178776 197628
rect 178828 197616 178834 197668
rect 166074 197548 166080 197600
rect 166132 197588 166138 197600
rect 170030 197588 170036 197600
rect 166132 197560 170036 197588
rect 166132 197548 166138 197560
rect 170030 197548 170036 197560
rect 170088 197548 170094 197600
rect 135990 197480 135996 197532
rect 136048 197520 136054 197532
rect 141878 197520 141884 197532
rect 136048 197492 141884 197520
rect 136048 197480 136054 197492
rect 141878 197480 141884 197492
rect 141936 197480 141942 197532
rect 163866 197480 163872 197532
rect 163924 197520 163930 197532
rect 172054 197520 172060 197532
rect 163924 197492 172060 197520
rect 163924 197480 163930 197492
rect 172054 197480 172060 197492
rect 172112 197480 172118 197532
rect 173802 197480 173808 197532
rect 173860 197520 173866 197532
rect 179874 197520 179880 197532
rect 173860 197492 179880 197520
rect 173860 197480 173866 197492
rect 179874 197480 179880 197492
rect 179932 197480 179938 197532
rect 133046 197412 133052 197464
rect 133104 197452 133110 197464
rect 137922 197452 137928 197464
rect 133104 197424 137928 197452
rect 133104 197412 133110 197424
rect 137922 197412 137928 197424
rect 137980 197412 137986 197464
rect 170490 197412 170496 197464
rect 170548 197452 170554 197464
rect 174630 197452 174636 197464
rect 170548 197424 174636 197452
rect 170548 197412 170554 197424
rect 174630 197412 174636 197424
rect 174688 197412 174694 197464
rect 134886 197344 134892 197396
rect 134944 197384 134950 197396
rect 138198 197384 138204 197396
rect 134944 197356 138204 197384
rect 134944 197344 134950 197356
rect 138198 197344 138204 197356
rect 138256 197344 138262 197396
rect 163590 197344 163596 197396
rect 163648 197384 163654 197396
rect 173802 197384 173808 197396
rect 163648 197356 173808 197384
rect 163648 197344 163654 197356
rect 173802 197344 173808 197356
rect 173860 197344 173866 197396
rect 176654 197344 176660 197396
rect 176712 197384 176718 197396
rect 176930 197384 176936 197396
rect 176712 197356 176936 197384
rect 176712 197344 176718 197356
rect 176930 197344 176936 197356
rect 176988 197344 176994 197396
rect 121270 197276 121276 197328
rect 121328 197316 121334 197328
rect 124858 197316 124864 197328
rect 121328 197288 124864 197316
rect 121328 197276 121334 197288
rect 124858 197276 124864 197288
rect 124916 197276 124922 197328
rect 127710 197276 127716 197328
rect 127768 197316 127774 197328
rect 151170 197316 151176 197328
rect 127768 197288 151176 197316
rect 127768 197276 127774 197288
rect 151170 197276 151176 197288
rect 151228 197276 151234 197328
rect 168282 197276 168288 197328
rect 168340 197316 168346 197328
rect 185486 197316 185492 197328
rect 168340 197288 185492 197316
rect 168340 197276 168346 197288
rect 185486 197276 185492 197288
rect 185544 197276 185550 197328
rect 121362 197208 121368 197260
rect 121420 197248 121426 197260
rect 127986 197248 127992 197260
rect 121420 197220 127992 197248
rect 121420 197208 121426 197220
rect 127986 197208 127992 197220
rect 128044 197208 128050 197260
rect 128078 197208 128084 197260
rect 128136 197248 128142 197260
rect 141878 197248 141884 197260
rect 128136 197220 141884 197248
rect 128136 197208 128142 197220
rect 141878 197208 141884 197220
rect 141936 197208 141942 197260
rect 142062 197208 142068 197260
rect 142120 197248 142126 197260
rect 144914 197248 144920 197260
rect 142120 197220 144920 197248
rect 142120 197208 142126 197220
rect 144914 197208 144920 197220
rect 144972 197208 144978 197260
rect 163038 197208 163044 197260
rect 163096 197248 163102 197260
rect 197722 197248 197728 197260
rect 163096 197220 197728 197248
rect 163096 197208 163102 197220
rect 197722 197208 197728 197220
rect 197780 197208 197786 197260
rect 119246 197140 119252 197192
rect 119304 197180 119310 197192
rect 124950 197180 124956 197192
rect 119304 197152 124956 197180
rect 119304 197140 119310 197152
rect 124950 197140 124956 197152
rect 125008 197140 125014 197192
rect 126330 197140 126336 197192
rect 126388 197180 126394 197192
rect 151262 197180 151268 197192
rect 126388 197152 151268 197180
rect 126388 197140 126394 197152
rect 151262 197140 151268 197152
rect 151320 197140 151326 197192
rect 155310 197140 155316 197192
rect 155368 197180 155374 197192
rect 163866 197180 163872 197192
rect 155368 197152 163872 197180
rect 155368 197140 155374 197152
rect 163866 197140 163872 197152
rect 163924 197140 163930 197192
rect 168742 197140 168748 197192
rect 168800 197180 168806 197192
rect 198826 197180 198832 197192
rect 168800 197152 198832 197180
rect 168800 197140 168806 197152
rect 198826 197140 198832 197152
rect 198884 197140 198890 197192
rect 120994 197072 121000 197124
rect 121052 197112 121058 197124
rect 128078 197112 128084 197124
rect 121052 197084 128084 197112
rect 121052 197072 121058 197084
rect 128078 197072 128084 197084
rect 128136 197072 128142 197124
rect 128170 197072 128176 197124
rect 128228 197112 128234 197124
rect 149146 197112 149152 197124
rect 128228 197084 149152 197112
rect 128228 197072 128234 197084
rect 149146 197072 149152 197084
rect 149204 197072 149210 197124
rect 150434 197072 150440 197124
rect 150492 197112 150498 197124
rect 151170 197112 151176 197124
rect 150492 197084 151176 197112
rect 150492 197072 150498 197084
rect 151170 197072 151176 197084
rect 151228 197072 151234 197124
rect 154850 197072 154856 197124
rect 154908 197112 154914 197124
rect 156414 197112 156420 197124
rect 154908 197084 156420 197112
rect 154908 197072 154914 197084
rect 156414 197072 156420 197084
rect 156472 197072 156478 197124
rect 158070 197072 158076 197124
rect 158128 197112 158134 197124
rect 192018 197112 192024 197124
rect 158128 197084 192024 197112
rect 158128 197072 158134 197084
rect 192018 197072 192024 197084
rect 192076 197072 192082 197124
rect 107378 197004 107384 197056
rect 107436 197044 107442 197056
rect 137646 197044 137652 197056
rect 107436 197016 137652 197044
rect 107436 197004 107442 197016
rect 137646 197004 137652 197016
rect 137704 197004 137710 197056
rect 141878 197004 141884 197056
rect 141936 197044 141942 197056
rect 145742 197044 145748 197056
rect 141936 197016 145748 197044
rect 141936 197004 141942 197016
rect 145742 197004 145748 197016
rect 145800 197004 145806 197056
rect 161474 197004 161480 197056
rect 161532 197044 161538 197056
rect 167822 197044 167828 197056
rect 161532 197016 167828 197044
rect 161532 197004 161538 197016
rect 167822 197004 167828 197016
rect 167880 197004 167886 197056
rect 168650 197004 168656 197056
rect 168708 197044 168714 197056
rect 203150 197044 203156 197056
rect 168708 197016 203156 197044
rect 168708 197004 168714 197016
rect 203150 197004 203156 197016
rect 203208 197004 203214 197056
rect 111702 196936 111708 196988
rect 111760 196976 111766 196988
rect 132954 196976 132960 196988
rect 111760 196948 132960 196976
rect 111760 196936 111766 196948
rect 132954 196936 132960 196948
rect 133012 196936 133018 196988
rect 160278 196936 160284 196988
rect 160336 196976 160342 196988
rect 193306 196976 193312 196988
rect 160336 196948 193312 196976
rect 160336 196936 160342 196948
rect 193306 196936 193312 196948
rect 193364 196936 193370 196988
rect 123478 196868 123484 196920
rect 123536 196908 123542 196920
rect 148410 196908 148416 196920
rect 123536 196880 148416 196908
rect 123536 196868 123542 196880
rect 148410 196868 148416 196880
rect 148468 196868 148474 196920
rect 159266 196868 159272 196920
rect 159324 196908 159330 196920
rect 193490 196908 193496 196920
rect 159324 196880 193496 196908
rect 159324 196868 159330 196880
rect 193490 196868 193496 196880
rect 193548 196868 193554 196920
rect 114002 196800 114008 196852
rect 114060 196840 114066 196852
rect 145650 196840 145656 196852
rect 114060 196812 145656 196840
rect 114060 196800 114066 196812
rect 145650 196800 145656 196812
rect 145708 196800 145714 196852
rect 150526 196800 150532 196852
rect 150584 196840 150590 196852
rect 150802 196840 150808 196852
rect 150584 196812 150808 196840
rect 150584 196800 150590 196812
rect 150802 196800 150808 196812
rect 150860 196800 150866 196852
rect 153194 196800 153200 196852
rect 153252 196840 153258 196852
rect 153654 196840 153660 196852
rect 153252 196812 153660 196840
rect 153252 196800 153258 196812
rect 153654 196800 153660 196812
rect 153712 196800 153718 196852
rect 163498 196800 163504 196852
rect 163556 196840 163562 196852
rect 197630 196840 197636 196852
rect 163556 196812 197636 196840
rect 163556 196800 163562 196812
rect 197630 196800 197636 196812
rect 197688 196800 197694 196852
rect 111610 196732 111616 196784
rect 111668 196772 111674 196784
rect 133138 196772 133144 196784
rect 111668 196744 133144 196772
rect 111668 196732 111674 196744
rect 133138 196732 133144 196744
rect 133196 196732 133202 196784
rect 135438 196732 135444 196784
rect 135496 196772 135502 196784
rect 135806 196772 135812 196784
rect 135496 196744 135812 196772
rect 135496 196732 135502 196744
rect 135806 196732 135812 196744
rect 135864 196732 135870 196784
rect 139394 196732 139400 196784
rect 139452 196772 139458 196784
rect 139762 196772 139768 196784
rect 139452 196744 139768 196772
rect 139452 196732 139458 196744
rect 139762 196732 139768 196744
rect 139820 196732 139826 196784
rect 149330 196732 149336 196784
rect 149388 196772 149394 196784
rect 149882 196772 149888 196784
rect 149388 196744 149888 196772
rect 149388 196732 149394 196744
rect 149882 196732 149888 196744
rect 149940 196732 149946 196784
rect 150342 196732 150348 196784
rect 150400 196772 150406 196784
rect 154022 196772 154028 196784
rect 150400 196744 154028 196772
rect 150400 196732 150406 196744
rect 154022 196732 154028 196744
rect 154080 196732 154086 196784
rect 161106 196732 161112 196784
rect 161164 196772 161170 196784
rect 161658 196772 161664 196784
rect 161164 196744 161664 196772
rect 161164 196732 161170 196744
rect 161658 196732 161664 196744
rect 161716 196732 161722 196784
rect 161842 196732 161848 196784
rect 161900 196772 161906 196784
rect 162394 196772 162400 196784
rect 161900 196744 162400 196772
rect 161900 196732 161906 196744
rect 162394 196732 162400 196744
rect 162452 196732 162458 196784
rect 164050 196732 164056 196784
rect 164108 196772 164114 196784
rect 197538 196772 197544 196784
rect 164108 196744 197544 196772
rect 164108 196732 164114 196744
rect 197538 196732 197544 196744
rect 197596 196732 197602 196784
rect 107286 196664 107292 196716
rect 107344 196704 107350 196716
rect 139854 196704 139860 196716
rect 107344 196676 139860 196704
rect 107344 196664 107350 196676
rect 139854 196664 139860 196676
rect 139912 196664 139918 196716
rect 140866 196664 140872 196716
rect 140924 196704 140930 196716
rect 141786 196704 141792 196716
rect 140924 196676 141792 196704
rect 140924 196664 140930 196676
rect 141786 196664 141792 196676
rect 141844 196664 141850 196716
rect 146294 196664 146300 196716
rect 146352 196704 146358 196716
rect 146846 196704 146852 196716
rect 146352 196676 146852 196704
rect 146352 196664 146358 196676
rect 146846 196664 146852 196676
rect 146904 196664 146910 196716
rect 147030 196664 147036 196716
rect 147088 196704 147094 196716
rect 149698 196704 149704 196716
rect 147088 196676 149704 196704
rect 147088 196664 147094 196676
rect 149698 196664 149704 196676
rect 149756 196664 149762 196716
rect 153378 196664 153384 196716
rect 153436 196704 153442 196716
rect 153436 196676 154620 196704
rect 153436 196664 153442 196676
rect 104710 196596 104716 196648
rect 104768 196636 104774 196648
rect 136818 196636 136824 196648
rect 104768 196608 136824 196636
rect 104768 196596 104774 196608
rect 136818 196596 136824 196608
rect 136876 196596 136882 196648
rect 137370 196596 137376 196648
rect 137428 196636 137434 196648
rect 137830 196636 137836 196648
rect 137428 196608 137836 196636
rect 137428 196596 137434 196608
rect 137830 196596 137836 196608
rect 137888 196596 137894 196648
rect 140958 196596 140964 196648
rect 141016 196636 141022 196648
rect 142154 196636 142160 196648
rect 141016 196608 142160 196636
rect 141016 196596 141022 196608
rect 142154 196596 142160 196608
rect 142212 196596 142218 196648
rect 147490 196596 147496 196648
rect 147548 196636 147554 196648
rect 153654 196636 153660 196648
rect 147548 196608 153660 196636
rect 147548 196596 147554 196608
rect 153654 196596 153660 196608
rect 153712 196596 153718 196648
rect 154592 196636 154620 196676
rect 157702 196664 157708 196716
rect 157760 196704 157766 196716
rect 158530 196704 158536 196716
rect 157760 196676 158536 196704
rect 157760 196664 157766 196676
rect 158530 196664 158536 196676
rect 158588 196664 158594 196716
rect 161474 196664 161480 196716
rect 161532 196704 161538 196716
rect 162946 196704 162952 196716
rect 161532 196676 162952 196704
rect 161532 196664 161538 196676
rect 162946 196664 162952 196676
rect 163004 196664 163010 196716
rect 165706 196664 165712 196716
rect 165764 196704 165770 196716
rect 166350 196704 166356 196716
rect 165764 196676 166356 196704
rect 165764 196664 165770 196676
rect 166350 196664 166356 196676
rect 166408 196664 166414 196716
rect 167178 196664 167184 196716
rect 167236 196704 167242 196716
rect 201770 196704 201776 196716
rect 167236 196676 201776 196704
rect 167236 196664 167242 196676
rect 201770 196664 201776 196676
rect 201828 196664 201834 196716
rect 220814 196636 220820 196648
rect 154592 196608 220820 196636
rect 220814 196596 220820 196608
rect 220872 196596 220878 196648
rect 119522 196528 119528 196580
rect 119580 196568 119586 196580
rect 126514 196568 126520 196580
rect 119580 196540 126520 196568
rect 119580 196528 119586 196540
rect 126514 196528 126520 196540
rect 126572 196528 126578 196580
rect 129090 196528 129096 196580
rect 129148 196568 129154 196580
rect 150710 196568 150716 196580
rect 129148 196540 150716 196568
rect 129148 196528 129154 196540
rect 150710 196528 150716 196540
rect 150768 196528 150774 196580
rect 165614 196528 165620 196580
rect 165672 196568 165678 196580
rect 166442 196568 166448 196580
rect 165672 196540 166448 196568
rect 165672 196528 165678 196540
rect 166442 196528 166448 196540
rect 166500 196528 166506 196580
rect 117038 196460 117044 196512
rect 117096 196500 117102 196512
rect 123478 196500 123484 196512
rect 117096 196472 123484 196500
rect 117096 196460 117102 196472
rect 123478 196460 123484 196472
rect 123536 196460 123542 196512
rect 129734 196460 129740 196512
rect 129792 196500 129798 196512
rect 132586 196500 132592 196512
rect 129792 196472 132592 196500
rect 129792 196460 129798 196472
rect 132586 196460 132592 196472
rect 132644 196460 132650 196512
rect 157886 196460 157892 196512
rect 157944 196500 157950 196512
rect 163682 196500 163688 196512
rect 157944 196472 163688 196500
rect 157944 196460 157950 196472
rect 163682 196460 163688 196472
rect 163740 196460 163746 196512
rect 165338 196460 165344 196512
rect 165396 196500 165402 196512
rect 165890 196500 165896 196512
rect 165396 196472 165896 196500
rect 165396 196460 165402 196472
rect 165890 196460 165896 196472
rect 165948 196460 165954 196512
rect 127802 196392 127808 196444
rect 127860 196432 127866 196444
rect 140038 196432 140044 196444
rect 127860 196404 140044 196432
rect 127860 196392 127866 196404
rect 140038 196392 140044 196404
rect 140096 196392 140102 196444
rect 120350 196324 120356 196376
rect 120408 196364 120414 196376
rect 128170 196364 128176 196376
rect 120408 196336 128176 196364
rect 120408 196324 120414 196336
rect 128170 196324 128176 196336
rect 128228 196324 128234 196376
rect 150710 196324 150716 196376
rect 150768 196364 150774 196376
rect 151538 196364 151544 196376
rect 150768 196336 151544 196364
rect 150768 196324 150774 196336
rect 151538 196324 151544 196336
rect 151596 196324 151602 196376
rect 119614 196256 119620 196308
rect 119672 196296 119678 196308
rect 128078 196296 128084 196308
rect 119672 196268 128084 196296
rect 119672 196256 119678 196268
rect 128078 196256 128084 196268
rect 128136 196256 128142 196308
rect 133138 196256 133144 196308
rect 133196 196296 133202 196308
rect 138842 196296 138848 196308
rect 133196 196268 138848 196296
rect 133196 196256 133202 196268
rect 138842 196256 138848 196268
rect 138900 196256 138906 196308
rect 141234 196256 141240 196308
rect 141292 196296 141298 196308
rect 142062 196296 142068 196308
rect 141292 196268 142068 196296
rect 141292 196256 141298 196268
rect 142062 196256 142068 196268
rect 142120 196256 142126 196308
rect 143994 196256 144000 196308
rect 144052 196296 144058 196308
rect 144730 196296 144736 196308
rect 144052 196268 144736 196296
rect 144052 196256 144058 196268
rect 144730 196256 144736 196268
rect 144788 196256 144794 196308
rect 132954 196188 132960 196240
rect 133012 196228 133018 196240
rect 143074 196228 143080 196240
rect 133012 196200 143080 196228
rect 133012 196188 133018 196200
rect 143074 196188 143080 196200
rect 143132 196188 143138 196240
rect 157794 196188 157800 196240
rect 157852 196228 157858 196240
rect 157978 196228 157984 196240
rect 157852 196200 157984 196228
rect 157852 196188 157858 196200
rect 157978 196188 157984 196200
rect 158036 196188 158042 196240
rect 174446 196188 174452 196240
rect 174504 196228 174510 196240
rect 180610 196228 180616 196240
rect 174504 196200 180616 196228
rect 174504 196188 174510 196200
rect 180610 196188 180616 196200
rect 180668 196188 180674 196240
rect 177114 196120 177120 196172
rect 177172 196160 177178 196172
rect 177758 196160 177764 196172
rect 177172 196132 177764 196160
rect 177172 196120 177178 196132
rect 177758 196120 177764 196132
rect 177816 196120 177822 196172
rect 131758 196052 131764 196104
rect 131816 196092 131822 196104
rect 138934 196092 138940 196104
rect 131816 196064 138940 196092
rect 131816 196052 131822 196064
rect 138934 196052 138940 196064
rect 138992 196052 138998 196104
rect 157334 196052 157340 196104
rect 157392 196092 157398 196104
rect 157392 196064 162854 196092
rect 157392 196052 157398 196064
rect 126238 195916 126244 195968
rect 126296 195956 126302 195968
rect 145834 195956 145840 195968
rect 126296 195928 145840 195956
rect 126296 195916 126302 195928
rect 145834 195916 145840 195928
rect 145892 195916 145898 195968
rect 154022 195916 154028 195968
rect 154080 195956 154086 195968
rect 154666 195956 154672 195968
rect 154080 195928 154672 195956
rect 154080 195916 154086 195928
rect 154666 195916 154672 195928
rect 154724 195916 154730 195968
rect 154758 195916 154764 195968
rect 154816 195956 154822 195968
rect 155862 195956 155868 195968
rect 154816 195928 155868 195956
rect 154816 195916 154822 195928
rect 155862 195916 155868 195928
rect 155920 195916 155926 195968
rect 157334 195916 157340 195968
rect 157392 195956 157398 195968
rect 157518 195956 157524 195968
rect 157392 195928 157524 195956
rect 157392 195916 157398 195928
rect 157518 195916 157524 195928
rect 157576 195916 157582 195968
rect 122282 195848 122288 195900
rect 122340 195888 122346 195900
rect 140222 195888 140228 195900
rect 122340 195860 140228 195888
rect 122340 195848 122346 195860
rect 140222 195848 140228 195860
rect 140280 195848 140286 195900
rect 143442 195888 143448 195900
rect 140332 195860 143448 195888
rect 108482 195780 108488 195832
rect 108540 195820 108546 195832
rect 133046 195820 133052 195832
rect 108540 195792 133052 195820
rect 108540 195780 108546 195792
rect 133046 195780 133052 195792
rect 133104 195780 133110 195832
rect 135898 195780 135904 195832
rect 135956 195820 135962 195832
rect 136726 195820 136732 195832
rect 135956 195792 136732 195820
rect 135956 195780 135962 195792
rect 136726 195780 136732 195792
rect 136784 195780 136790 195832
rect 140332 195820 140360 195860
rect 143442 195848 143448 195860
rect 143500 195848 143506 195900
rect 152090 195848 152096 195900
rect 152148 195888 152154 195900
rect 152366 195888 152372 195900
rect 152148 195860 152372 195888
rect 152148 195848 152154 195860
rect 152366 195848 152372 195860
rect 152424 195848 152430 195900
rect 162826 195888 162854 196064
rect 162946 196052 162952 196104
rect 163004 196092 163010 196104
rect 163406 196092 163412 196104
rect 163004 196064 163412 196092
rect 163004 196052 163010 196064
rect 163406 196052 163412 196064
rect 163464 196052 163470 196104
rect 165706 195984 165712 196036
rect 165764 196024 165770 196036
rect 166718 196024 166724 196036
rect 165764 195996 166724 196024
rect 165764 195984 165770 195996
rect 166718 195984 166724 195996
rect 166776 195984 166782 196036
rect 171226 195984 171232 196036
rect 171284 196024 171290 196036
rect 171410 196024 171416 196036
rect 171284 195996 171416 196024
rect 171284 195984 171290 195996
rect 171410 195984 171416 195996
rect 171468 195984 171474 196036
rect 176930 195984 176936 196036
rect 176988 196024 176994 196036
rect 177482 196024 177488 196036
rect 176988 195996 177488 196024
rect 176988 195984 176994 195996
rect 177482 195984 177488 195996
rect 177540 195984 177546 196036
rect 164510 195916 164516 195968
rect 164568 195956 164574 195968
rect 164786 195956 164792 195968
rect 164568 195928 164792 195956
rect 164568 195916 164574 195928
rect 164786 195916 164792 195928
rect 164844 195916 164850 195968
rect 165522 195916 165528 195968
rect 165580 195956 165586 195968
rect 166166 195956 166172 195968
rect 165580 195928 166172 195956
rect 165580 195916 165586 195928
rect 166166 195916 166172 195928
rect 166224 195916 166230 195968
rect 168558 195916 168564 195968
rect 168616 195956 168622 195968
rect 185762 195956 185768 195968
rect 168616 195928 185768 195956
rect 168616 195916 168622 195928
rect 185762 195916 185768 195928
rect 185820 195916 185826 195968
rect 180426 195888 180432 195900
rect 162826 195860 180432 195888
rect 180426 195848 180432 195860
rect 180484 195848 180490 195900
rect 137940 195792 140360 195820
rect 118234 195712 118240 195764
rect 118292 195752 118298 195764
rect 135806 195752 135812 195764
rect 118292 195724 135812 195752
rect 118292 195712 118298 195724
rect 135806 195712 135812 195724
rect 135864 195712 135870 195764
rect 110230 195644 110236 195696
rect 110288 195684 110294 195696
rect 137940 195684 137968 195792
rect 140866 195780 140872 195832
rect 140924 195820 140930 195832
rect 147950 195820 147956 195832
rect 140924 195792 147956 195820
rect 140924 195780 140930 195792
rect 147950 195780 147956 195792
rect 148008 195780 148014 195832
rect 157518 195780 157524 195832
rect 157576 195820 157582 195832
rect 158438 195820 158444 195832
rect 157576 195792 158444 195820
rect 157576 195780 157582 195792
rect 158438 195780 158444 195792
rect 158496 195780 158502 195832
rect 161382 195780 161388 195832
rect 161440 195820 161446 195832
rect 161440 195792 167684 195820
rect 161440 195780 161446 195792
rect 138014 195712 138020 195764
rect 138072 195752 138078 195764
rect 149054 195752 149060 195764
rect 138072 195724 149060 195752
rect 138072 195712 138078 195724
rect 149054 195712 149060 195724
rect 149112 195712 149118 195764
rect 154666 195712 154672 195764
rect 154724 195752 154730 195764
rect 155954 195752 155960 195764
rect 154724 195724 155960 195752
rect 154724 195712 154730 195724
rect 155954 195712 155960 195724
rect 156012 195712 156018 195764
rect 156230 195712 156236 195764
rect 156288 195752 156294 195764
rect 157058 195752 157064 195764
rect 156288 195724 157064 195752
rect 156288 195712 156294 195724
rect 157058 195712 157064 195724
rect 157116 195712 157122 195764
rect 110288 195656 137968 195684
rect 110288 195644 110294 195656
rect 140222 195644 140228 195696
rect 140280 195684 140286 195696
rect 146478 195684 146484 195696
rect 140280 195656 146484 195684
rect 140280 195644 140286 195656
rect 146478 195644 146484 195656
rect 146536 195644 146542 195696
rect 167656 195684 167684 195792
rect 170030 195780 170036 195832
rect 170088 195820 170094 195832
rect 200298 195820 200304 195832
rect 170088 195792 200304 195820
rect 170088 195780 170094 195792
rect 200298 195780 200304 195792
rect 200356 195780 200362 195832
rect 171594 195712 171600 195764
rect 171652 195752 171658 195764
rect 192662 195752 192668 195764
rect 171652 195724 192668 195752
rect 171652 195712 171658 195724
rect 192662 195712 192668 195724
rect 192720 195712 192726 195764
rect 196066 195684 196072 195696
rect 167656 195656 196072 195684
rect 196066 195644 196072 195656
rect 196124 195644 196130 195696
rect 109862 195576 109868 195628
rect 109920 195616 109926 195628
rect 142890 195616 142896 195628
rect 109920 195588 142896 195616
rect 109920 195576 109926 195588
rect 142890 195576 142896 195588
rect 142948 195576 142954 195628
rect 162302 195576 162308 195628
rect 162360 195616 162366 195628
rect 171594 195616 171600 195628
rect 162360 195588 171600 195616
rect 162360 195576 162366 195588
rect 171594 195576 171600 195588
rect 171652 195576 171658 195628
rect 171704 195588 172514 195616
rect 105814 195508 105820 195560
rect 105872 195548 105878 195560
rect 133138 195548 133144 195560
rect 105872 195520 133144 195548
rect 105872 195508 105878 195520
rect 133138 195508 133144 195520
rect 133196 195508 133202 195560
rect 135806 195508 135812 195560
rect 135864 195548 135870 195560
rect 138014 195548 138020 195560
rect 135864 195520 138020 195548
rect 135864 195508 135870 195520
rect 138014 195508 138020 195520
rect 138072 195508 138078 195560
rect 159726 195508 159732 195560
rect 159784 195548 159790 195560
rect 171704 195548 171732 195588
rect 159784 195520 171732 195548
rect 172486 195548 172514 195588
rect 174446 195576 174452 195628
rect 174504 195616 174510 195628
rect 174814 195616 174820 195628
rect 174504 195588 174820 195616
rect 174504 195576 174510 195588
rect 174814 195576 174820 195588
rect 174872 195576 174878 195628
rect 179506 195576 179512 195628
rect 179564 195616 179570 195628
rect 211338 195616 211344 195628
rect 179564 195588 211344 195616
rect 179564 195576 179570 195588
rect 211338 195576 211344 195588
rect 211396 195576 211402 195628
rect 193214 195548 193220 195560
rect 172486 195520 193220 195548
rect 159784 195508 159790 195520
rect 193214 195508 193220 195520
rect 193272 195508 193278 195560
rect 112438 195440 112444 195492
rect 112496 195480 112502 195492
rect 145558 195480 145564 195492
rect 112496 195452 145564 195480
rect 112496 195440 112502 195452
rect 145558 195440 145564 195452
rect 145616 195440 145622 195492
rect 151906 195440 151912 195492
rect 151964 195480 151970 195492
rect 152090 195480 152096 195492
rect 151964 195452 152096 195480
rect 151964 195440 151970 195452
rect 152090 195440 152096 195452
rect 152148 195440 152154 195492
rect 158714 195440 158720 195492
rect 158772 195480 158778 195492
rect 159818 195480 159824 195492
rect 158772 195452 159824 195480
rect 158772 195440 158778 195452
rect 159818 195440 159824 195452
rect 159876 195440 159882 195492
rect 165062 195440 165068 195492
rect 165120 195480 165126 195492
rect 198918 195480 198924 195492
rect 165120 195452 198924 195480
rect 165120 195440 165126 195452
rect 198918 195440 198924 195452
rect 198976 195440 198982 195492
rect 114370 195372 114376 195424
rect 114428 195412 114434 195424
rect 148778 195412 148784 195424
rect 114428 195384 148784 195412
rect 114428 195372 114434 195384
rect 148778 195372 148784 195384
rect 148836 195372 148842 195424
rect 149514 195372 149520 195424
rect 149572 195412 149578 195424
rect 149974 195412 149980 195424
rect 149572 195384 149980 195412
rect 149572 195372 149578 195384
rect 149974 195372 149980 195384
rect 150032 195372 150038 195424
rect 161198 195372 161204 195424
rect 161256 195412 161262 195424
rect 194686 195412 194692 195424
rect 161256 195384 194692 195412
rect 161256 195372 161262 195384
rect 194686 195372 194692 195384
rect 194744 195372 194750 195424
rect 111242 195304 111248 195356
rect 111300 195344 111306 195356
rect 145926 195344 145932 195356
rect 111300 195316 145932 195344
rect 111300 195304 111306 195316
rect 145926 195304 145932 195316
rect 145984 195304 145990 195356
rect 149606 195304 149612 195356
rect 149664 195344 149670 195356
rect 150158 195344 150164 195356
rect 149664 195316 150164 195344
rect 149664 195304 149670 195316
rect 150158 195304 150164 195316
rect 150216 195304 150222 195356
rect 156046 195304 156052 195356
rect 156104 195344 156110 195356
rect 156506 195344 156512 195356
rect 156104 195316 156512 195344
rect 156104 195304 156110 195316
rect 156506 195304 156512 195316
rect 156564 195304 156570 195356
rect 160370 195304 160376 195356
rect 160428 195344 160434 195356
rect 160428 195316 164234 195344
rect 160428 195304 160434 195316
rect 111334 195236 111340 195288
rect 111392 195276 111398 195288
rect 144270 195276 144276 195288
rect 111392 195248 144276 195276
rect 111392 195236 111398 195248
rect 144270 195236 144276 195248
rect 144328 195236 144334 195288
rect 146938 195236 146944 195288
rect 146996 195276 147002 195288
rect 152734 195276 152740 195288
rect 146996 195248 152740 195276
rect 146996 195236 147002 195248
rect 152734 195236 152740 195248
rect 152792 195236 152798 195288
rect 158898 195236 158904 195288
rect 158956 195276 158962 195288
rect 159910 195276 159916 195288
rect 158956 195248 159916 195276
rect 158956 195236 158962 195248
rect 159910 195236 159916 195248
rect 159968 195236 159974 195288
rect 164206 195276 164234 195316
rect 175182 195304 175188 195356
rect 175240 195344 175246 195356
rect 175366 195344 175372 195356
rect 175240 195316 175372 195344
rect 175240 195304 175246 195316
rect 175366 195304 175372 195316
rect 175424 195304 175430 195356
rect 180518 195304 180524 195356
rect 180576 195344 180582 195356
rect 210326 195344 210332 195356
rect 180576 195316 210332 195344
rect 180576 195304 180582 195316
rect 210326 195304 210332 195316
rect 210384 195304 210390 195356
rect 214558 195276 214564 195288
rect 164206 195248 214564 195276
rect 214558 195236 214564 195248
rect 214616 195236 214622 195288
rect 129274 195168 129280 195220
rect 129332 195208 129338 195220
rect 140866 195208 140872 195220
rect 129332 195180 140872 195208
rect 129332 195168 129338 195180
rect 140866 195168 140872 195180
rect 140924 195168 140930 195220
rect 166534 195168 166540 195220
rect 166592 195208 166598 195220
rect 181438 195208 181444 195220
rect 166592 195180 181444 195208
rect 166592 195168 166598 195180
rect 181438 195168 181444 195180
rect 181496 195168 181502 195220
rect 140498 195100 140504 195152
rect 140556 195140 140562 195152
rect 143626 195140 143632 195152
rect 140556 195112 143632 195140
rect 140556 195100 140562 195112
rect 143626 195100 143632 195112
rect 143684 195100 143690 195152
rect 160462 195100 160468 195152
rect 160520 195140 160526 195152
rect 161290 195140 161296 195152
rect 160520 195112 161296 195140
rect 160520 195100 160526 195112
rect 161290 195100 161296 195112
rect 161348 195100 161354 195152
rect 168374 195100 168380 195152
rect 168432 195140 168438 195152
rect 169386 195140 169392 195152
rect 168432 195112 169392 195140
rect 168432 195100 168438 195112
rect 169386 195100 169392 195112
rect 169444 195100 169450 195152
rect 171318 195100 171324 195152
rect 171376 195140 171382 195152
rect 172238 195140 172244 195152
rect 171376 195112 172244 195140
rect 171376 195100 171382 195112
rect 172238 195100 172244 195112
rect 172296 195100 172302 195152
rect 132402 195032 132408 195084
rect 132460 195072 132466 195084
rect 144178 195072 144184 195084
rect 132460 195044 144184 195072
rect 132460 195032 132466 195044
rect 144178 195032 144184 195044
rect 144236 195032 144242 195084
rect 152182 195032 152188 195084
rect 152240 195072 152246 195084
rect 152918 195072 152924 195084
rect 152240 195044 152924 195072
rect 152240 195032 152246 195044
rect 152918 195032 152924 195044
rect 152976 195032 152982 195084
rect 160186 194896 160192 194948
rect 160244 194936 160250 194948
rect 160738 194936 160744 194948
rect 160244 194908 160744 194936
rect 160244 194896 160250 194908
rect 160738 194896 160744 194908
rect 160796 194896 160802 194948
rect 166626 194896 166632 194948
rect 166684 194936 166690 194948
rect 183094 194936 183100 194948
rect 166684 194908 183100 194936
rect 166684 194896 166690 194908
rect 183094 194896 183100 194908
rect 183152 194896 183158 194948
rect 156322 194828 156328 194880
rect 156380 194868 156386 194880
rect 156966 194868 156972 194880
rect 156380 194840 156972 194868
rect 156380 194828 156386 194840
rect 156966 194828 156972 194840
rect 157024 194828 157030 194880
rect 133138 194760 133144 194812
rect 133196 194800 133202 194812
rect 139118 194800 139124 194812
rect 133196 194772 139124 194800
rect 133196 194760 133202 194772
rect 139118 194760 139124 194772
rect 139176 194760 139182 194812
rect 164326 194760 164332 194812
rect 164384 194800 164390 194812
rect 164878 194800 164884 194812
rect 164384 194772 164884 194800
rect 164384 194760 164390 194772
rect 164878 194760 164884 194772
rect 164936 194760 164942 194812
rect 132218 194692 132224 194744
rect 132276 194732 132282 194744
rect 138474 194732 138480 194744
rect 132276 194704 138480 194732
rect 132276 194692 132282 194704
rect 138474 194692 138480 194704
rect 138532 194692 138538 194744
rect 151906 194692 151912 194744
rect 151964 194732 151970 194744
rect 152642 194732 152648 194744
rect 151964 194704 152648 194732
rect 151964 194692 151970 194704
rect 152642 194692 152648 194704
rect 152700 194692 152706 194744
rect 117774 194488 117780 194540
rect 117832 194528 117838 194540
rect 120810 194528 120816 194540
rect 117832 194500 120816 194528
rect 117832 194488 117838 194500
rect 120810 194488 120816 194500
rect 120868 194488 120874 194540
rect 141050 194488 141056 194540
rect 141108 194528 141114 194540
rect 143534 194528 143540 194540
rect 141108 194500 143540 194528
rect 141108 194488 141114 194500
rect 143534 194488 143540 194500
rect 143592 194488 143598 194540
rect 165522 194488 165528 194540
rect 165580 194528 165586 194540
rect 167362 194528 167368 194540
rect 165580 194500 167368 194528
rect 165580 194488 165586 194500
rect 167362 194488 167368 194500
rect 167420 194488 167426 194540
rect 147766 194420 147772 194472
rect 147824 194460 147830 194472
rect 148226 194460 148232 194472
rect 147824 194432 148232 194460
rect 147824 194420 147830 194432
rect 148226 194420 148232 194432
rect 148284 194420 148290 194472
rect 130378 194352 130384 194404
rect 130436 194392 130442 194404
rect 147674 194392 147680 194404
rect 130436 194364 147680 194392
rect 130436 194352 130442 194364
rect 147674 194352 147680 194364
rect 147732 194352 147738 194404
rect 173158 194352 173164 194404
rect 173216 194392 173222 194404
rect 207198 194392 207204 194404
rect 173216 194364 207204 194392
rect 173216 194352 173222 194364
rect 207198 194352 207204 194364
rect 207256 194352 207262 194404
rect 108666 194284 108672 194336
rect 108724 194324 108730 194336
rect 140682 194324 140688 194336
rect 108724 194296 140688 194324
rect 108724 194284 108730 194296
rect 140682 194284 140688 194296
rect 140740 194284 140746 194336
rect 175090 194284 175096 194336
rect 175148 194324 175154 194336
rect 208670 194324 208676 194336
rect 175148 194296 208676 194324
rect 175148 194284 175154 194296
rect 208670 194284 208676 194296
rect 208728 194284 208734 194336
rect 109678 194216 109684 194268
rect 109736 194256 109742 194268
rect 109736 194228 140452 194256
rect 109736 194216 109742 194228
rect 108298 194148 108304 194200
rect 108356 194188 108362 194200
rect 140314 194188 140320 194200
rect 108356 194160 140320 194188
rect 108356 194148 108362 194160
rect 140314 194148 140320 194160
rect 140372 194148 140378 194200
rect 140424 194188 140452 194228
rect 147950 194216 147956 194268
rect 148008 194256 148014 194268
rect 148594 194256 148600 194268
rect 148008 194228 148600 194256
rect 148008 194216 148014 194228
rect 148594 194216 148600 194228
rect 148652 194216 148658 194268
rect 175734 194216 175740 194268
rect 175792 194256 175798 194268
rect 210142 194256 210148 194268
rect 175792 194228 210148 194256
rect 175792 194216 175798 194228
rect 210142 194216 210148 194228
rect 210200 194216 210206 194268
rect 141878 194188 141884 194200
rect 140424 194160 141884 194188
rect 141878 194148 141884 194160
rect 141936 194148 141942 194200
rect 179874 194148 179880 194200
rect 179932 194188 179938 194200
rect 207382 194188 207388 194200
rect 179932 194160 207388 194188
rect 179932 194148 179938 194160
rect 207382 194148 207388 194160
rect 207440 194148 207446 194200
rect 100478 194080 100484 194132
rect 100536 194120 100542 194132
rect 126974 194120 126980 194132
rect 100536 194092 126980 194120
rect 100536 194080 100542 194092
rect 126974 194080 126980 194092
rect 127032 194080 127038 194132
rect 174078 194080 174084 194132
rect 174136 194120 174142 194132
rect 208762 194120 208768 194132
rect 174136 194092 208768 194120
rect 174136 194080 174142 194092
rect 208762 194080 208768 194092
rect 208820 194080 208826 194132
rect 103330 194012 103336 194064
rect 103388 194052 103394 194064
rect 135530 194052 135536 194064
rect 103388 194024 135536 194052
rect 103388 194012 103394 194024
rect 135530 194012 135536 194024
rect 135588 194012 135594 194064
rect 158990 194012 158996 194064
rect 159048 194052 159054 194064
rect 176010 194052 176016 194064
rect 159048 194024 176016 194052
rect 159048 194012 159054 194024
rect 176010 194012 176016 194024
rect 176068 194012 176074 194064
rect 177022 194012 177028 194064
rect 177080 194052 177086 194064
rect 177574 194052 177580 194064
rect 177080 194024 177580 194052
rect 177080 194012 177086 194024
rect 177574 194012 177580 194024
rect 177632 194012 177638 194064
rect 179414 194012 179420 194064
rect 179472 194052 179478 194064
rect 211798 194052 211804 194064
rect 179472 194024 211804 194052
rect 179472 194012 179478 194024
rect 211798 194012 211804 194024
rect 211856 194012 211862 194064
rect 108758 193944 108764 193996
rect 108816 193984 108822 193996
rect 143166 193984 143172 193996
rect 108816 193956 143172 193984
rect 108816 193944 108822 193956
rect 143166 193944 143172 193956
rect 143224 193944 143230 193996
rect 158806 193944 158812 193996
rect 158864 193984 158870 193996
rect 159542 193984 159548 193996
rect 158864 193956 159548 193984
rect 158864 193944 158870 193956
rect 159542 193944 159548 193956
rect 159600 193944 159606 193996
rect 162118 193944 162124 193996
rect 162176 193984 162182 193996
rect 174814 193984 174820 193996
rect 162176 193956 174820 193984
rect 162176 193944 162182 193956
rect 174814 193944 174820 193956
rect 174872 193944 174878 193996
rect 175458 193944 175464 193996
rect 175516 193984 175522 193996
rect 210510 193984 210516 193996
rect 175516 193956 210516 193984
rect 175516 193944 175522 193956
rect 210510 193944 210516 193956
rect 210568 193944 210574 193996
rect 104342 193876 104348 193928
rect 104400 193916 104406 193928
rect 139302 193916 139308 193928
rect 104400 193888 139308 193916
rect 104400 193876 104406 193888
rect 139302 193876 139308 193888
rect 139360 193876 139366 193928
rect 151814 193876 151820 193928
rect 151872 193916 151878 193928
rect 171594 193916 171600 193928
rect 151872 193888 171600 193916
rect 151872 193876 151878 193888
rect 171594 193876 171600 193888
rect 171652 193876 171658 193928
rect 174538 193876 174544 193928
rect 174596 193916 174602 193928
rect 214374 193916 214380 193928
rect 174596 193888 214380 193916
rect 174596 193876 174602 193888
rect 214374 193876 214380 193888
rect 214432 193876 214438 193928
rect 96430 193808 96436 193860
rect 96488 193848 96494 193860
rect 135990 193848 135996 193860
rect 96488 193820 135996 193848
rect 96488 193808 96494 193820
rect 135990 193808 135996 193820
rect 136048 193808 136054 193860
rect 141326 193808 141332 193860
rect 141384 193848 141390 193860
rect 143902 193848 143908 193860
rect 141384 193820 143908 193848
rect 141384 193808 141390 193820
rect 143902 193808 143908 193820
rect 143960 193808 143966 193860
rect 169570 193808 169576 193860
rect 169628 193848 169634 193860
rect 221366 193848 221372 193860
rect 169628 193820 221372 193848
rect 169628 193808 169634 193820
rect 221366 193808 221372 193820
rect 221424 193808 221430 193860
rect 156506 193332 156512 193384
rect 156564 193372 156570 193384
rect 157242 193372 157248 193384
rect 156564 193344 157248 193372
rect 156564 193332 156570 193344
rect 157242 193332 157248 193344
rect 157300 193332 157306 193384
rect 119522 193128 119528 193180
rect 119580 193168 119586 193180
rect 143718 193168 143724 193180
rect 119580 193140 143724 193168
rect 119580 193128 119586 193140
rect 143718 193128 143724 193140
rect 143776 193128 143782 193180
rect 157702 193128 157708 193180
rect 157760 193168 157766 193180
rect 158254 193168 158260 193180
rect 157760 193140 158260 193168
rect 157760 193128 157766 193140
rect 158254 193128 158260 193140
rect 158312 193128 158318 193180
rect 166810 193128 166816 193180
rect 166868 193168 166874 193180
rect 200206 193168 200212 193180
rect 166868 193140 200212 193168
rect 166868 193128 166874 193140
rect 200206 193128 200212 193140
rect 200264 193128 200270 193180
rect 119430 193060 119436 193112
rect 119488 193100 119494 193112
rect 145282 193100 145288 193112
rect 119488 193072 145288 193100
rect 119488 193060 119494 193072
rect 145282 193060 145288 193072
rect 145340 193060 145346 193112
rect 163130 193060 163136 193112
rect 163188 193100 163194 193112
rect 163958 193100 163964 193112
rect 163188 193072 163964 193100
rect 163188 193060 163194 193072
rect 163958 193060 163964 193072
rect 164016 193060 164022 193112
rect 167454 193060 167460 193112
rect 167512 193100 167518 193112
rect 201678 193100 201684 193112
rect 167512 193072 201684 193100
rect 167512 193060 167518 193072
rect 201678 193060 201684 193072
rect 201736 193060 201742 193112
rect 123938 192992 123944 193044
rect 123996 193032 124002 193044
rect 153194 193032 153200 193044
rect 123996 193004 153200 193032
rect 123996 192992 124002 193004
rect 153194 192992 153200 193004
rect 153252 192992 153258 193044
rect 170398 192992 170404 193044
rect 170456 193032 170462 193044
rect 204254 193032 204260 193044
rect 170456 193004 204260 193032
rect 170456 192992 170462 193004
rect 204254 192992 204260 193004
rect 204312 192992 204318 193044
rect 112714 192924 112720 192976
rect 112772 192964 112778 192976
rect 146202 192964 146208 192976
rect 112772 192936 146208 192964
rect 112772 192924 112778 192936
rect 146202 192924 146208 192936
rect 146260 192924 146266 192976
rect 153286 192924 153292 192976
rect 153344 192964 153350 192976
rect 153470 192964 153476 192976
rect 153344 192936 153476 192964
rect 153344 192924 153350 192936
rect 153470 192924 153476 192936
rect 153528 192924 153534 192976
rect 169202 192924 169208 192976
rect 169260 192964 169266 192976
rect 203058 192964 203064 192976
rect 169260 192936 203064 192964
rect 169260 192924 169266 192936
rect 203058 192924 203064 192936
rect 203116 192924 203122 192976
rect 101674 192856 101680 192908
rect 101732 192896 101738 192908
rect 135162 192896 135168 192908
rect 101732 192868 135168 192896
rect 101732 192856 101738 192868
rect 135162 192856 135168 192868
rect 135220 192856 135226 192908
rect 169938 192856 169944 192908
rect 169996 192896 170002 192908
rect 204438 192896 204444 192908
rect 169996 192868 204444 192896
rect 169996 192856 170002 192868
rect 204438 192856 204444 192868
rect 204496 192856 204502 192908
rect 101766 192788 101772 192840
rect 101824 192828 101830 192840
rect 134978 192828 134984 192840
rect 101824 192800 134984 192828
rect 101824 192788 101830 192800
rect 134978 192788 134984 192800
rect 135036 192788 135042 192840
rect 171502 192788 171508 192840
rect 171560 192828 171566 192840
rect 205634 192828 205640 192840
rect 171560 192800 205640 192828
rect 171560 192788 171566 192800
rect 205634 192788 205640 192800
rect 205692 192788 205698 192840
rect 108574 192720 108580 192772
rect 108632 192760 108638 192772
rect 142798 192760 142804 192772
rect 108632 192732 142804 192760
rect 108632 192720 108638 192732
rect 142798 192720 142804 192732
rect 142856 192720 142862 192772
rect 170122 192720 170128 192772
rect 170180 192760 170186 192772
rect 204346 192760 204352 192772
rect 170180 192732 204352 192760
rect 170180 192720 170186 192732
rect 204346 192720 204352 192732
rect 204404 192720 204410 192772
rect 108206 192652 108212 192704
rect 108264 192692 108270 192704
rect 142614 192692 142620 192704
rect 108264 192664 142620 192692
rect 108264 192652 108270 192664
rect 142614 192652 142620 192664
rect 142672 192652 142678 192704
rect 170674 192652 170680 192704
rect 170732 192692 170738 192704
rect 204530 192692 204536 192704
rect 170732 192664 204536 192692
rect 170732 192652 170738 192664
rect 204530 192652 204536 192664
rect 204588 192652 204594 192704
rect 112254 192584 112260 192636
rect 112312 192624 112318 192636
rect 146570 192624 146576 192636
rect 112312 192596 146576 192624
rect 112312 192584 112318 192596
rect 146570 192584 146576 192596
rect 146628 192584 146634 192636
rect 172146 192584 172152 192636
rect 172204 192624 172210 192636
rect 205818 192624 205824 192636
rect 172204 192596 205824 192624
rect 172204 192584 172210 192596
rect 205818 192584 205824 192596
rect 205876 192584 205882 192636
rect 97810 192516 97816 192568
rect 97868 192556 97874 192568
rect 143810 192556 143816 192568
rect 97868 192528 143816 192556
rect 97868 192516 97874 192528
rect 143810 192516 143816 192528
rect 143868 192516 143874 192568
rect 162486 192516 162492 192568
rect 162544 192556 162550 192568
rect 171962 192556 171968 192568
rect 162544 192528 171968 192556
rect 162544 192516 162550 192528
rect 171962 192516 171968 192528
rect 172020 192516 172026 192568
rect 172974 192516 172980 192568
rect 173032 192556 173038 192568
rect 207474 192556 207480 192568
rect 173032 192528 207480 192556
rect 173032 192516 173038 192528
rect 207474 192516 207480 192528
rect 207532 192516 207538 192568
rect 97442 192448 97448 192500
rect 97500 192488 97506 192500
rect 150526 192488 150532 192500
rect 97500 192460 150532 192488
rect 97500 192448 97506 192460
rect 150526 192448 150532 192460
rect 150584 192448 150590 192500
rect 155218 192448 155224 192500
rect 155276 192488 155282 192500
rect 216858 192488 216864 192500
rect 155276 192460 216864 192488
rect 155276 192448 155282 192460
rect 216858 192448 216864 192460
rect 216916 192448 216922 192500
rect 129366 192380 129372 192432
rect 129424 192420 129430 192432
rect 150250 192420 150256 192432
rect 129424 192392 150256 192420
rect 129424 192380 129430 192392
rect 150250 192380 150256 192392
rect 150308 192380 150314 192432
rect 164970 192380 164976 192432
rect 165028 192420 165034 192432
rect 174538 192420 174544 192432
rect 165028 192392 174544 192420
rect 165028 192380 165034 192392
rect 174538 192380 174544 192392
rect 174596 192380 174602 192432
rect 174630 192380 174636 192432
rect 174688 192420 174694 192432
rect 202414 192420 202420 192432
rect 174688 192392 202420 192420
rect 174688 192380 174694 192392
rect 202414 192380 202420 192392
rect 202472 192380 202478 192432
rect 130470 192312 130476 192364
rect 130528 192352 130534 192364
rect 149146 192352 149152 192364
rect 130528 192324 149152 192352
rect 130528 192312 130534 192324
rect 149146 192312 149152 192324
rect 149204 192312 149210 192364
rect 171778 192312 171784 192364
rect 171836 192352 171842 192364
rect 183186 192352 183192 192364
rect 171836 192324 183192 192352
rect 171836 192312 171842 192324
rect 183186 192312 183192 192324
rect 183244 192312 183250 192364
rect 130746 192244 130752 192296
rect 130804 192284 130810 192296
rect 147490 192284 147496 192296
rect 130804 192256 147496 192284
rect 130804 192244 130810 192256
rect 147490 192244 147496 192256
rect 147548 192244 147554 192296
rect 108850 191564 108856 191616
rect 108908 191604 108914 191616
rect 141050 191604 141056 191616
rect 108908 191576 141056 191604
rect 108908 191564 108914 191576
rect 141050 191564 141056 191576
rect 141108 191564 141114 191616
rect 104802 191496 104808 191548
rect 104860 191536 104866 191548
rect 137646 191536 137652 191548
rect 104860 191508 137652 191536
rect 104860 191496 104866 191508
rect 137646 191496 137652 191508
rect 137704 191496 137710 191548
rect 153286 191496 153292 191548
rect 153344 191536 153350 191548
rect 154298 191536 154304 191548
rect 153344 191508 154304 191536
rect 153344 191496 153350 191508
rect 154298 191496 154304 191508
rect 154356 191496 154362 191548
rect 107470 191428 107476 191480
rect 107528 191468 107534 191480
rect 139486 191468 139492 191480
rect 107528 191440 139492 191468
rect 107528 191428 107534 191440
rect 139486 191428 139492 191440
rect 139544 191428 139550 191480
rect 166966 191440 176654 191468
rect 116762 191360 116768 191412
rect 116820 191400 116826 191412
rect 149790 191400 149796 191412
rect 116820 191372 149796 191400
rect 116820 191360 116826 191372
rect 149790 191360 149796 191372
rect 149848 191360 149854 191412
rect 99190 191292 99196 191344
rect 99248 191332 99254 191344
rect 132770 191332 132776 191344
rect 99248 191304 132776 191332
rect 99248 191292 99254 191304
rect 132770 191292 132776 191304
rect 132828 191292 132834 191344
rect 160830 191292 160836 191344
rect 160888 191332 160894 191344
rect 166966 191332 166994 191440
rect 160888 191304 166994 191332
rect 160888 191292 160894 191304
rect 167086 191292 167092 191344
rect 167144 191332 167150 191344
rect 176626 191332 176654 191440
rect 188338 191332 188344 191344
rect 167144 191304 176516 191332
rect 176626 191304 188344 191332
rect 167144 191292 167150 191304
rect 103054 191224 103060 191276
rect 103112 191264 103118 191276
rect 137462 191264 137468 191276
rect 103112 191236 137468 191264
rect 103112 191224 103118 191236
rect 137462 191224 137468 191236
rect 137520 191224 137526 191276
rect 167178 191224 167184 191276
rect 167236 191264 167242 191276
rect 168006 191264 168012 191276
rect 167236 191236 168012 191264
rect 167236 191224 167242 191236
rect 168006 191224 168012 191236
rect 168064 191224 168070 191276
rect 171410 191224 171416 191276
rect 171468 191264 171474 191276
rect 172238 191264 172244 191276
rect 171468 191236 172244 191264
rect 171468 191224 171474 191236
rect 172238 191224 172244 191236
rect 172296 191224 172302 191276
rect 175550 191224 175556 191276
rect 175608 191264 175614 191276
rect 176378 191264 176384 191276
rect 175608 191236 176384 191264
rect 175608 191224 175614 191236
rect 176378 191224 176384 191236
rect 176436 191224 176442 191276
rect 176488 191264 176516 191304
rect 188338 191292 188344 191304
rect 188396 191292 188402 191344
rect 201494 191264 201500 191276
rect 176488 191236 201500 191264
rect 201494 191224 201500 191236
rect 201552 191224 201558 191276
rect 99098 191156 99104 191208
rect 99156 191196 99162 191208
rect 146754 191196 146760 191208
rect 99156 191168 146760 191196
rect 99156 191156 99162 191168
rect 146754 191156 146760 191168
rect 146812 191156 146818 191208
rect 166350 191156 166356 191208
rect 166408 191196 166414 191208
rect 200482 191196 200488 191208
rect 166408 191168 200488 191196
rect 166408 191156 166414 191168
rect 200482 191156 200488 191168
rect 200540 191156 200546 191208
rect 99006 191088 99012 191140
rect 99064 191128 99070 191140
rect 99064 191100 138014 191128
rect 99064 191088 99070 191100
rect 133046 191020 133052 191072
rect 133104 191060 133110 191072
rect 133782 191060 133788 191072
rect 133104 191032 133788 191060
rect 133104 191020 133110 191032
rect 133782 191020 133788 191032
rect 133840 191020 133846 191072
rect 135714 191020 135720 191072
rect 135772 191060 135778 191072
rect 136082 191060 136088 191072
rect 135772 191032 136088 191060
rect 135772 191020 135778 191032
rect 136082 191020 136088 191032
rect 136140 191020 136146 191072
rect 137986 191060 138014 191100
rect 138382 191088 138388 191140
rect 138440 191128 138446 191140
rect 139210 191128 139216 191140
rect 138440 191100 139216 191128
rect 138440 191088 138446 191100
rect 139210 191088 139216 191100
rect 139268 191088 139274 191140
rect 140222 191088 140228 191140
rect 140280 191128 140286 191140
rect 140590 191128 140596 191140
rect 140280 191100 140596 191128
rect 140280 191088 140286 191100
rect 140590 191088 140596 191100
rect 140648 191088 140654 191140
rect 163222 191088 163228 191140
rect 163280 191128 163286 191140
rect 211614 191128 211620 191140
rect 163280 191100 211620 191128
rect 163280 191088 163286 191100
rect 211614 191088 211620 191100
rect 211672 191088 211678 191140
rect 146846 191060 146852 191072
rect 137986 191032 146852 191060
rect 146846 191020 146852 191032
rect 146904 191020 146910 191072
rect 167822 191020 167828 191072
rect 167880 191060 167886 191072
rect 168006 191060 168012 191072
rect 167880 191032 168012 191060
rect 167880 191020 167886 191032
rect 168006 191020 168012 191032
rect 168064 191020 168070 191072
rect 169754 191020 169760 191072
rect 169812 191060 169818 191072
rect 170858 191060 170864 191072
rect 169812 191032 170864 191060
rect 169812 191020 169818 191032
rect 170858 191020 170864 191032
rect 170916 191020 170922 191072
rect 171134 191020 171140 191072
rect 171192 191060 171198 191072
rect 171686 191060 171692 191072
rect 171192 191032 171692 191060
rect 171192 191020 171198 191032
rect 171686 191020 171692 191032
rect 171744 191020 171750 191072
rect 172606 191020 172612 191072
rect 172664 191060 172670 191072
rect 173618 191060 173624 191072
rect 172664 191032 173624 191060
rect 172664 191020 172670 191032
rect 173618 191020 173624 191032
rect 173676 191020 173682 191072
rect 175458 191020 175464 191072
rect 175516 191060 175522 191072
rect 176102 191060 176108 191072
rect 175516 191032 176108 191060
rect 175516 191020 175522 191032
rect 176102 191020 176108 191032
rect 176160 191020 176166 191072
rect 167086 190952 167092 191004
rect 167144 190992 167150 191004
rect 168098 190992 168104 191004
rect 167144 190964 168104 190992
rect 167144 190952 167150 190964
rect 168098 190952 168104 190964
rect 168156 190952 168162 191004
rect 142614 190884 142620 190936
rect 142672 190924 142678 190936
rect 142982 190924 142988 190936
rect 142672 190896 142988 190924
rect 142672 190884 142678 190896
rect 142982 190884 142988 190896
rect 143040 190884 143046 190936
rect 167638 190884 167644 190936
rect 167696 190924 167702 190936
rect 168282 190924 168288 190936
rect 167696 190896 168288 190924
rect 167696 190884 167702 190896
rect 168282 190884 168288 190896
rect 168340 190884 168346 190936
rect 174170 190884 174176 190936
rect 174228 190924 174234 190936
rect 174722 190924 174728 190936
rect 174228 190896 174728 190924
rect 174228 190884 174234 190896
rect 174722 190884 174728 190896
rect 174780 190884 174786 190936
rect 132126 190680 132132 190732
rect 132184 190680 132190 190732
rect 132144 190528 132172 190680
rect 132126 190476 132132 190528
rect 132184 190476 132190 190528
rect 155494 190408 155500 190460
rect 155552 190448 155558 190460
rect 185670 190448 185676 190460
rect 155552 190420 185676 190448
rect 155552 190408 155558 190420
rect 185670 190408 185676 190420
rect 185728 190408 185734 190460
rect 132034 190340 132040 190392
rect 132092 190380 132098 190392
rect 132218 190380 132224 190392
rect 132092 190352 132224 190380
rect 132092 190340 132098 190352
rect 132218 190340 132224 190352
rect 132276 190340 132282 190392
rect 132310 190340 132316 190392
rect 132368 190380 132374 190392
rect 132494 190380 132500 190392
rect 132368 190352 132500 190380
rect 132368 190340 132374 190352
rect 132494 190340 132500 190352
rect 132552 190340 132558 190392
rect 173710 190340 173716 190392
rect 173768 190380 173774 190392
rect 205726 190380 205732 190392
rect 173768 190352 205732 190380
rect 173768 190340 173774 190352
rect 205726 190340 205732 190352
rect 205784 190340 205790 190392
rect 120810 190272 120816 190324
rect 120868 190312 120874 190324
rect 151078 190312 151084 190324
rect 120868 190284 151084 190312
rect 120868 190272 120874 190284
rect 151078 190272 151084 190284
rect 151136 190272 151142 190324
rect 174446 190272 174452 190324
rect 174504 190312 174510 190324
rect 208578 190312 208584 190324
rect 174504 190284 208584 190312
rect 174504 190272 174510 190284
rect 208578 190272 208584 190284
rect 208636 190272 208642 190324
rect 106090 190204 106096 190256
rect 106148 190244 106154 190256
rect 137186 190244 137192 190256
rect 106148 190216 137192 190244
rect 106148 190204 106154 190216
rect 137186 190204 137192 190216
rect 137244 190204 137250 190256
rect 176470 190204 176476 190256
rect 176528 190244 176534 190256
rect 210234 190244 210240 190256
rect 176528 190216 210240 190244
rect 176528 190204 176534 190216
rect 210234 190204 210240 190216
rect 210292 190204 210298 190256
rect 103238 190136 103244 190188
rect 103296 190176 103302 190188
rect 136358 190176 136364 190188
rect 103296 190148 136364 190176
rect 103296 190136 103302 190148
rect 136358 190136 136364 190148
rect 136416 190136 136422 190188
rect 177298 190136 177304 190188
rect 177356 190176 177362 190188
rect 211706 190176 211712 190188
rect 177356 190148 211712 190176
rect 177356 190136 177362 190148
rect 211706 190136 211712 190148
rect 211764 190136 211770 190188
rect 110138 190068 110144 190120
rect 110196 190108 110202 190120
rect 144546 190108 144552 190120
rect 110196 190080 144552 190108
rect 110196 190068 110202 190080
rect 144546 190068 144552 190080
rect 144604 190068 144610 190120
rect 157886 190068 157892 190120
rect 157944 190108 157950 190120
rect 202322 190108 202328 190120
rect 157944 190080 202328 190108
rect 157944 190068 157950 190080
rect 202322 190068 202328 190080
rect 202380 190068 202386 190120
rect 110046 190000 110052 190052
rect 110104 190040 110110 190052
rect 144086 190040 144092 190052
rect 110104 190012 144092 190040
rect 110104 190000 110110 190012
rect 144086 190000 144092 190012
rect 144144 190000 144150 190052
rect 158990 190000 158996 190052
rect 159048 190040 159054 190052
rect 207014 190040 207020 190052
rect 159048 190012 207020 190040
rect 159048 190000 159054 190012
rect 207014 190000 207020 190012
rect 207072 190000 207078 190052
rect 101858 189932 101864 189984
rect 101916 189972 101922 189984
rect 135990 189972 135996 189984
rect 101916 189944 135996 189972
rect 101916 189932 101922 189944
rect 135990 189932 135996 189944
rect 136048 189932 136054 189984
rect 137278 189932 137284 189984
rect 137336 189972 137342 189984
rect 137462 189972 137468 189984
rect 137336 189944 137468 189972
rect 137336 189932 137342 189944
rect 137462 189932 137468 189944
rect 137520 189932 137526 189984
rect 157794 189932 157800 189984
rect 157852 189972 157858 189984
rect 219618 189972 219624 189984
rect 157852 189944 219624 189972
rect 157852 189932 157858 189944
rect 219618 189932 219624 189944
rect 219676 189932 219682 189984
rect 108114 189864 108120 189916
rect 108172 189904 108178 189916
rect 143902 189904 143908 189916
rect 108172 189876 143908 189904
rect 108172 189864 108178 189876
rect 143902 189864 143908 189876
rect 143960 189864 143966 189916
rect 157978 189864 157984 189916
rect 158036 189904 158042 189916
rect 221090 189904 221096 189916
rect 158036 189876 221096 189904
rect 158036 189864 158042 189876
rect 221090 189864 221096 189876
rect 221148 189864 221154 189916
rect 97350 189796 97356 189848
rect 97408 189836 97414 189848
rect 144822 189836 144828 189848
rect 97408 189808 144828 189836
rect 97408 189796 97414 189808
rect 144822 189796 144828 189808
rect 144880 189796 144886 189848
rect 156506 189796 156512 189848
rect 156564 189836 156570 189848
rect 220998 189836 221004 189848
rect 156564 189808 221004 189836
rect 156564 189796 156570 189808
rect 220998 189796 221004 189808
rect 221056 189796 221062 189848
rect 96338 189728 96344 189780
rect 96396 189768 96402 189780
rect 149514 189768 149520 189780
rect 96396 189740 149520 189768
rect 96396 189728 96402 189740
rect 149514 189728 149520 189740
rect 149572 189728 149578 189780
rect 156414 189728 156420 189780
rect 156472 189768 156478 189780
rect 221182 189768 221188 189780
rect 156472 189740 221188 189768
rect 156472 189728 156478 189740
rect 221182 189728 221188 189740
rect 221240 189728 221246 189780
rect 159634 189660 159640 189712
rect 159692 189700 159698 189712
rect 185854 189700 185860 189712
rect 159692 189672 185860 189700
rect 159692 189660 159698 189672
rect 185854 189660 185860 189672
rect 185912 189660 185918 189712
rect 137186 188640 137192 188692
rect 137244 188680 137250 188692
rect 137554 188680 137560 188692
rect 137244 188652 137560 188680
rect 137244 188640 137250 188652
rect 137554 188640 137560 188652
rect 137612 188640 137618 188692
rect 132218 188368 132224 188420
rect 132276 188408 132282 188420
rect 132402 188408 132408 188420
rect 132276 188380 132408 188408
rect 132276 188368 132282 188380
rect 132402 188368 132408 188380
rect 132460 188368 132466 188420
rect 142522 188368 142528 188420
rect 142580 188408 142586 188420
rect 143258 188408 143264 188420
rect 142580 188380 143264 188408
rect 142580 188368 142586 188380
rect 143258 188368 143264 188380
rect 143316 188368 143322 188420
rect 168558 188368 168564 188420
rect 168616 188408 168622 188420
rect 168742 188408 168748 188420
rect 168616 188380 168748 188408
rect 168616 188368 168622 188380
rect 168742 188368 168748 188380
rect 168800 188368 168806 188420
rect 168466 188096 168472 188148
rect 168524 188136 168530 188148
rect 169662 188136 169668 188148
rect 168524 188108 169668 188136
rect 168524 188096 168530 188108
rect 169662 188096 169668 188108
rect 169720 188096 169726 188148
rect 135714 187688 135720 187740
rect 135772 187728 135778 187740
rect 136542 187728 136548 187740
rect 135772 187700 136548 187728
rect 135772 187688 135778 187700
rect 136542 187688 136548 187700
rect 136600 187688 136606 187740
rect 172514 187552 172520 187604
rect 172572 187592 172578 187604
rect 173342 187592 173348 187604
rect 172572 187564 173348 187592
rect 172572 187552 172578 187564
rect 173342 187552 173348 187564
rect 173400 187552 173406 187604
rect 101950 187484 101956 187536
rect 102008 187524 102014 187536
rect 135622 187524 135628 187536
rect 102008 187496 135628 187524
rect 102008 187484 102014 187496
rect 135622 187484 135628 187496
rect 135680 187484 135686 187536
rect 166166 187484 166172 187536
rect 166224 187524 166230 187536
rect 212718 187524 212724 187536
rect 166224 187496 212724 187524
rect 166224 187484 166230 187496
rect 212718 187484 212724 187496
rect 212776 187484 212782 187536
rect 100294 187416 100300 187468
rect 100352 187456 100358 187468
rect 133966 187456 133972 187468
rect 100352 187428 133972 187456
rect 100352 187416 100358 187428
rect 133966 187416 133972 187428
rect 134024 187416 134030 187468
rect 161934 187416 161940 187468
rect 161992 187456 161998 187468
rect 210418 187456 210424 187468
rect 161992 187428 210424 187456
rect 161992 187416 161998 187428
rect 210418 187416 210424 187428
rect 210476 187416 210482 187468
rect 105906 187348 105912 187400
rect 105964 187388 105970 187400
rect 139946 187388 139952 187400
rect 105964 187360 139952 187388
rect 105964 187348 105970 187360
rect 139946 187348 139952 187360
rect 140004 187348 140010 187400
rect 160462 187348 160468 187400
rect 160520 187388 160526 187400
rect 208946 187388 208952 187400
rect 160520 187360 208952 187388
rect 160520 187348 160526 187360
rect 208946 187348 208952 187360
rect 209004 187348 209010 187400
rect 100386 187280 100392 187332
rect 100444 187320 100450 187332
rect 134334 187320 134340 187332
rect 100444 187292 134340 187320
rect 100444 187280 100450 187292
rect 134334 187280 134340 187292
rect 134392 187280 134398 187332
rect 160370 187280 160376 187332
rect 160428 187320 160434 187332
rect 208854 187320 208860 187332
rect 160428 187292 208860 187320
rect 160428 187280 160434 187292
rect 208854 187280 208860 187292
rect 208912 187280 208918 187332
rect 104434 187212 104440 187264
rect 104492 187252 104498 187264
rect 138290 187252 138296 187264
rect 104492 187224 138296 187252
rect 104492 187212 104498 187224
rect 138290 187212 138296 187224
rect 138348 187212 138354 187264
rect 163866 187212 163872 187264
rect 163924 187252 163930 187264
rect 215662 187252 215668 187264
rect 163924 187224 215668 187252
rect 163924 187212 163930 187224
rect 215662 187212 215668 187224
rect 215720 187212 215726 187264
rect 98914 187144 98920 187196
rect 98972 187184 98978 187196
rect 133506 187184 133512 187196
rect 98972 187156 133512 187184
rect 98972 187144 98978 187156
rect 133506 187144 133512 187156
rect 133564 187144 133570 187196
rect 168190 187144 168196 187196
rect 168248 187184 168254 187196
rect 219710 187184 219716 187196
rect 168248 187156 219716 187184
rect 168248 187144 168254 187156
rect 219710 187144 219716 187156
rect 219768 187144 219774 187196
rect 98730 187076 98736 187128
rect 98788 187116 98794 187128
rect 133230 187116 133236 187128
rect 98788 187088 133236 187116
rect 98788 187076 98794 187088
rect 133230 187076 133236 187088
rect 133288 187076 133294 187128
rect 156322 187076 156328 187128
rect 156380 187116 156386 187128
rect 210050 187116 210056 187128
rect 156380 187088 210056 187116
rect 156380 187076 156386 187088
rect 210050 187076 210056 187088
rect 210108 187076 210114 187128
rect 106918 187008 106924 187060
rect 106976 187048 106982 187060
rect 141602 187048 141608 187060
rect 106976 187020 141608 187048
rect 106976 187008 106982 187020
rect 141602 187008 141608 187020
rect 141660 187008 141666 187060
rect 158898 187008 158904 187060
rect 158956 187048 158962 187060
rect 218238 187048 218244 187060
rect 158956 187020 218244 187048
rect 158956 187008 158962 187020
rect 218238 187008 218244 187020
rect 218296 187008 218302 187060
rect 98822 186940 98828 186992
rect 98880 186980 98886 186992
rect 145374 186980 145380 186992
rect 98880 186952 145380 186980
rect 98880 186940 98886 186952
rect 145374 186940 145380 186952
rect 145432 186940 145438 186992
rect 152366 186940 152372 186992
rect 152424 186980 152430 186992
rect 217410 186980 217416 186992
rect 152424 186952 217416 186980
rect 152424 186940 152430 186952
rect 217410 186940 217416 186952
rect 217468 186940 217474 186992
rect 134242 186464 134248 186516
rect 134300 186504 134306 186516
rect 135070 186504 135076 186516
rect 134300 186476 135076 186504
rect 134300 186464 134306 186476
rect 135070 186464 135076 186476
rect 135128 186464 135134 186516
rect 189810 165588 189816 165640
rect 189868 165628 189874 165640
rect 580166 165628 580172 165640
rect 189868 165600 580172 165628
rect 189868 165588 189874 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 164786 158652 164792 158704
rect 164844 158692 164850 158704
rect 197906 158692 197912 158704
rect 164844 158664 197912 158692
rect 164844 158652 164850 158664
rect 197906 158652 197912 158664
rect 197964 158652 197970 158704
rect 177114 158584 177120 158636
rect 177172 158624 177178 158636
rect 210602 158624 210608 158636
rect 177172 158596 210608 158624
rect 177172 158584 177178 158596
rect 210602 158584 210608 158596
rect 210660 158584 210666 158636
rect 165982 158516 165988 158568
rect 166040 158556 166046 158568
rect 201218 158556 201224 158568
rect 166040 158528 201224 158556
rect 166040 158516 166046 158528
rect 201218 158516 201224 158528
rect 201276 158516 201282 158568
rect 168742 158448 168748 158500
rect 168800 158488 168806 158500
rect 203426 158488 203432 158500
rect 168800 158460 203432 158488
rect 168800 158448 168806 158460
rect 203426 158448 203432 158460
rect 203484 158448 203490 158500
rect 168006 158380 168012 158432
rect 168064 158420 168070 158432
rect 216030 158420 216036 158432
rect 168064 158392 216036 158420
rect 168064 158380 168070 158392
rect 216030 158380 216036 158392
rect 216088 158380 216094 158432
rect 166074 158312 166080 158364
rect 166132 158352 166138 158364
rect 217502 158352 217508 158364
rect 166132 158324 217508 158352
rect 166132 158312 166138 158324
rect 217502 158312 217508 158324
rect 217560 158312 217566 158364
rect 152366 158244 152372 158296
rect 152424 158284 152430 158296
rect 204714 158284 204720 158296
rect 152424 158256 204720 158284
rect 152424 158244 152430 158256
rect 204714 158244 204720 158256
rect 204772 158244 204778 158296
rect 164694 158176 164700 158228
rect 164752 158216 164758 158228
rect 219894 158216 219900 158228
rect 164752 158188 219900 158216
rect 164752 158176 164758 158188
rect 219894 158176 219900 158188
rect 219952 158176 219958 158228
rect 164602 158108 164608 158160
rect 164660 158148 164666 158160
rect 219986 158148 219992 158160
rect 164660 158120 219992 158148
rect 164660 158108 164666 158120
rect 219986 158108 219992 158120
rect 220044 158108 220050 158160
rect 163130 158040 163136 158092
rect 163188 158080 163194 158092
rect 219802 158080 219808 158092
rect 163188 158052 219808 158080
rect 163188 158040 163194 158052
rect 219802 158040 219808 158052
rect 219860 158040 219866 158092
rect 152274 157972 152280 158024
rect 152332 158012 152338 158024
rect 218054 158012 218060 158024
rect 152332 157984 218060 158012
rect 152332 157972 152338 157984
rect 218054 157972 218060 157984
rect 218112 157972 218118 158024
rect 168834 157904 168840 157956
rect 168892 157944 168898 157956
rect 197998 157944 198004 157956
rect 168892 157916 198004 157944
rect 168892 157904 168898 157916
rect 197998 157904 198004 157916
rect 198056 157904 198062 157956
rect 168926 157836 168932 157888
rect 168984 157876 168990 157888
rect 196618 157876 196624 157888
rect 168984 157848 196624 157876
rect 168984 157836 168990 157848
rect 196618 157836 196624 157848
rect 196676 157836 196682 157888
rect 177206 157768 177212 157820
rect 177264 157808 177270 157820
rect 203334 157808 203340 157820
rect 177264 157780 203340 157808
rect 177264 157768 177270 157780
rect 203334 157768 203340 157780
rect 203392 157768 203398 157820
rect 163038 155864 163044 155916
rect 163096 155904 163102 155916
rect 184382 155904 184388 155916
rect 163096 155876 184388 155904
rect 163096 155864 163102 155876
rect 184382 155864 184388 155876
rect 184440 155864 184446 155916
rect 161842 155796 161848 155848
rect 161900 155836 161906 155848
rect 184290 155836 184296 155848
rect 161900 155808 184296 155836
rect 161900 155796 161906 155808
rect 184290 155796 184296 155808
rect 184348 155796 184354 155848
rect 162946 155728 162952 155780
rect 163004 155768 163010 155780
rect 186038 155768 186044 155780
rect 163004 155740 186044 155768
rect 163004 155728 163010 155740
rect 186038 155728 186044 155740
rect 186096 155728 186102 155780
rect 164326 155660 164332 155712
rect 164384 155700 164390 155712
rect 188522 155700 188528 155712
rect 164384 155672 188528 155700
rect 164384 155660 164390 155672
rect 188522 155660 188528 155672
rect 188580 155660 188586 155712
rect 171502 155592 171508 155644
rect 171560 155632 171566 155644
rect 200574 155632 200580 155644
rect 171560 155604 200580 155632
rect 171560 155592 171566 155604
rect 200574 155592 200580 155604
rect 200632 155592 200638 155644
rect 158806 155524 158812 155576
rect 158864 155564 158870 155576
rect 188430 155564 188436 155576
rect 158864 155536 188436 155564
rect 158864 155524 158870 155536
rect 188430 155524 188436 155536
rect 188488 155524 188494 155576
rect 157702 155456 157708 155508
rect 157760 155496 157766 155508
rect 188614 155496 188620 155508
rect 157760 155468 188620 155496
rect 157760 155456 157766 155468
rect 188614 155456 188620 155468
rect 188672 155456 188678 155508
rect 165890 155388 165896 155440
rect 165948 155428 165954 155440
rect 200666 155428 200672 155440
rect 165948 155400 200672 155428
rect 165948 155388 165954 155400
rect 200666 155388 200672 155400
rect 200724 155388 200730 155440
rect 165798 155320 165804 155372
rect 165856 155360 165862 155372
rect 200758 155360 200764 155372
rect 165856 155332 200764 155360
rect 165856 155320 165862 155332
rect 200758 155320 200764 155332
rect 200816 155320 200822 155372
rect 165706 155252 165712 155304
rect 165764 155292 165770 155304
rect 211890 155292 211896 155304
rect 165764 155264 211896 155292
rect 165764 155252 165770 155264
rect 211890 155252 211896 155264
rect 211948 155252 211954 155304
rect 164510 155184 164516 155236
rect 164568 155224 164574 155236
rect 212994 155224 213000 155236
rect 164568 155196 213000 155224
rect 164568 155184 164574 155196
rect 212994 155184 213000 155196
rect 213052 155184 213058 155236
rect 164418 155116 164424 155168
rect 164476 155156 164482 155168
rect 184198 155156 184204 155168
rect 164476 155128 184204 155156
rect 164476 155116 164482 155128
rect 184198 155116 184204 155128
rect 184256 155116 184262 155168
rect 119338 154164 119344 154216
rect 119396 154204 119402 154216
rect 133966 154204 133972 154216
rect 119396 154176 133972 154204
rect 119396 154164 119402 154176
rect 133966 154164 133972 154176
rect 134024 154164 134030 154216
rect 96246 154096 96252 154148
rect 96304 154136 96310 154148
rect 134518 154136 134524 154148
rect 96304 154108 134524 154136
rect 96304 154096 96310 154108
rect 134518 154096 134524 154108
rect 134576 154096 134582 154148
rect 97166 154028 97172 154080
rect 97224 154068 97230 154080
rect 140222 154068 140228 154080
rect 97224 154040 140228 154068
rect 97224 154028 97230 154040
rect 140222 154028 140228 154040
rect 140280 154028 140286 154080
rect 96154 153960 96160 154012
rect 96212 154000 96218 154012
rect 140406 154000 140412 154012
rect 96212 153972 140412 154000
rect 96212 153960 96218 153972
rect 140406 153960 140412 153972
rect 140464 153960 140470 154012
rect 165706 153960 165712 154012
rect 165764 154000 165770 154012
rect 203242 154000 203248 154012
rect 165764 153972 203248 154000
rect 165764 153960 165770 153972
rect 203242 153960 203248 153972
rect 203300 153960 203306 154012
rect 96982 153892 96988 153944
rect 97040 153932 97046 153944
rect 145282 153932 145288 153944
rect 97040 153904 145288 153932
rect 97040 153892 97046 153904
rect 145282 153892 145288 153904
rect 145340 153892 145346 153944
rect 162946 153892 162952 153944
rect 163004 153932 163010 153944
rect 204622 153932 204628 153944
rect 163004 153904 204628 153932
rect 163004 153892 163010 153904
rect 204622 153892 204628 153904
rect 204680 153892 204686 153944
rect 120902 153824 120908 153876
rect 120960 153864 120966 153876
rect 170122 153864 170128 153876
rect 120960 153836 170128 153864
rect 120960 153824 120966 153836
rect 170122 153824 170128 153836
rect 170180 153824 170186 153876
rect 173710 153824 173716 153876
rect 173768 153864 173774 153876
rect 214742 153864 214748 153876
rect 173768 153836 214748 153864
rect 173768 153824 173774 153836
rect 214742 153824 214748 153836
rect 214800 153824 214806 153876
rect 95878 153212 95884 153264
rect 95936 153252 95942 153264
rect 184934 153252 184940 153264
rect 95936 153224 184940 153252
rect 95936 153212 95942 153224
rect 184934 153212 184940 153224
rect 184992 153252 184998 153264
rect 192570 153252 192576 153264
rect 184992 153224 192576 153252
rect 184992 153212 184998 153224
rect 192570 153212 192576 153224
rect 192628 153212 192634 153264
rect 158530 153144 158536 153196
rect 158588 153184 158594 153196
rect 187326 153184 187332 153196
rect 158588 153156 187332 153184
rect 158588 153144 158594 153156
rect 187326 153144 187332 153156
rect 187384 153144 187390 153196
rect 156230 153076 156236 153128
rect 156288 153116 156294 153128
rect 187142 153116 187148 153128
rect 156288 153088 187148 153116
rect 156288 153076 156294 153088
rect 187142 153076 187148 153088
rect 187200 153076 187206 153128
rect 157610 153008 157616 153060
rect 157668 153048 157674 153060
rect 188706 153048 188712 153060
rect 157668 153020 188712 153048
rect 157668 153008 157674 153020
rect 188706 153008 188712 153020
rect 188764 153008 188770 153060
rect 160186 152940 160192 152992
rect 160244 152980 160250 152992
rect 184658 152980 184664 152992
rect 160244 152952 184664 152980
rect 160244 152940 160250 152952
rect 184658 152940 184664 152952
rect 184716 152940 184722 152992
rect 186958 152940 186964 152992
rect 187016 152980 187022 152992
rect 218422 152980 218428 152992
rect 187016 152952 218428 152980
rect 187016 152940 187022 152952
rect 218422 152940 218428 152952
rect 218480 152940 218486 152992
rect 175550 152872 175556 152924
rect 175608 152912 175614 152924
rect 207934 152912 207940 152924
rect 175608 152884 207940 152912
rect 175608 152872 175614 152884
rect 207934 152872 207940 152884
rect 207992 152872 207998 152924
rect 176746 152804 176752 152856
rect 176804 152844 176810 152856
rect 209130 152844 209136 152856
rect 176804 152816 209136 152844
rect 176804 152804 176810 152816
rect 209130 152804 209136 152816
rect 209188 152804 209194 152856
rect 176654 152736 176660 152788
rect 176712 152776 176718 152788
rect 209038 152776 209044 152788
rect 176712 152748 209044 152776
rect 176712 152736 176718 152748
rect 209038 152736 209044 152748
rect 209096 152736 209102 152788
rect 157518 152668 157524 152720
rect 157576 152708 157582 152720
rect 191374 152708 191380 152720
rect 157576 152680 191380 152708
rect 157576 152668 157582 152680
rect 191374 152668 191380 152680
rect 191432 152668 191438 152720
rect 160278 152600 160284 152652
rect 160336 152640 160342 152652
rect 209222 152640 209228 152652
rect 160336 152612 209228 152640
rect 160336 152600 160342 152612
rect 209222 152600 209228 152612
rect 209280 152600 209286 152652
rect 158714 152532 158720 152584
rect 158772 152572 158778 152584
rect 218330 152572 218336 152584
rect 158772 152544 218336 152572
rect 158772 152532 158778 152544
rect 218330 152532 218336 152544
rect 218388 152532 218394 152584
rect 111150 152464 111156 152516
rect 111208 152504 111214 152516
rect 142890 152504 142896 152516
rect 111208 152476 142896 152504
rect 111208 152464 111214 152476
rect 142890 152464 142896 152476
rect 142948 152464 142954 152516
rect 154942 152464 154948 152516
rect 155000 152504 155006 152516
rect 218606 152504 218612 152516
rect 155000 152476 218612 152504
rect 155000 152464 155006 152476
rect 218606 152464 218612 152476
rect 218664 152464 218670 152516
rect 157426 152396 157432 152448
rect 157484 152436 157490 152448
rect 187234 152436 187240 152448
rect 157484 152408 187240 152436
rect 157484 152396 157490 152408
rect 187234 152396 187240 152408
rect 187292 152396 187298 152448
rect 183462 152328 183468 152380
rect 183520 152368 183526 152380
rect 207658 152368 207664 152380
rect 183520 152340 207664 152368
rect 183520 152328 183526 152340
rect 207658 152328 207664 152340
rect 207716 152328 207722 152380
rect 187970 151784 187976 151836
rect 188028 151824 188034 151836
rect 580074 151824 580080 151836
rect 188028 151796 580080 151824
rect 188028 151784 188034 151796
rect 580074 151784 580080 151796
rect 580132 151784 580138 151836
rect 114922 151716 114928 151768
rect 114980 151756 114986 151768
rect 140958 151756 140964 151768
rect 114980 151728 140964 151756
rect 114980 151716 114986 151728
rect 140958 151716 140964 151728
rect 141016 151716 141022 151768
rect 101398 151648 101404 151700
rect 101456 151688 101462 151700
rect 134242 151688 134248 151700
rect 101456 151660 134248 151688
rect 101456 151648 101462 151660
rect 134242 151648 134248 151660
rect 134300 151648 134306 151700
rect 102778 151580 102784 151632
rect 102836 151620 102842 151632
rect 135806 151620 135812 151632
rect 102836 151592 135812 151620
rect 102836 151580 102842 151592
rect 135806 151580 135812 151592
rect 135864 151580 135870 151632
rect 98638 151512 98644 151564
rect 98696 151552 98702 151564
rect 133046 151552 133052 151564
rect 98696 151524 133052 151552
rect 98696 151512 98702 151524
rect 133046 151512 133052 151524
rect 133104 151512 133110 151564
rect 102962 151444 102968 151496
rect 103020 151484 103026 151496
rect 137370 151484 137376 151496
rect 103020 151456 137376 151484
rect 103020 151444 103026 151456
rect 137370 151444 137376 151456
rect 137428 151444 137434 151496
rect 100018 151376 100024 151428
rect 100076 151416 100082 151428
rect 134334 151416 134340 151428
rect 100076 151388 134340 151416
rect 100076 151376 100082 151388
rect 134334 151376 134340 151388
rect 134392 151376 134398 151428
rect 174538 151376 174544 151428
rect 174596 151416 174602 151428
rect 199470 151416 199476 151428
rect 174596 151388 199476 151416
rect 174596 151376 174602 151388
rect 199470 151376 199476 151388
rect 199528 151376 199534 151428
rect 100110 151308 100116 151360
rect 100168 151348 100174 151360
rect 134058 151348 134064 151360
rect 100168 151320 134064 151348
rect 100168 151308 100174 151320
rect 134058 151308 134064 151320
rect 134116 151308 134122 151360
rect 171962 151308 171968 151360
rect 172020 151348 172026 151360
rect 206002 151348 206008 151360
rect 172020 151320 206008 151348
rect 172020 151308 172026 151320
rect 206002 151308 206008 151320
rect 206060 151308 206066 151360
rect 101490 151240 101496 151292
rect 101548 151280 101554 151292
rect 136082 151280 136088 151292
rect 101548 151252 136088 151280
rect 101548 151240 101554 151252
rect 136082 151240 136088 151252
rect 136140 151240 136146 151292
rect 168650 151240 168656 151292
rect 168708 151280 168714 151292
rect 203518 151280 203524 151292
rect 168708 151252 203524 151280
rect 168708 151240 168714 151252
rect 203518 151240 203524 151252
rect 203576 151240 203582 151292
rect 98546 151172 98552 151224
rect 98604 151212 98610 151224
rect 133138 151212 133144 151224
rect 98604 151184 133144 151212
rect 98604 151172 98610 151184
rect 133138 151172 133144 151184
rect 133196 151172 133202 151224
rect 167270 151172 167276 151224
rect 167328 151212 167334 151224
rect 206094 151212 206100 151224
rect 167328 151184 206100 151212
rect 167328 151172 167334 151184
rect 206094 151172 206100 151184
rect 206152 151172 206158 151224
rect 101306 151104 101312 151156
rect 101364 151144 101370 151156
rect 135530 151144 135536 151156
rect 101364 151116 135536 151144
rect 101364 151104 101370 151116
rect 135530 151104 135536 151116
rect 135588 151104 135594 151156
rect 154942 151104 154948 151156
rect 155000 151144 155006 151156
rect 207566 151144 207572 151156
rect 155000 151116 207572 151144
rect 155000 151104 155006 151116
rect 207566 151104 207572 151116
rect 207624 151104 207630 151156
rect 96062 151036 96068 151088
rect 96120 151076 96126 151088
rect 139302 151076 139308 151088
rect 96120 151048 139308 151076
rect 96120 151036 96126 151048
rect 139302 151036 139308 151048
rect 139360 151036 139366 151088
rect 153562 151036 153568 151088
rect 153620 151076 153626 151088
rect 207106 151076 207112 151088
rect 153620 151048 207112 151076
rect 153620 151036 153626 151048
rect 207106 151036 207112 151048
rect 207164 151036 207170 151088
rect 118970 150968 118976 151020
rect 119028 151008 119034 151020
rect 144914 151008 144920 151020
rect 119028 150980 144920 151008
rect 119028 150968 119034 150980
rect 144914 150968 144920 150980
rect 144972 150968 144978 151020
rect 124030 150900 124036 150952
rect 124088 150940 124094 150952
rect 141878 150940 141884 150952
rect 124088 150912 141884 150940
rect 124088 150900 124094 150912
rect 141878 150900 141884 150912
rect 141936 150900 141942 150952
rect 125042 150424 125048 150476
rect 125100 150464 125106 150476
rect 580534 150464 580540 150476
rect 125100 150436 580540 150464
rect 125100 150424 125106 150436
rect 580534 150424 580540 150436
rect 580592 150424 580598 150476
rect 182082 150356 182088 150408
rect 182140 150396 182146 150408
rect 195054 150396 195060 150408
rect 182140 150368 195060 150396
rect 182140 150356 182146 150368
rect 195054 150356 195060 150368
rect 195112 150356 195118 150408
rect 171870 150288 171876 150340
rect 171928 150328 171934 150340
rect 191282 150328 191288 150340
rect 171928 150300 191288 150328
rect 171928 150288 171934 150300
rect 191282 150288 191288 150300
rect 191340 150288 191346 150340
rect 175366 150220 175372 150272
rect 175424 150260 175430 150272
rect 204898 150260 204904 150272
rect 175424 150232 204904 150260
rect 175424 150220 175430 150232
rect 204898 150220 204904 150232
rect 204956 150220 204962 150272
rect 172882 150152 172888 150204
rect 172940 150192 172946 150204
rect 206186 150192 206192 150204
rect 172940 150164 206192 150192
rect 172940 150152 172946 150164
rect 206186 150152 206192 150164
rect 206244 150152 206250 150204
rect 174170 150084 174176 150136
rect 174228 150124 174234 150136
rect 207566 150124 207572 150136
rect 174228 150096 207572 150124
rect 174228 150084 174234 150096
rect 207566 150084 207572 150096
rect 207624 150084 207630 150136
rect 172698 150016 172704 150068
rect 172756 150056 172762 150068
rect 206278 150056 206284 150068
rect 172756 150028 206284 150056
rect 172756 150016 172762 150028
rect 206278 150016 206284 150028
rect 206336 150016 206342 150068
rect 173894 149948 173900 150000
rect 173952 149988 173958 150000
rect 207750 149988 207756 150000
rect 173952 149960 207756 149988
rect 173952 149948 173958 149960
rect 207750 149948 207756 149960
rect 207808 149948 207814 150000
rect 173986 149880 173992 149932
rect 174044 149920 174050 149932
rect 207658 149920 207664 149932
rect 174044 149892 207664 149920
rect 174044 149880 174050 149892
rect 207658 149880 207664 149892
rect 207716 149880 207722 149932
rect 171318 149812 171324 149864
rect 171376 149852 171382 149864
rect 204990 149852 204996 149864
rect 171376 149824 204996 149852
rect 171376 149812 171382 149824
rect 204990 149812 204996 149824
rect 205048 149812 205054 149864
rect 175182 149744 175188 149796
rect 175240 149784 175246 149796
rect 207842 149784 207848 149796
rect 175240 149756 207848 149784
rect 175240 149744 175246 149756
rect 207842 149744 207848 149756
rect 207900 149744 207906 149796
rect 99834 149676 99840 149728
rect 99892 149716 99898 149728
rect 148042 149716 148048 149728
rect 99892 149688 148048 149716
rect 99892 149676 99898 149688
rect 148042 149676 148048 149688
rect 148100 149676 148106 149728
rect 171410 149676 171416 149728
rect 171468 149716 171474 149728
rect 206094 149716 206100 149728
rect 171468 149688 206100 149716
rect 171468 149676 171474 149688
rect 206094 149676 206100 149688
rect 206152 149676 206158 149728
rect 3142 149132 3148 149184
rect 3200 149172 3206 149184
rect 180886 149172 180892 149184
rect 3200 149144 180892 149172
rect 3200 149132 3206 149144
rect 180886 149132 180892 149144
rect 180944 149172 180950 149184
rect 182082 149172 182088 149184
rect 180944 149144 182088 149172
rect 180944 149132 180950 149144
rect 182082 149132 182088 149144
rect 182140 149132 182146 149184
rect 125686 149064 125692 149116
rect 125744 149104 125750 149116
rect 126514 149104 126520 149116
rect 125744 149076 126520 149104
rect 125744 149064 125750 149076
rect 126514 149064 126520 149076
rect 126572 149104 126578 149116
rect 580626 149104 580632 149116
rect 126572 149076 580632 149104
rect 126572 149064 126578 149076
rect 580626 149064 580632 149076
rect 580684 149064 580690 149116
rect 118878 148996 118884 149048
rect 118936 149036 118942 149048
rect 147030 149036 147036 149048
rect 118936 149008 147036 149036
rect 118936 148996 118942 149008
rect 147030 148996 147036 149008
rect 147088 148996 147094 149048
rect 171042 148996 171048 149048
rect 171100 149036 171106 149048
rect 195054 149036 195060 149048
rect 171100 149008 195060 149036
rect 171100 148996 171106 149008
rect 195054 148996 195060 149008
rect 195112 148996 195118 149048
rect 104158 148928 104164 148980
rect 104216 148968 104222 148980
rect 131942 148968 131948 148980
rect 104216 148940 131948 148968
rect 104216 148928 104222 148940
rect 131942 148928 131948 148940
rect 132000 148928 132006 148980
rect 161750 148928 161756 148980
rect 161808 148968 161814 148980
rect 188798 148968 188804 148980
rect 161808 148940 188804 148968
rect 161808 148928 161814 148940
rect 188798 148928 188804 148940
rect 188856 148928 188862 148980
rect 110782 148860 110788 148912
rect 110840 148900 110846 148912
rect 142522 148900 142528 148912
rect 110840 148872 142528 148900
rect 110840 148860 110846 148872
rect 142522 148860 142528 148872
rect 142580 148860 142586 148912
rect 162762 148860 162768 148912
rect 162820 148900 162826 148912
rect 198366 148900 198372 148912
rect 162820 148872 198372 148900
rect 162820 148860 162826 148872
rect 198366 148860 198372 148872
rect 198424 148860 198430 148912
rect 122466 148792 122472 148844
rect 122524 148832 122530 148844
rect 153470 148832 153476 148844
rect 122524 148804 153476 148832
rect 122524 148792 122530 148804
rect 153470 148792 153476 148804
rect 153528 148792 153534 148844
rect 161014 148792 161020 148844
rect 161072 148832 161078 148844
rect 195606 148832 195612 148844
rect 161072 148804 195612 148832
rect 161072 148792 161078 148804
rect 195606 148792 195612 148804
rect 195664 148792 195670 148844
rect 111058 148724 111064 148776
rect 111116 148764 111122 148776
rect 142614 148764 142620 148776
rect 111116 148736 142620 148764
rect 111116 148724 111122 148736
rect 142614 148724 142620 148736
rect 142672 148724 142678 148776
rect 161290 148724 161296 148776
rect 161348 148764 161354 148776
rect 196894 148764 196900 148776
rect 161348 148736 196900 148764
rect 161348 148724 161354 148736
rect 196894 148724 196900 148736
rect 196952 148724 196958 148776
rect 98454 148656 98460 148708
rect 98512 148696 98518 148708
rect 130654 148696 130660 148708
rect 98512 148668 130660 148696
rect 98512 148656 98518 148668
rect 130654 148656 130660 148668
rect 130712 148656 130718 148708
rect 164234 148656 164240 148708
rect 164292 148696 164298 148708
rect 199746 148696 199752 148708
rect 164292 148668 199752 148696
rect 164292 148656 164298 148668
rect 199746 148656 199752 148668
rect 199804 148656 199810 148708
rect 118786 148588 118792 148640
rect 118844 148628 118850 148640
rect 152182 148628 152188 148640
rect 118844 148600 152188 148628
rect 118844 148588 118850 148600
rect 152182 148588 152188 148600
rect 152240 148588 152246 148640
rect 168282 148588 168288 148640
rect 168340 148628 168346 148640
rect 202046 148628 202052 148640
rect 168340 148600 202052 148628
rect 168340 148588 168346 148600
rect 202046 148588 202052 148600
rect 202104 148588 202110 148640
rect 99926 148520 99932 148572
rect 99984 148560 99990 148572
rect 132310 148560 132316 148572
rect 99984 148532 132316 148560
rect 99984 148520 99990 148532
rect 132310 148520 132316 148532
rect 132368 148520 132374 148572
rect 169662 148520 169668 148572
rect 169720 148560 169726 148572
rect 203702 148560 203708 148572
rect 169720 148532 203708 148560
rect 169720 148520 169726 148532
rect 203702 148520 203708 148532
rect 203760 148520 203766 148572
rect 114830 148452 114836 148504
rect 114888 148492 114894 148504
rect 149330 148492 149336 148504
rect 114888 148464 149336 148492
rect 114888 148452 114894 148464
rect 149330 148452 149336 148464
rect 149388 148452 149394 148504
rect 160002 148452 160008 148504
rect 160060 148492 160066 148504
rect 195146 148492 195152 148504
rect 160060 148464 195152 148492
rect 160060 148452 160066 148464
rect 195146 148452 195152 148464
rect 195204 148452 195210 148504
rect 97074 148384 97080 148436
rect 97132 148424 97138 148436
rect 152090 148424 152096 148436
rect 97132 148396 152096 148424
rect 97132 148384 97138 148396
rect 152090 148384 152096 148396
rect 152148 148384 152154 148436
rect 165614 148384 165620 148436
rect 165672 148424 165678 148436
rect 200850 148424 200856 148436
rect 165672 148396 200856 148424
rect 165672 148384 165678 148396
rect 200850 148384 200856 148396
rect 200908 148384 200914 148436
rect 112346 148316 112352 148368
rect 112404 148356 112410 148368
rect 128906 148356 128912 148368
rect 112404 148328 128912 148356
rect 112404 148316 112410 148328
rect 128906 148316 128912 148328
rect 128964 148356 128970 148368
rect 187970 148356 187976 148368
rect 128964 148328 187976 148356
rect 128964 148316 128970 148328
rect 187970 148316 187976 148328
rect 188028 148316 188034 148368
rect 120902 148248 120908 148300
rect 120960 148288 120966 148300
rect 147950 148288 147956 148300
rect 120960 148260 147956 148288
rect 120960 148248 120966 148260
rect 147950 148248 147956 148260
rect 148008 148248 148014 148300
rect 177666 148248 177672 148300
rect 177724 148288 177730 148300
rect 199654 148288 199660 148300
rect 177724 148260 199660 148288
rect 177724 148248 177730 148260
rect 199654 148248 199660 148260
rect 199712 148248 199718 148300
rect 106734 148180 106740 148232
rect 106792 148220 106798 148232
rect 131850 148220 131856 148232
rect 106792 148192 131856 148220
rect 106792 148180 106798 148192
rect 131850 148180 131856 148192
rect 131908 148180 131914 148232
rect 179598 147568 179604 147620
rect 179656 147608 179662 147620
rect 196434 147608 196440 147620
rect 179656 147580 196440 147608
rect 179656 147568 179662 147580
rect 196434 147568 196440 147580
rect 196492 147568 196498 147620
rect 179782 147500 179788 147552
rect 179840 147540 179846 147552
rect 199194 147540 199200 147552
rect 179840 147512 199200 147540
rect 179840 147500 179846 147512
rect 199194 147500 199200 147512
rect 199252 147500 199258 147552
rect 178586 147432 178592 147484
rect 178644 147472 178650 147484
rect 199286 147472 199292 147484
rect 178644 147444 199292 147472
rect 178644 147432 178650 147444
rect 199286 147432 199292 147444
rect 199344 147432 199350 147484
rect 176654 147364 176660 147416
rect 176712 147404 176718 147416
rect 197814 147404 197820 147416
rect 176712 147376 197820 147404
rect 176712 147364 176718 147376
rect 197814 147364 197820 147376
rect 197872 147364 197878 147416
rect 109586 147296 109592 147348
rect 109644 147336 109650 147348
rect 138566 147336 138572 147348
rect 109644 147308 138572 147336
rect 109644 147296 109650 147308
rect 138566 147296 138572 147308
rect 138624 147296 138630 147348
rect 170030 147296 170036 147348
rect 170088 147336 170094 147348
rect 195698 147336 195704 147348
rect 170088 147308 195704 147336
rect 170088 147296 170094 147308
rect 195698 147296 195704 147308
rect 195756 147296 195762 147348
rect 105354 147228 105360 147280
rect 105412 147268 105418 147280
rect 137186 147268 137192 147280
rect 105412 147240 137192 147268
rect 105412 147228 105418 147240
rect 137186 147228 137192 147240
rect 137244 147228 137250 147280
rect 169846 147228 169852 147280
rect 169904 147268 169910 147280
rect 199286 147268 199292 147280
rect 169904 147240 199292 147268
rect 169904 147228 169910 147240
rect 199286 147228 199292 147240
rect 199344 147228 199350 147280
rect 110690 147160 110696 147212
rect 110748 147200 110754 147212
rect 143994 147200 144000 147212
rect 110748 147172 144000 147200
rect 110748 147160 110754 147172
rect 143994 147160 144000 147172
rect 144052 147160 144058 147212
rect 157334 147160 157340 147212
rect 157392 147200 157398 147212
rect 182726 147200 182732 147212
rect 157392 147172 182732 147200
rect 157392 147160 157398 147172
rect 182726 147160 182732 147172
rect 182784 147160 182790 147212
rect 182910 147160 182916 147212
rect 182968 147200 182974 147212
rect 183186 147200 183192 147212
rect 182968 147172 183192 147200
rect 182968 147160 182974 147172
rect 183186 147160 183192 147172
rect 183244 147160 183250 147212
rect 102870 147092 102876 147144
rect 102928 147132 102934 147144
rect 135714 147132 135720 147144
rect 102928 147104 135720 147132
rect 102928 147092 102934 147104
rect 135714 147092 135720 147104
rect 135772 147092 135778 147144
rect 172514 147092 172520 147144
rect 172572 147132 172578 147144
rect 206370 147132 206376 147144
rect 172572 147104 182772 147132
rect 172572 147092 172578 147104
rect 104066 147024 104072 147076
rect 104124 147064 104130 147076
rect 137278 147064 137284 147076
rect 104124 147036 137284 147064
rect 104124 147024 104130 147036
rect 137278 147024 137284 147036
rect 137336 147024 137342 147076
rect 156138 147024 156144 147076
rect 156196 147064 156202 147076
rect 182634 147064 182640 147076
rect 156196 147036 182640 147064
rect 156196 147024 156202 147036
rect 182634 147024 182640 147036
rect 182692 147024 182698 147076
rect 182744 147064 182772 147104
rect 182928 147104 206376 147132
rect 182928 147064 182956 147104
rect 206370 147092 206376 147104
rect 206428 147092 206434 147144
rect 182744 147036 182956 147064
rect 109402 146956 109408 147008
rect 109460 146996 109466 147008
rect 143626 146996 143632 147008
rect 109460 146968 143632 146996
rect 109460 146956 109466 146968
rect 143626 146956 143632 146968
rect 143684 146956 143690 147008
rect 171134 146956 171140 147008
rect 171192 146996 171198 147008
rect 205082 146996 205088 147008
rect 171192 146968 205088 146996
rect 171192 146956 171198 146968
rect 205082 146956 205088 146968
rect 205140 146956 205146 147008
rect 105446 146888 105452 146940
rect 105504 146928 105510 146940
rect 140130 146928 140136 146940
rect 105504 146900 140136 146928
rect 105504 146888 105510 146900
rect 140130 146888 140136 146900
rect 140188 146888 140194 146940
rect 161382 146888 161388 146940
rect 161440 146928 161446 146940
rect 197906 146928 197912 146940
rect 161440 146900 197912 146928
rect 161440 146888 161446 146900
rect 197906 146888 197912 146900
rect 197964 146888 197970 146940
rect 179506 146820 179512 146872
rect 179564 146860 179570 146872
rect 197354 146860 197360 146872
rect 179564 146832 197360 146860
rect 179564 146820 179570 146832
rect 197354 146820 197360 146832
rect 197412 146820 197418 146872
rect 181530 146752 181536 146804
rect 181588 146792 181594 146804
rect 190086 146792 190092 146804
rect 181588 146764 190092 146792
rect 181588 146752 181594 146764
rect 190086 146752 190092 146764
rect 190144 146752 190150 146804
rect 182726 146684 182732 146736
rect 182784 146724 182790 146736
rect 189718 146724 189724 146736
rect 182784 146696 189724 146724
rect 182784 146684 182790 146696
rect 189718 146684 189724 146696
rect 189776 146684 189782 146736
rect 182634 146616 182640 146668
rect 182692 146656 182698 146668
rect 189994 146656 190000 146668
rect 182692 146628 190000 146656
rect 182692 146616 182698 146628
rect 189994 146616 190000 146628
rect 190052 146616 190058 146668
rect 113818 146208 113824 146260
rect 113876 146248 113882 146260
rect 129734 146248 129740 146260
rect 113876 146220 129740 146248
rect 113876 146208 113882 146220
rect 129734 146208 129740 146220
rect 129792 146208 129798 146260
rect 180150 146208 180156 146260
rect 180208 146248 180214 146260
rect 193582 146248 193588 146260
rect 180208 146220 193588 146248
rect 180208 146208 180214 146220
rect 193582 146208 193588 146220
rect 193640 146208 193646 146260
rect 112622 146140 112628 146192
rect 112680 146180 112686 146192
rect 130010 146180 130016 146192
rect 112680 146152 130016 146180
rect 112680 146140 112686 146152
rect 130010 146140 130016 146152
rect 130068 146140 130074 146192
rect 178126 146140 178132 146192
rect 178184 146180 178190 146192
rect 193950 146180 193956 146192
rect 178184 146152 193956 146180
rect 178184 146140 178190 146152
rect 193950 146140 193956 146152
rect 194008 146140 194014 146192
rect 110966 146072 110972 146124
rect 111024 146112 111030 146124
rect 132218 146112 132224 146124
rect 111024 146084 132224 146112
rect 111024 146072 111030 146084
rect 132218 146072 132224 146084
rect 132276 146072 132282 146124
rect 178034 146072 178040 146124
rect 178092 146112 178098 146124
rect 194962 146112 194968 146124
rect 178092 146084 194968 146112
rect 178092 146072 178098 146084
rect 194962 146072 194968 146084
rect 195020 146072 195026 146124
rect 119890 146004 119896 146056
rect 119948 146044 119954 146056
rect 149238 146044 149244 146056
rect 119948 146016 149244 146044
rect 119948 146004 119954 146016
rect 149238 146004 149244 146016
rect 149296 146004 149302 146056
rect 167914 146004 167920 146056
rect 167972 146044 167978 146056
rect 194226 146044 194232 146056
rect 167972 146016 194232 146044
rect 167972 146004 167978 146016
rect 194226 146004 194232 146016
rect 194284 146004 194290 146056
rect 111426 145936 111432 145988
rect 111484 145976 111490 145988
rect 142154 145976 142160 145988
rect 111484 145948 142160 145976
rect 111484 145936 111490 145948
rect 142154 145936 142160 145948
rect 142212 145936 142218 145988
rect 165522 145936 165528 145988
rect 165580 145976 165586 145988
rect 192570 145976 192576 145988
rect 165580 145948 192576 145976
rect 165580 145936 165586 145948
rect 192570 145936 192576 145948
rect 192628 145936 192634 145988
rect 116394 145868 116400 145920
rect 116452 145908 116458 145920
rect 149054 145908 149060 145920
rect 116452 145880 149060 145908
rect 116452 145868 116458 145880
rect 149054 145868 149060 145880
rect 149112 145868 149118 145920
rect 161658 145868 161664 145920
rect 161716 145908 161722 145920
rect 196986 145908 196992 145920
rect 161716 145880 196992 145908
rect 161716 145868 161722 145880
rect 196986 145868 196992 145880
rect 197044 145868 197050 145920
rect 116210 145800 116216 145852
rect 116268 145840 116274 145852
rect 149698 145840 149704 145852
rect 116268 145812 149704 145840
rect 116268 145800 116274 145812
rect 149698 145800 149704 145812
rect 149756 145800 149762 145852
rect 157610 145800 157616 145852
rect 157668 145840 157674 145852
rect 192202 145840 192208 145852
rect 157668 145812 192208 145840
rect 157668 145800 157674 145812
rect 192202 145800 192208 145812
rect 192260 145800 192266 145852
rect 117774 145732 117780 145784
rect 117832 145772 117838 145784
rect 151814 145772 151820 145784
rect 117832 145744 151820 145772
rect 117832 145732 117838 145744
rect 151814 145732 151820 145744
rect 151872 145732 151878 145784
rect 161566 145732 161572 145784
rect 161624 145772 161630 145784
rect 197078 145772 197084 145784
rect 161624 145744 197084 145772
rect 161624 145732 161630 145744
rect 197078 145732 197084 145744
rect 197136 145732 197142 145784
rect 116302 145664 116308 145716
rect 116360 145704 116366 145716
rect 150710 145704 150716 145716
rect 116360 145676 150716 145704
rect 116360 145664 116366 145676
rect 150710 145664 150716 145676
rect 150768 145664 150774 145716
rect 157242 145664 157248 145716
rect 157300 145704 157306 145716
rect 192202 145704 192208 145716
rect 157300 145676 192208 145704
rect 157300 145664 157306 145676
rect 192202 145664 192208 145676
rect 192260 145664 192266 145716
rect 113818 145596 113824 145648
rect 113876 145636 113882 145648
rect 148410 145636 148416 145648
rect 113876 145608 148416 145636
rect 113876 145596 113882 145608
rect 148410 145596 148416 145608
rect 148468 145596 148474 145648
rect 150342 145596 150348 145648
rect 150400 145636 150406 145648
rect 190178 145636 190184 145648
rect 150400 145608 190184 145636
rect 150400 145596 150406 145608
rect 190178 145596 190184 145608
rect 190236 145596 190242 145648
rect 3510 145528 3516 145580
rect 3568 145568 3574 145580
rect 3568 145540 161474 145568
rect 3568 145528 3574 145540
rect 116486 145460 116492 145512
rect 116544 145500 116550 145512
rect 130102 145500 130108 145512
rect 116544 145472 130108 145500
rect 116544 145460 116550 145472
rect 130102 145460 130108 145472
rect 130160 145460 130166 145512
rect 161446 145500 161474 145540
rect 179414 145528 179420 145580
rect 179472 145568 179478 145580
rect 196526 145568 196532 145580
rect 179472 145540 196532 145568
rect 179472 145528 179478 145540
rect 196526 145528 196532 145540
rect 196584 145528 196590 145580
rect 179690 145500 179696 145512
rect 161446 145472 179696 145500
rect 179690 145460 179696 145472
rect 179748 145500 179754 145512
rect 189626 145500 189632 145512
rect 179748 145472 189632 145500
rect 179748 145460 179754 145472
rect 189626 145460 189632 145472
rect 189684 145460 189690 145512
rect 115474 144848 115480 144900
rect 115532 144888 115538 144900
rect 135346 144888 135352 144900
rect 115532 144860 135352 144888
rect 115532 144848 115538 144860
rect 135346 144848 135352 144860
rect 135404 144848 135410 144900
rect 174354 144848 174360 144900
rect 174412 144888 174418 144900
rect 196250 144888 196256 144900
rect 174412 144860 196256 144888
rect 174412 144848 174418 144860
rect 196250 144848 196256 144860
rect 196308 144848 196314 144900
rect 114186 144780 114192 144832
rect 114244 144820 114250 144832
rect 136174 144820 136180 144832
rect 114244 144792 136180 144820
rect 114244 144780 114250 144792
rect 136174 144780 136180 144792
rect 136232 144780 136238 144832
rect 168466 144780 168472 144832
rect 168524 144820 168530 144832
rect 194502 144820 194508 144832
rect 168524 144792 194508 144820
rect 168524 144780 168530 144792
rect 194502 144780 194508 144792
rect 194560 144780 194566 144832
rect 110874 144712 110880 144764
rect 110932 144752 110938 144764
rect 132034 144752 132040 144764
rect 110932 144724 132040 144752
rect 110932 144712 110938 144724
rect 132034 144712 132040 144724
rect 132092 144712 132098 144764
rect 171042 144712 171048 144764
rect 171100 144752 171106 144764
rect 196158 144752 196164 144764
rect 171100 144724 196164 144752
rect 171100 144712 171106 144724
rect 196158 144712 196164 144724
rect 196216 144712 196222 144764
rect 115290 144644 115296 144696
rect 115348 144684 115354 144696
rect 138014 144684 138020 144696
rect 115348 144656 138020 144684
rect 115348 144644 115354 144656
rect 138014 144644 138020 144656
rect 138072 144644 138078 144696
rect 165798 144644 165804 144696
rect 165856 144684 165862 144696
rect 192386 144684 192392 144696
rect 165856 144656 192392 144684
rect 165856 144644 165862 144656
rect 192386 144644 192392 144656
rect 192444 144644 192450 144696
rect 111518 144576 111524 144628
rect 111576 144616 111582 144628
rect 137278 144616 137284 144628
rect 111576 144588 137284 144616
rect 111576 144576 111582 144588
rect 137278 144576 137284 144588
rect 137336 144576 137342 144628
rect 156690 144576 156696 144628
rect 156748 144616 156754 144628
rect 189350 144616 189356 144628
rect 156748 144588 189356 144616
rect 156748 144576 156754 144588
rect 189350 144576 189356 144588
rect 189408 144576 189414 144628
rect 119982 144508 119988 144560
rect 120040 144548 120046 144560
rect 147766 144548 147772 144560
rect 120040 144520 147772 144548
rect 120040 144508 120046 144520
rect 147766 144508 147772 144520
rect 147824 144508 147830 144560
rect 159450 144508 159456 144560
rect 159508 144548 159514 144560
rect 192478 144548 192484 144560
rect 159508 144520 192484 144548
rect 159508 144508 159514 144520
rect 192478 144508 192484 144520
rect 192536 144508 192542 144560
rect 109770 144440 109776 144492
rect 109828 144480 109834 144492
rect 138934 144480 138940 144492
rect 109828 144452 138940 144480
rect 109828 144440 109834 144452
rect 138934 144440 138940 144452
rect 138992 144440 138998 144492
rect 155678 144440 155684 144492
rect 155736 144480 155742 144492
rect 189074 144480 189080 144492
rect 155736 144452 189080 144480
rect 155736 144440 155742 144452
rect 189074 144440 189080 144452
rect 189132 144440 189138 144492
rect 119706 144372 119712 144424
rect 119764 144412 119770 144424
rect 150526 144412 150532 144424
rect 119764 144384 150532 144412
rect 119764 144372 119770 144384
rect 150526 144372 150532 144384
rect 150584 144372 150590 144424
rect 155862 144372 155868 144424
rect 155920 144412 155926 144424
rect 191466 144412 191472 144424
rect 155920 144384 191472 144412
rect 155920 144372 155926 144384
rect 191466 144372 191472 144384
rect 191524 144372 191530 144424
rect 112530 144304 112536 144356
rect 112588 144344 112594 144356
rect 143902 144344 143908 144356
rect 112588 144316 143908 144344
rect 112588 144304 112594 144316
rect 143902 144304 143908 144316
rect 143960 144304 143966 144356
rect 160002 144304 160008 144356
rect 160060 144344 160066 144356
rect 193766 144344 193772 144356
rect 160060 144316 193772 144344
rect 160060 144304 160066 144316
rect 193766 144304 193772 144316
rect 193824 144304 193830 144356
rect 119338 144236 119344 144288
rect 119396 144276 119402 144288
rect 129182 144276 129188 144288
rect 119396 144248 129188 144276
rect 119396 144236 119402 144248
rect 129182 144236 129188 144248
rect 129240 144236 129246 144288
rect 130286 144236 130292 144288
rect 130344 144276 130350 144288
rect 189810 144276 189816 144288
rect 130344 144248 189816 144276
rect 130344 144236 130350 144248
rect 189810 144236 189816 144248
rect 189868 144236 189874 144288
rect 124950 144168 124956 144220
rect 125008 144208 125014 144220
rect 131482 144208 131488 144220
rect 125008 144180 131488 144208
rect 125008 144168 125014 144180
rect 131482 144168 131488 144180
rect 131540 144208 131546 144220
rect 580350 144208 580356 144220
rect 131540 144180 580356 144208
rect 131540 144168 131546 144180
rect 580350 144168 580356 144180
rect 580408 144168 580414 144220
rect 117682 144100 117688 144152
rect 117740 144140 117746 144152
rect 127894 144140 127900 144152
rect 117740 144112 127900 144140
rect 117740 144100 117746 144112
rect 127894 144100 127900 144112
rect 127952 144100 127958 144152
rect 175918 144100 175924 144152
rect 175976 144140 175982 144152
rect 194870 144140 194876 144152
rect 175976 144112 194876 144140
rect 175976 144100 175982 144112
rect 194870 144100 194876 144112
rect 194928 144100 194934 144152
rect 113726 144032 113732 144084
rect 113784 144072 113790 144084
rect 130286 144072 130292 144084
rect 113784 144044 130292 144072
rect 113784 144032 113790 144044
rect 130286 144032 130292 144044
rect 130344 144032 130350 144084
rect 180242 144032 180248 144084
rect 180300 144072 180306 144084
rect 189350 144072 189356 144084
rect 180300 144044 189356 144072
rect 180300 144032 180306 144044
rect 189350 144032 189356 144044
rect 189408 144032 189414 144084
rect 185854 143760 185860 143812
rect 185912 143800 185918 143812
rect 192386 143800 192392 143812
rect 185912 143772 192392 143800
rect 185912 143760 185918 143772
rect 192386 143760 192392 143772
rect 192444 143760 192450 143812
rect 115382 143488 115388 143540
rect 115440 143528 115446 143540
rect 124214 143528 124220 143540
rect 115440 143500 124220 143528
rect 115440 143488 115446 143500
rect 124214 143488 124220 143500
rect 124272 143488 124278 143540
rect 174906 143488 174912 143540
rect 174964 143528 174970 143540
rect 179506 143528 179512 143540
rect 174964 143500 179512 143528
rect 174964 143488 174970 143500
rect 179506 143488 179512 143500
rect 179564 143488 179570 143540
rect 185670 143488 185676 143540
rect 185728 143528 185734 143540
rect 189626 143528 189632 143540
rect 185728 143500 189632 143528
rect 185728 143488 185734 143500
rect 189626 143488 189632 143500
rect 189684 143488 189690 143540
rect 124858 143420 124864 143472
rect 124916 143460 124922 143472
rect 132862 143460 132868 143472
rect 124916 143432 132868 143460
rect 124916 143420 124922 143432
rect 132862 143420 132868 143432
rect 132920 143420 132926 143472
rect 176562 143420 176568 143472
rect 176620 143460 176626 143472
rect 178586 143460 178592 143472
rect 176620 143432 178592 143460
rect 176620 143420 176626 143432
rect 178586 143420 178592 143432
rect 178644 143420 178650 143472
rect 186222 143420 186228 143472
rect 186280 143460 186286 143472
rect 187786 143460 187792 143472
rect 186280 143432 187792 143460
rect 186280 143420 186286 143432
rect 187786 143420 187792 143432
rect 187844 143420 187850 143472
rect 118142 143352 118148 143404
rect 118200 143392 118206 143404
rect 127434 143392 127440 143404
rect 118200 143364 127440 143392
rect 118200 143352 118206 143364
rect 127434 143352 127440 143364
rect 127492 143352 127498 143404
rect 177482 143352 177488 143404
rect 177540 143392 177546 143404
rect 179414 143392 179420 143404
rect 177540 143364 179420 143392
rect 177540 143352 177546 143364
rect 179414 143352 179420 143364
rect 179472 143352 179478 143404
rect 116854 143284 116860 143336
rect 116912 143324 116918 143336
rect 128722 143324 128728 143336
rect 116912 143296 128728 143324
rect 116912 143284 116918 143296
rect 128722 143284 128728 143296
rect 128780 143284 128786 143336
rect 171410 143284 171416 143336
rect 171468 143324 171474 143336
rect 179782 143324 179788 143336
rect 171468 143296 179788 143324
rect 171468 143284 171474 143296
rect 179782 143284 179788 143296
rect 179840 143284 179846 143336
rect 114186 143216 114192 143268
rect 114244 143256 114250 143268
rect 129274 143256 129280 143268
rect 114244 143228 129280 143256
rect 114244 143216 114250 143228
rect 129274 143216 129280 143228
rect 129332 143216 129338 143268
rect 185578 143216 185584 143268
rect 185636 143256 185642 143268
rect 196342 143256 196348 143268
rect 185636 143228 196348 143256
rect 185636 143216 185642 143228
rect 196342 143216 196348 143228
rect 196400 143216 196406 143268
rect 118050 143148 118056 143200
rect 118108 143188 118114 143200
rect 131758 143188 131764 143200
rect 118108 143160 131764 143188
rect 118108 143148 118114 143160
rect 131758 143148 131764 143160
rect 131816 143148 131822 143200
rect 131850 143148 131856 143200
rect 131908 143188 131914 143200
rect 141142 143188 141148 143200
rect 131908 143160 141148 143188
rect 131908 143148 131914 143160
rect 141142 143148 141148 143160
rect 141200 143148 141206 143200
rect 165522 143148 165528 143200
rect 165580 143188 165586 143200
rect 189534 143188 189540 143200
rect 165580 143160 189540 143188
rect 165580 143148 165586 143160
rect 189534 143148 189540 143160
rect 189592 143148 189598 143200
rect 113910 143080 113916 143132
rect 113968 143120 113974 143132
rect 133414 143120 133420 143132
rect 113968 143092 133420 143120
rect 113968 143080 113974 143092
rect 133414 143080 133420 143092
rect 133472 143080 133478 143132
rect 160554 143080 160560 143132
rect 160612 143120 160618 143132
rect 190730 143120 190736 143132
rect 160612 143092 190736 143120
rect 160612 143080 160618 143092
rect 190730 143080 190736 143092
rect 190788 143080 190794 143132
rect 117958 143012 117964 143064
rect 118016 143052 118022 143064
rect 141694 143052 141700 143064
rect 118016 143024 141700 143052
rect 118016 143012 118022 143024
rect 141694 143012 141700 143024
rect 141752 143012 141758 143064
rect 156046 143012 156052 143064
rect 156104 143052 156110 143064
rect 191834 143052 191840 143064
rect 156104 143024 191840 143052
rect 156104 143012 156110 143024
rect 191834 143012 191840 143024
rect 191892 143012 191898 143064
rect 116670 142944 116676 142996
rect 116728 142984 116734 142996
rect 140038 142984 140044 142996
rect 116728 142956 140044 142984
rect 116728 142944 116734 142956
rect 140038 142944 140044 142956
rect 140096 142944 140102 142996
rect 154850 142944 154856 142996
rect 154908 142984 154914 142996
rect 191098 142984 191104 142996
rect 154908 142956 191104 142984
rect 154908 142944 154914 142956
rect 191098 142944 191104 142956
rect 191156 142944 191162 142996
rect 115198 142876 115204 142928
rect 115256 142916 115262 142928
rect 140774 142916 140780 142928
rect 115256 142888 140780 142916
rect 115256 142876 115262 142888
rect 140774 142876 140780 142888
rect 140832 142876 140838 142928
rect 168374 142876 168380 142928
rect 168432 142916 168438 142928
rect 211982 142916 211988 142928
rect 168432 142888 211988 142916
rect 168432 142876 168438 142888
rect 211982 142876 211988 142888
rect 212040 142876 212046 142928
rect 116578 142808 116584 142860
rect 116636 142848 116642 142860
rect 143534 142848 143540 142860
rect 116636 142820 143540 142848
rect 116636 142808 116642 142820
rect 143534 142808 143540 142820
rect 143592 142808 143598 142860
rect 150618 142808 150624 142860
rect 150676 142848 150682 142860
rect 213086 142848 213092 142860
rect 150676 142820 213092 142848
rect 150676 142808 150682 142820
rect 213086 142808 213092 142820
rect 213144 142808 213150 142860
rect 183462 142672 183468 142724
rect 183520 142712 183526 142724
rect 184474 142712 184480 142724
rect 183520 142684 184480 142712
rect 183520 142672 183526 142684
rect 184474 142672 184480 142684
rect 184532 142672 184538 142724
rect 128722 142468 128728 142520
rect 128780 142508 128786 142520
rect 137002 142508 137008 142520
rect 128780 142480 137008 142508
rect 128780 142468 128786 142480
rect 137002 142468 137008 142480
rect 137060 142468 137066 142520
rect 184842 142468 184848 142520
rect 184900 142508 184906 142520
rect 190822 142508 190828 142520
rect 184900 142480 190828 142508
rect 184900 142468 184906 142480
rect 190822 142468 190828 142480
rect 190880 142468 190886 142520
rect 129918 142400 129924 142452
rect 129976 142440 129982 142452
rect 133506 142440 133512 142452
rect 129976 142412 133512 142440
rect 129976 142400 129982 142412
rect 133506 142400 133512 142412
rect 133564 142400 133570 142452
rect 120626 142332 120632 142384
rect 120684 142372 120690 142384
rect 186222 142372 186228 142384
rect 120684 142344 186228 142372
rect 120684 142332 120690 142344
rect 186222 142332 186228 142344
rect 186280 142332 186286 142384
rect 128078 142264 128084 142316
rect 128136 142304 128142 142316
rect 549898 142304 549904 142316
rect 128136 142276 549904 142304
rect 128136 142264 128142 142276
rect 549898 142264 549904 142276
rect 549956 142264 549962 142316
rect 130102 142196 130108 142248
rect 130160 142236 130166 142248
rect 130160 142208 133460 142236
rect 130160 142196 130166 142208
rect 127986 142128 127992 142180
rect 128044 142168 128050 142180
rect 129826 142168 129832 142180
rect 128044 142140 129832 142168
rect 128044 142128 128050 142140
rect 129826 142128 129832 142140
rect 129884 142128 129890 142180
rect 130010 142128 130016 142180
rect 130068 142168 130074 142180
rect 132494 142168 132500 142180
rect 130068 142140 132500 142168
rect 130068 142128 130074 142140
rect 132494 142128 132500 142140
rect 132552 142128 132558 142180
rect 133432 142168 133460 142208
rect 133506 142196 133512 142248
rect 133564 142236 133570 142248
rect 579798 142236 579804 142248
rect 133564 142208 579804 142236
rect 133564 142196 133570 142208
rect 579798 142196 579804 142208
rect 579856 142196 579862 142248
rect 134518 142168 134524 142180
rect 133432 142140 134524 142168
rect 134518 142128 134524 142140
rect 134576 142128 134582 142180
rect 137002 142128 137008 142180
rect 137060 142168 137066 142180
rect 580810 142168 580816 142180
rect 137060 142140 580816 142168
rect 137060 142128 137066 142140
rect 580810 142128 580816 142140
rect 580868 142128 580874 142180
rect 112806 142060 112812 142112
rect 112864 142100 112870 142112
rect 125502 142100 125508 142112
rect 112864 142072 125508 142100
rect 112864 142060 112870 142072
rect 125502 142060 125508 142072
rect 125560 142060 125566 142112
rect 182726 142060 182732 142112
rect 182784 142100 182790 142112
rect 199102 142100 199108 142112
rect 182784 142072 199108 142100
rect 182784 142060 182790 142072
rect 199102 142060 199108 142072
rect 199160 142060 199166 142112
rect 112898 141992 112904 142044
rect 112956 142032 112962 142044
rect 127526 142032 127532 142044
rect 112956 142004 127532 142032
rect 112956 141992 112962 142004
rect 127526 141992 127532 142004
rect 127584 141992 127590 142044
rect 176010 141992 176016 142044
rect 176068 142032 176074 142044
rect 193950 142032 193956 142044
rect 176068 142004 193956 142032
rect 176068 141992 176074 142004
rect 193950 141992 193956 142004
rect 194008 141992 194014 142044
rect 115474 141924 115480 141976
rect 115532 141964 115538 141976
rect 130470 141964 130476 141976
rect 115532 141936 130476 141964
rect 115532 141924 115538 141936
rect 130470 141924 130476 141936
rect 130528 141924 130534 141976
rect 173802 141924 173808 141976
rect 173860 141964 173866 141976
rect 190638 141964 190644 141976
rect 173860 141936 190644 141964
rect 173860 141924 173866 141936
rect 190638 141924 190644 141936
rect 190696 141924 190702 141976
rect 114094 141856 114100 141908
rect 114152 141896 114158 141908
rect 135622 141896 135628 141908
rect 114152 141868 135628 141896
rect 114152 141856 114158 141868
rect 135622 141856 135628 141868
rect 135680 141856 135686 141908
rect 175090 141856 175096 141908
rect 175148 141896 175154 141908
rect 193858 141896 193864 141908
rect 175148 141868 193864 141896
rect 175148 141856 175154 141868
rect 193858 141856 193864 141868
rect 193916 141856 193922 141908
rect 115566 141788 115572 141840
rect 115624 141828 115630 141840
rect 138382 141828 138388 141840
rect 115624 141800 138388 141828
rect 115624 141788 115630 141800
rect 138382 141788 138388 141800
rect 138440 141788 138446 141840
rect 168742 141788 168748 141840
rect 168800 141828 168806 141840
rect 189258 141828 189264 141840
rect 168800 141800 189264 141828
rect 168800 141788 168806 141800
rect 189258 141788 189264 141800
rect 189316 141788 189322 141840
rect 112622 141720 112628 141772
rect 112680 141760 112686 141772
rect 141602 141760 141608 141772
rect 112680 141732 141608 141760
rect 112680 141720 112686 141732
rect 141602 141720 141608 141732
rect 141660 141720 141666 141772
rect 166810 141720 166816 141772
rect 166868 141760 166874 141772
rect 190914 141760 190920 141772
rect 166868 141732 190920 141760
rect 166868 141720 166874 141732
rect 190914 141720 190920 141732
rect 190972 141720 190978 141772
rect 116394 141652 116400 141704
rect 116452 141692 116458 141704
rect 147214 141692 147220 141704
rect 116452 141664 147220 141692
rect 116452 141652 116458 141664
rect 147214 141652 147220 141664
rect 147272 141652 147278 141704
rect 156966 141652 156972 141704
rect 157024 141692 157030 141704
rect 189902 141692 189908 141704
rect 157024 141664 189908 141692
rect 157024 141652 157030 141664
rect 189902 141652 189908 141664
rect 189960 141652 189966 141704
rect 115106 141584 115112 141636
rect 115164 141624 115170 141636
rect 146846 141624 146852 141636
rect 115164 141596 146852 141624
rect 115164 141584 115170 141596
rect 146846 141584 146852 141596
rect 146904 141584 146910 141636
rect 157426 141584 157432 141636
rect 157484 141624 157490 141636
rect 192294 141624 192300 141636
rect 157484 141596 192300 141624
rect 157484 141584 157490 141596
rect 192294 141584 192300 141596
rect 192352 141584 192358 141636
rect 116854 141516 116860 141568
rect 116912 141556 116918 141568
rect 149606 141556 149612 141568
rect 116912 141528 149612 141556
rect 116912 141516 116918 141528
rect 149606 141516 149612 141528
rect 149664 141516 149670 141568
rect 154758 141516 154764 141568
rect 154816 141556 154822 141568
rect 190822 141556 190828 141568
rect 154816 141528 190828 141556
rect 154816 141516 154822 141528
rect 190822 141516 190828 141528
rect 190880 141516 190886 141568
rect 113726 141448 113732 141500
rect 113784 141488 113790 141500
rect 148226 141488 148232 141500
rect 113784 141460 148232 141488
rect 113784 141448 113790 141460
rect 148226 141448 148232 141460
rect 148284 141448 148290 141500
rect 163774 141448 163780 141500
rect 163832 141488 163838 141500
rect 204622 141488 204628 141500
rect 163832 141460 204628 141488
rect 163832 141448 163838 141460
rect 204622 141448 204628 141460
rect 204680 141448 204686 141500
rect 112806 141380 112812 141432
rect 112864 141420 112870 141432
rect 153654 141420 153660 141432
rect 112864 141392 153660 141420
rect 112864 141380 112870 141392
rect 153654 141380 153660 141392
rect 153712 141380 153718 141432
rect 154666 141380 154672 141432
rect 154724 141420 154730 141432
rect 213178 141420 213184 141432
rect 154724 141392 213184 141420
rect 154724 141380 154730 141392
rect 213178 141380 213184 141392
rect 213236 141380 213242 141432
rect 118326 141312 118332 141364
rect 118384 141352 118390 141364
rect 129366 141352 129372 141364
rect 118384 141324 129372 141352
rect 118384 141312 118390 141324
rect 129366 141312 129372 141324
rect 129424 141312 129430 141364
rect 179506 141312 179512 141364
rect 179564 141352 179570 141364
rect 180610 141352 180616 141364
rect 179564 141324 180616 141352
rect 179564 141312 179570 141324
rect 180610 141312 180616 141324
rect 180668 141352 180674 141364
rect 193674 141352 193680 141364
rect 180668 141324 193680 141352
rect 180668 141312 180674 141324
rect 193674 141312 193680 141324
rect 193732 141312 193738 141364
rect 184290 141244 184296 141296
rect 184348 141284 184354 141296
rect 196526 141284 196532 141296
rect 184348 141256 196532 141284
rect 184348 141244 184354 141256
rect 196526 141244 196532 141256
rect 196584 141244 196590 141296
rect 186038 141176 186044 141228
rect 186096 141216 186102 141228
rect 197998 141216 198004 141228
rect 186096 141188 198004 141216
rect 186096 141176 186102 141188
rect 197998 141176 198004 141188
rect 198056 141176 198062 141228
rect 119062 140836 119068 140888
rect 119120 140876 119126 140888
rect 179506 140876 179512 140888
rect 119120 140848 179512 140876
rect 119120 140836 119126 140848
rect 179506 140836 179512 140848
rect 179564 140836 179570 140888
rect 8938 140768 8944 140820
rect 8996 140808 9002 140820
rect 183186 140808 183192 140820
rect 8996 140780 183192 140808
rect 8996 140768 9002 140780
rect 183186 140768 183192 140780
rect 183244 140768 183250 140820
rect 129734 140700 129740 140752
rect 129792 140740 129798 140752
rect 130654 140740 130660 140752
rect 129792 140712 130660 140740
rect 129792 140700 129798 140712
rect 130654 140700 130660 140712
rect 130712 140700 130718 140752
rect 142154 140700 142160 140752
rect 142212 140740 142218 140752
rect 142798 140740 142804 140752
rect 142212 140712 142804 140740
rect 142212 140700 142218 140712
rect 142798 140700 142804 140712
rect 142856 140700 142862 140752
rect 149238 140700 149244 140752
rect 149296 140740 149302 140752
rect 149514 140740 149520 140752
rect 149296 140712 149520 140740
rect 149296 140700 149302 140712
rect 149514 140700 149520 140712
rect 149572 140700 149578 140752
rect 151814 140700 151820 140752
rect 151872 140740 151878 140752
rect 152734 140740 152740 140752
rect 151872 140712 152740 140740
rect 151872 140700 151878 140712
rect 152734 140700 152740 140712
rect 152792 140700 152798 140752
rect 157334 140700 157340 140752
rect 157392 140740 157398 140752
rect 158254 140740 158260 140752
rect 157392 140712 158260 140740
rect 157392 140700 157398 140712
rect 158254 140700 158260 140712
rect 158312 140700 158318 140752
rect 166994 140700 167000 140752
rect 167052 140740 167058 140752
rect 167638 140740 167644 140752
rect 167052 140712 167644 140740
rect 167052 140700 167058 140712
rect 167638 140700 167644 140712
rect 167696 140700 167702 140752
rect 168834 140700 168840 140752
rect 168892 140740 168898 140752
rect 169294 140740 169300 140752
rect 168892 140712 169300 140740
rect 168892 140700 168898 140712
rect 169294 140700 169300 140712
rect 169352 140700 169358 140752
rect 169754 140700 169760 140752
rect 169812 140740 169818 140752
rect 193674 140740 193680 140752
rect 169812 140712 193680 140740
rect 169812 140700 169818 140712
rect 193674 140700 193680 140712
rect 193732 140700 193738 140752
rect 117958 140632 117964 140684
rect 118016 140672 118022 140684
rect 127710 140672 127716 140684
rect 118016 140644 127716 140672
rect 118016 140632 118022 140644
rect 127710 140632 127716 140644
rect 127768 140632 127774 140684
rect 176654 140632 176660 140684
rect 176712 140672 176718 140684
rect 177574 140672 177580 140684
rect 176712 140644 177580 140672
rect 176712 140632 176718 140644
rect 177574 140632 177580 140644
rect 177632 140632 177638 140684
rect 178034 140632 178040 140684
rect 178092 140672 178098 140684
rect 178678 140672 178684 140684
rect 178092 140644 178684 140672
rect 178092 140632 178098 140644
rect 178678 140632 178684 140644
rect 178736 140632 178742 140684
rect 118050 140564 118056 140616
rect 118108 140604 118114 140616
rect 127802 140604 127808 140616
rect 118108 140576 127808 140604
rect 118108 140564 118114 140576
rect 127802 140564 127808 140576
rect 127860 140564 127866 140616
rect 112898 140496 112904 140548
rect 112956 140536 112962 140548
rect 123386 140536 123392 140548
rect 112956 140508 123392 140536
rect 112956 140496 112962 140508
rect 123386 140496 123392 140508
rect 123444 140496 123450 140548
rect 117866 140428 117872 140480
rect 117924 140468 117930 140480
rect 129090 140468 129096 140480
rect 117924 140440 129096 140468
rect 117924 140428 117930 140440
rect 129090 140428 129096 140440
rect 129148 140428 129154 140480
rect 116670 140360 116676 140412
rect 116728 140400 116734 140412
rect 128998 140400 129004 140412
rect 116728 140372 129004 140400
rect 116728 140360 116734 140372
rect 128998 140360 129004 140372
rect 129056 140360 129062 140412
rect 114094 140292 114100 140344
rect 114152 140332 114158 140344
rect 130378 140332 130384 140344
rect 114152 140304 130384 140332
rect 114152 140292 114158 140304
rect 130378 140292 130384 140304
rect 130436 140292 130442 140344
rect 180058 140292 180064 140344
rect 180116 140332 180122 140344
rect 189166 140332 189172 140344
rect 180116 140304 189172 140332
rect 180116 140292 180122 140304
rect 189166 140292 189172 140304
rect 189224 140292 189230 140344
rect 120718 140224 120724 140276
rect 120776 140264 120782 140276
rect 151170 140264 151176 140276
rect 120776 140236 151176 140264
rect 120776 140224 120782 140236
rect 151170 140224 151176 140236
rect 151228 140224 151234 140276
rect 183094 140224 183100 140276
rect 183152 140264 183158 140276
rect 193766 140264 193772 140276
rect 183152 140236 193772 140264
rect 183152 140224 183158 140236
rect 193766 140224 193772 140236
rect 193824 140224 193830 140276
rect 115290 140156 115296 140208
rect 115348 140196 115354 140208
rect 148134 140196 148140 140208
rect 115348 140168 148140 140196
rect 115348 140156 115354 140168
rect 148134 140156 148140 140168
rect 148192 140156 148198 140208
rect 176194 140156 176200 140208
rect 176252 140196 176258 140208
rect 188154 140196 188160 140208
rect 176252 140168 188160 140196
rect 176252 140156 176258 140168
rect 188154 140156 188160 140168
rect 188212 140156 188218 140208
rect 188706 140156 188712 140208
rect 188764 140196 188770 140208
rect 191006 140196 191012 140208
rect 188764 140168 191012 140196
rect 188764 140156 188770 140168
rect 191006 140156 191012 140168
rect 191064 140156 191070 140208
rect 117774 140088 117780 140140
rect 117832 140128 117838 140140
rect 151262 140128 151268 140140
rect 117832 140100 151268 140128
rect 117832 140088 117838 140100
rect 151262 140088 151268 140100
rect 151320 140088 151326 140140
rect 155770 140088 155776 140140
rect 155828 140088 155834 140140
rect 178586 140088 178592 140140
rect 178644 140128 178650 140140
rect 206002 140128 206008 140140
rect 178644 140100 206008 140128
rect 178644 140088 178650 140100
rect 206002 140088 206008 140100
rect 206060 140088 206066 140140
rect 104250 140020 104256 140072
rect 104308 140060 104314 140072
rect 138290 140060 138296 140072
rect 104308 140032 138296 140060
rect 104308 140020 104314 140032
rect 138290 140020 138296 140032
rect 138348 140020 138354 140072
rect 155788 140060 155816 140088
rect 155788 140032 180794 140060
rect 119246 139952 119252 140004
rect 119304 139992 119310 140004
rect 126422 139992 126428 140004
rect 119304 139964 126428 139992
rect 119304 139952 119310 139964
rect 126422 139952 126428 139964
rect 126480 139952 126486 140004
rect 180766 139992 180794 140032
rect 189994 140020 190000 140072
rect 190052 140060 190058 140072
rect 190914 140060 190920 140072
rect 190052 140032 190920 140060
rect 190052 140020 190058 140032
rect 190914 140020 190920 140032
rect 190972 140020 190978 140072
rect 191190 139992 191196 140004
rect 180766 139964 191196 139992
rect 191190 139952 191196 139964
rect 191248 139952 191254 140004
rect 125686 139884 125692 139936
rect 125744 139924 125750 139936
rect 126330 139924 126336 139936
rect 125744 139896 126336 139924
rect 125744 139884 125750 139896
rect 126330 139884 126336 139896
rect 126388 139884 126394 139936
rect 187326 139884 187332 139936
rect 187384 139924 187390 139936
rect 192294 139924 192300 139936
rect 187384 139896 192300 139924
rect 187384 139884 187390 139896
rect 192294 139884 192300 139896
rect 192352 139884 192358 139936
rect 187142 139816 187148 139868
rect 187200 139856 187206 139868
rect 189442 139856 189448 139868
rect 187200 139828 189448 139856
rect 187200 139816 187206 139828
rect 189442 139816 189448 139828
rect 189500 139816 189506 139868
rect 192846 139856 192852 139868
rect 190426 139828 192852 139856
rect 187234 139748 187240 139800
rect 187292 139788 187298 139800
rect 190426 139788 190454 139828
rect 192846 139816 192852 139828
rect 192904 139816 192910 139868
rect 187292 139760 190454 139788
rect 187292 139748 187298 139760
rect 173250 139680 173256 139732
rect 173308 139720 173314 139732
rect 199010 139720 199016 139732
rect 173308 139692 199016 139720
rect 173308 139680 173314 139692
rect 199010 139680 199016 139692
rect 199068 139680 199074 139732
rect 161474 139612 161480 139664
rect 161532 139652 161538 139664
rect 194778 139652 194784 139664
rect 161532 139624 194784 139652
rect 161532 139612 161538 139624
rect 194778 139612 194784 139624
rect 194836 139612 194842 139664
rect 95970 139544 95976 139596
rect 96028 139584 96034 139596
rect 182174 139584 182180 139596
rect 96028 139556 182180 139584
rect 96028 139544 96034 139556
rect 182174 139544 182180 139556
rect 182232 139544 182238 139596
rect 4798 139476 4804 139528
rect 4856 139516 4862 139528
rect 180794 139516 180800 139528
rect 4856 139488 180800 139516
rect 4856 139476 4862 139488
rect 180794 139476 180800 139488
rect 180852 139516 180858 139528
rect 181438 139516 181444 139528
rect 180852 139488 181444 139516
rect 180852 139476 180858 139488
rect 181438 139476 181444 139488
rect 181496 139476 181502 139528
rect 182634 139476 182640 139528
rect 182692 139516 182698 139528
rect 192110 139516 192116 139528
rect 182692 139488 192116 139516
rect 182692 139476 182698 139488
rect 192110 139476 192116 139488
rect 192168 139476 192174 139528
rect 113634 139408 113640 139460
rect 113692 139448 113698 139460
rect 122190 139448 122196 139460
rect 113692 139420 122196 139448
rect 113692 139408 113698 139420
rect 122190 139408 122196 139420
rect 122248 139408 122254 139460
rect 126146 139408 126152 139460
rect 126204 139448 126210 139460
rect 327718 139448 327724 139460
rect 126204 139420 327724 139448
rect 126204 139408 126210 139420
rect 327718 139408 327724 139420
rect 327776 139408 327782 139460
rect 184658 139340 184664 139392
rect 184716 139380 184722 139392
rect 186498 139380 186504 139392
rect 184716 139352 186504 139380
rect 184716 139340 184722 139352
rect 186498 139340 186504 139352
rect 186556 139340 186562 139392
rect 188430 139272 188436 139324
rect 188488 139312 188494 139324
rect 192478 139312 192484 139324
rect 188488 139284 192484 139312
rect 188488 139272 188494 139284
rect 192478 139272 192484 139284
rect 192536 139272 192542 139324
rect 188246 138864 188252 138916
rect 188304 138904 188310 138916
rect 195330 138904 195336 138916
rect 188304 138876 195336 138904
rect 188304 138864 188310 138876
rect 195330 138864 195336 138876
rect 195388 138864 195394 138916
rect 188798 138796 188804 138848
rect 188856 138836 188862 138848
rect 196434 138836 196440 138848
rect 188856 138808 196440 138836
rect 188856 138796 188862 138808
rect 196434 138796 196440 138808
rect 196492 138796 196498 138848
rect 188522 138728 188528 138780
rect 188580 138768 188586 138780
rect 199378 138768 199384 138780
rect 188580 138740 199384 138768
rect 188580 138728 188586 138740
rect 199378 138728 199384 138740
rect 199436 138728 199442 138780
rect 3418 138660 3424 138712
rect 3476 138700 3482 138712
rect 120626 138700 120632 138712
rect 3476 138672 120632 138700
rect 3476 138660 3482 138672
rect 120626 138660 120632 138672
rect 120684 138660 120690 138712
rect 188154 138660 188160 138712
rect 188212 138700 188218 138712
rect 203610 138700 203616 138712
rect 188212 138672 203616 138700
rect 188212 138660 188218 138672
rect 203610 138660 203616 138672
rect 203668 138660 203674 138712
rect 191282 138116 191288 138168
rect 191340 138156 191346 138168
rect 198182 138156 198188 138168
rect 191340 138128 198188 138156
rect 191340 138116 191346 138128
rect 198182 138116 198188 138128
rect 198240 138116 198246 138168
rect 188614 137980 188620 138032
rect 188672 138020 188678 138032
rect 189994 138020 190000 138032
rect 188672 137992 190000 138020
rect 188672 137980 188678 137992
rect 189994 137980 190000 137992
rect 190052 137980 190058 138032
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 119062 137952 119068 137964
rect 3292 137924 119068 137952
rect 3292 137912 3298 137924
rect 119062 137912 119068 137924
rect 119120 137912 119126 137964
rect 188154 137776 188160 137828
rect 188212 137816 188218 137828
rect 202138 137816 202144 137828
rect 188212 137788 202144 137816
rect 188212 137776 188218 137788
rect 202138 137776 202144 137788
rect 202196 137776 202202 137828
rect 188890 136688 188896 136740
rect 188948 136728 188954 136740
rect 202230 136728 202236 136740
rect 188948 136700 202236 136728
rect 188948 136688 188954 136700
rect 202230 136688 202236 136700
rect 202288 136688 202294 136740
rect 202322 136552 202328 136604
rect 202380 136592 202386 136604
rect 206462 136592 206468 136604
rect 202380 136564 206468 136592
rect 202380 136552 202386 136564
rect 206462 136552 206468 136564
rect 206520 136552 206526 136604
rect 195422 124856 195428 124908
rect 195480 124896 195486 124908
rect 204806 124896 204812 124908
rect 195480 124868 204812 124896
rect 195480 124856 195486 124868
rect 204806 124856 204812 124868
rect 204864 124856 204870 124908
rect 192570 122068 192576 122120
rect 192628 122108 192634 122120
rect 202322 122108 202328 122120
rect 192628 122080 202328 122108
rect 192628 122068 192634 122080
rect 202322 122068 202328 122080
rect 202380 122068 202386 122120
rect 191190 118668 191196 118720
rect 191248 118708 191254 118720
rect 191926 118708 191932 118720
rect 191248 118680 191932 118708
rect 191248 118668 191254 118680
rect 191926 118668 191932 118680
rect 191984 118668 191990 118720
rect 189718 114520 189724 114572
rect 189776 114560 189782 114572
rect 191098 114560 191104 114572
rect 189776 114532 191104 114560
rect 189776 114520 189782 114532
rect 191098 114520 191104 114532
rect 191156 114520 191162 114572
rect 189994 114384 190000 114436
rect 190052 114424 190058 114436
rect 192570 114424 192576 114436
rect 190052 114396 192576 114424
rect 190052 114384 190058 114396
rect 192570 114384 192576 114396
rect 192628 114384 192634 114436
rect 189902 113840 189908 113892
rect 189960 113880 189966 113892
rect 191190 113880 191196 113892
rect 189960 113852 191196 113880
rect 189960 113840 189966 113852
rect 191190 113840 191196 113852
rect 191248 113840 191254 113892
rect 189810 113704 189816 113756
rect 189868 113744 189874 113756
rect 191926 113744 191932 113756
rect 189868 113716 191932 113744
rect 189868 113704 189874 113716
rect 191926 113704 191932 113716
rect 191984 113704 191990 113756
rect 2774 110780 2780 110832
rect 2832 110820 2838 110832
rect 4798 110820 4804 110832
rect 2832 110792 4804 110820
rect 2832 110780 2838 110792
rect 4798 110780 4804 110792
rect 4856 110780 4862 110832
rect 115014 110440 115020 110492
rect 115072 110480 115078 110492
rect 120718 110480 120724 110492
rect 115072 110452 120724 110480
rect 115072 110440 115078 110452
rect 120718 110440 120724 110452
rect 120776 110440 120782 110492
rect 549898 100648 549904 100700
rect 549956 100688 549962 100700
rect 579614 100688 579620 100700
rect 549956 100660 579620 100688
rect 549956 100648 549962 100660
rect 579614 100648 579620 100660
rect 579672 100648 579678 100700
rect 105630 89088 105636 89140
rect 105688 89088 105694 89140
rect 105648 88924 105676 89088
rect 105722 88924 105728 88936
rect 105648 88896 105728 88924
rect 105722 88884 105728 88896
rect 105780 88884 105786 88936
rect 482278 86912 482284 86964
rect 482336 86952 482342 86964
rect 579614 86952 579620 86964
rect 482336 86924 579620 86952
rect 482336 86912 482342 86924
rect 579614 86912 579620 86924
rect 579672 86912 579678 86964
rect 197906 86776 197912 86828
rect 197964 86816 197970 86828
rect 197964 86788 198044 86816
rect 197964 86776 197970 86788
rect 198016 86624 198044 86788
rect 197998 86572 198004 86624
rect 198056 86572 198062 86624
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 95970 85524 95976 85536
rect 3568 85496 95976 85524
rect 3568 85484 3574 85496
rect 95970 85484 95976 85496
rect 96028 85484 96034 85536
rect 188890 82764 188896 82816
rect 188948 82804 188954 82816
rect 203702 82804 203708 82816
rect 188948 82776 203708 82804
rect 188948 82764 188954 82776
rect 203702 82764 203708 82776
rect 203760 82764 203766 82816
rect 188982 82084 188988 82136
rect 189040 82124 189046 82136
rect 196158 82124 196164 82136
rect 189040 82096 196164 82124
rect 189040 82084 189046 82096
rect 196158 82084 196164 82096
rect 196216 82084 196222 82136
rect 215846 81064 215852 81116
rect 215904 81104 215910 81116
rect 216122 81104 216128 81116
rect 215904 81076 216128 81104
rect 215904 81064 215910 81076
rect 216122 81064 216128 81076
rect 216180 81064 216186 81116
rect 114922 80996 114928 81048
rect 114980 81036 114986 81048
rect 120718 81036 120724 81048
rect 114980 81008 120724 81036
rect 114980 80996 114986 81008
rect 120718 80996 120724 81008
rect 120776 80996 120782 81048
rect 109494 80860 109500 80912
rect 109552 80900 109558 80912
rect 120810 80900 120816 80912
rect 109552 80872 120816 80900
rect 109552 80860 109558 80872
rect 120810 80860 120816 80872
rect 120868 80860 120874 80912
rect 105170 80792 105176 80844
rect 105228 80832 105234 80844
rect 120074 80832 120080 80844
rect 105228 80804 120080 80832
rect 105228 80792 105234 80804
rect 120074 80792 120080 80804
rect 120132 80792 120138 80844
rect 120994 80792 121000 80844
rect 121052 80832 121058 80844
rect 205082 80832 205088 80844
rect 121052 80804 146662 80832
rect 121052 80792 121058 80804
rect 112438 80724 112444 80776
rect 112496 80764 112502 80776
rect 112496 80736 145650 80764
rect 112496 80724 112502 80736
rect 112346 80656 112352 80708
rect 112404 80696 112410 80708
rect 112404 80668 145512 80696
rect 112404 80656 112410 80668
rect 118694 80588 118700 80640
rect 118752 80628 118758 80640
rect 118752 80600 141648 80628
rect 118752 80588 118758 80600
rect 121086 80520 121092 80572
rect 121144 80560 121150 80572
rect 121144 80532 141556 80560
rect 121144 80520 121150 80532
rect 121178 80452 121184 80504
rect 121236 80492 121242 80504
rect 121236 80464 141464 80492
rect 121236 80452 121242 80464
rect 102778 80384 102784 80436
rect 102836 80424 102842 80436
rect 124858 80424 124864 80436
rect 102836 80396 124864 80424
rect 102836 80384 102842 80396
rect 124858 80384 124864 80396
rect 124916 80384 124922 80436
rect 131942 80384 131948 80436
rect 132000 80424 132006 80436
rect 132000 80396 138658 80424
rect 132000 80384 132006 80396
rect 131758 80316 131764 80368
rect 131816 80356 131822 80368
rect 131816 80328 137738 80356
rect 131816 80316 131822 80328
rect 131666 80112 131672 80164
rect 131724 80152 131730 80164
rect 131724 80124 134978 80152
rect 131724 80112 131730 80124
rect 130378 80044 130384 80096
rect 130436 80084 130442 80096
rect 134950 80084 134978 80124
rect 130436 80056 133184 80084
rect 134950 80056 137508 80084
rect 130436 80044 130442 80056
rect 130470 79976 130476 80028
rect 130528 80016 130534 80028
rect 130528 79988 132494 80016
rect 130528 79976 130534 79988
rect 132466 79948 132494 79988
rect 133000 79948 133006 79960
rect 132466 79920 133006 79948
rect 133000 79908 133006 79920
rect 133058 79908 133064 79960
rect 132632 79880 132638 79892
rect 132604 79840 132638 79880
rect 132690 79840 132696 79892
rect 133156 79880 133184 80056
rect 134398 79988 134886 80016
rect 133644 79948 133650 79960
rect 133616 79908 133650 79948
rect 133702 79908 133708 79960
rect 134104 79908 134110 79960
rect 134162 79908 134168 79960
rect 133276 79880 133282 79892
rect 133156 79852 133282 79880
rect 133276 79840 133282 79852
rect 133334 79840 133340 79892
rect 133368 79840 133374 79892
rect 133426 79840 133432 79892
rect 133460 79840 133466 79892
rect 133518 79880 133524 79892
rect 133518 79840 133552 79880
rect 113726 79772 113732 79824
rect 113784 79812 113790 79824
rect 113784 79784 132448 79812
rect 113784 79772 113790 79784
rect 99834 79704 99840 79756
rect 99892 79744 99898 79756
rect 132310 79744 132316 79756
rect 99892 79716 132316 79744
rect 99892 79704 99898 79716
rect 132310 79704 132316 79716
rect 132368 79704 132374 79756
rect 120534 79636 120540 79688
rect 120592 79676 120598 79688
rect 130562 79676 130568 79688
rect 120592 79648 130568 79676
rect 120592 79636 120598 79648
rect 130562 79636 130568 79648
rect 130620 79676 130626 79688
rect 131022 79676 131028 79688
rect 130620 79648 131028 79676
rect 130620 79636 130626 79648
rect 131022 79636 131028 79648
rect 131080 79636 131086 79688
rect 132420 79676 132448 79784
rect 132604 79756 132632 79840
rect 133092 79772 133098 79824
rect 133150 79772 133156 79824
rect 132586 79704 132592 79756
rect 132644 79704 132650 79756
rect 133110 79688 133138 79772
rect 132770 79676 132776 79688
rect 132420 79648 132776 79676
rect 132770 79636 132776 79648
rect 132828 79636 132834 79688
rect 132954 79676 132960 79688
rect 132880 79648 132960 79676
rect 109678 79568 109684 79620
rect 109736 79608 109742 79620
rect 123754 79608 123760 79620
rect 109736 79580 123760 79608
rect 109736 79568 109742 79580
rect 123754 79568 123760 79580
rect 123812 79568 123818 79620
rect 127066 79568 127072 79620
rect 127124 79608 127130 79620
rect 132880 79608 132908 79648
rect 132954 79636 132960 79648
rect 133012 79636 133018 79688
rect 133046 79636 133052 79688
rect 133104 79648 133138 79688
rect 133104 79636 133110 79648
rect 127124 79580 132908 79608
rect 133386 79620 133414 79840
rect 133524 79688 133552 79840
rect 133506 79636 133512 79688
rect 133564 79636 133570 79688
rect 133386 79580 133420 79620
rect 127124 79568 127130 79580
rect 133414 79568 133420 79580
rect 133472 79568 133478 79620
rect 106918 79500 106924 79552
rect 106976 79540 106982 79552
rect 122834 79540 122840 79552
rect 106976 79512 122840 79540
rect 106976 79500 106982 79512
rect 122834 79500 122840 79512
rect 122892 79540 122898 79552
rect 124122 79540 124128 79552
rect 122892 79512 124128 79540
rect 122892 79500 122898 79512
rect 124122 79500 124128 79512
rect 124180 79500 124186 79552
rect 128630 79500 128636 79552
rect 128688 79540 128694 79552
rect 133138 79540 133144 79552
rect 128688 79512 133144 79540
rect 128688 79500 128694 79512
rect 133138 79500 133144 79512
rect 133196 79500 133202 79552
rect 108022 79432 108028 79484
rect 108080 79472 108086 79484
rect 108666 79472 108672 79484
rect 108080 79444 108672 79472
rect 108080 79432 108086 79444
rect 108666 79432 108672 79444
rect 108724 79432 108730 79484
rect 113634 79432 113640 79484
rect 113692 79472 113698 79484
rect 113692 79444 127572 79472
rect 113692 79432 113698 79444
rect 108390 79364 108396 79416
rect 108448 79404 108454 79416
rect 126974 79404 126980 79416
rect 108448 79376 126980 79404
rect 108448 79364 108454 79376
rect 126974 79364 126980 79376
rect 127032 79364 127038 79416
rect 127544 79404 127572 79444
rect 132494 79432 132500 79484
rect 132552 79472 132558 79484
rect 133616 79472 133644 79908
rect 133828 79840 133834 79892
rect 133886 79840 133892 79892
rect 133920 79840 133926 79892
rect 133978 79880 133984 79892
rect 133978 79840 134012 79880
rect 133846 79756 133874 79840
rect 133846 79716 133880 79756
rect 133874 79704 133880 79716
rect 133932 79704 133938 79756
rect 133782 79636 133788 79688
rect 133840 79676 133846 79688
rect 133984 79676 134012 79840
rect 134122 79744 134150 79908
rect 134122 79716 134196 79744
rect 133840 79648 134012 79676
rect 133840 79636 133846 79648
rect 133966 79568 133972 79620
rect 134024 79608 134030 79620
rect 134168 79608 134196 79716
rect 134024 79580 134196 79608
rect 134024 79568 134030 79580
rect 134398 79540 134426 79988
rect 134858 79960 134886 79988
rect 134472 79908 134478 79960
rect 134530 79908 134536 79960
rect 134840 79908 134846 79960
rect 134898 79908 134904 79960
rect 134932 79908 134938 79960
rect 134990 79908 134996 79960
rect 136036 79948 136042 79960
rect 135088 79920 136042 79948
rect 134490 79620 134518 79908
rect 134656 79840 134662 79892
rect 134714 79840 134720 79892
rect 134674 79812 134702 79840
rect 134628 79784 134702 79812
rect 134628 79620 134656 79784
rect 134950 79688 134978 79908
rect 135088 79688 135116 79920
rect 136036 79908 136042 79920
rect 136094 79908 136100 79960
rect 136192 79920 136450 79948
rect 135668 79840 135674 79892
rect 135726 79840 135732 79892
rect 135760 79840 135766 79892
rect 135818 79880 135824 79892
rect 135818 79852 136036 79880
rect 135818 79840 135824 79852
rect 135208 79812 135214 79824
rect 135180 79772 135214 79812
rect 135266 79772 135272 79824
rect 135392 79772 135398 79824
rect 135450 79772 135456 79824
rect 135484 79772 135490 79824
rect 135542 79772 135548 79824
rect 134886 79636 134892 79688
rect 134944 79648 134978 79688
rect 134944 79636 134950 79648
rect 135070 79636 135076 79688
rect 135128 79636 135134 79688
rect 135180 79620 135208 79772
rect 135410 79620 135438 79772
rect 135502 79688 135530 79772
rect 135502 79648 135536 79688
rect 135530 79636 135536 79648
rect 135588 79636 135594 79688
rect 134490 79580 134524 79620
rect 134518 79568 134524 79580
rect 134576 79568 134582 79620
rect 134610 79568 134616 79620
rect 134668 79568 134674 79620
rect 135162 79568 135168 79620
rect 135220 79568 135226 79620
rect 135346 79568 135352 79620
rect 135404 79580 135438 79620
rect 135404 79568 135410 79580
rect 134794 79540 134800 79552
rect 134398 79512 134800 79540
rect 134794 79500 134800 79512
rect 134852 79500 134858 79552
rect 132552 79444 133644 79472
rect 132552 79432 132558 79444
rect 130838 79404 130844 79416
rect 127544 79376 130844 79404
rect 130838 79364 130844 79376
rect 130896 79364 130902 79416
rect 131022 79364 131028 79416
rect 131080 79404 131086 79416
rect 131080 79376 132448 79404
rect 131080 79364 131086 79376
rect 96062 79296 96068 79348
rect 96120 79296 96126 79348
rect 108206 79296 108212 79348
rect 108264 79336 108270 79348
rect 131206 79336 131212 79348
rect 108264 79308 131212 79336
rect 108264 79296 108270 79308
rect 131206 79296 131212 79308
rect 131264 79336 131270 79348
rect 132310 79336 132316 79348
rect 131264 79308 132316 79336
rect 131264 79296 131270 79308
rect 132310 79296 132316 79308
rect 132368 79296 132374 79348
rect 132420 79336 132448 79376
rect 132770 79364 132776 79416
rect 132828 79404 132834 79416
rect 134242 79404 134248 79416
rect 132828 79376 134248 79404
rect 132828 79364 132834 79376
rect 134242 79364 134248 79376
rect 134300 79364 134306 79416
rect 135438 79364 135444 79416
rect 135496 79404 135502 79416
rect 135686 79404 135714 79840
rect 135852 79772 135858 79824
rect 135910 79772 135916 79824
rect 135870 79620 135898 79772
rect 135806 79568 135812 79620
rect 135864 79580 135898 79620
rect 135864 79568 135870 79580
rect 136008 79484 136036 79852
rect 136192 79552 136220 79920
rect 136422 79892 136450 79920
rect 136588 79908 136594 79960
rect 136646 79908 136652 79960
rect 136864 79908 136870 79960
rect 136922 79908 136928 79960
rect 137324 79908 137330 79960
rect 137382 79908 137388 79960
rect 136404 79840 136410 79892
rect 136462 79840 136468 79892
rect 136496 79840 136502 79892
rect 136554 79840 136560 79892
rect 136514 79756 136542 79840
rect 136450 79704 136456 79756
rect 136508 79716 136542 79756
rect 136508 79704 136514 79716
rect 136174 79500 136180 79552
rect 136232 79500 136238 79552
rect 135990 79432 135996 79484
rect 136048 79432 136054 79484
rect 136450 79432 136456 79484
rect 136508 79472 136514 79484
rect 136606 79472 136634 79908
rect 136882 79824 136910 79908
rect 137048 79840 137054 79892
rect 137106 79880 137112 79892
rect 137342 79880 137370 79908
rect 137480 79892 137508 80056
rect 137710 80016 137738 80328
rect 138630 80084 138658 80396
rect 138630 80056 140498 80084
rect 137710 79988 138566 80016
rect 138538 79960 138566 79988
rect 138630 79988 139026 80016
rect 137600 79908 137606 79960
rect 137658 79908 137664 79960
rect 137968 79908 137974 79960
rect 138026 79908 138032 79960
rect 138060 79908 138066 79960
rect 138118 79908 138124 79960
rect 138520 79908 138526 79960
rect 138578 79908 138584 79960
rect 137106 79840 137140 79880
rect 136882 79784 136916 79824
rect 136910 79772 136916 79784
rect 136968 79772 136974 79824
rect 137112 79756 137140 79840
rect 137204 79852 137370 79880
rect 137094 79704 137100 79756
rect 137152 79704 137158 79756
rect 137002 79636 137008 79688
rect 137060 79676 137066 79688
rect 137204 79676 137232 79852
rect 137416 79840 137422 79892
rect 137474 79852 137508 79892
rect 137474 79840 137480 79852
rect 137618 79688 137646 79908
rect 137986 79756 138014 79908
rect 137922 79704 137928 79756
rect 137980 79716 138014 79756
rect 137980 79704 137986 79716
rect 137060 79648 137232 79676
rect 137060 79636 137066 79648
rect 137554 79636 137560 79688
rect 137612 79648 137646 79688
rect 138078 79688 138106 79908
rect 138244 79840 138250 79892
rect 138302 79840 138308 79892
rect 138078 79648 138112 79688
rect 137612 79636 137618 79648
rect 138106 79636 138112 79648
rect 138164 79636 138170 79688
rect 137830 79500 137836 79552
rect 137888 79540 137894 79552
rect 138262 79540 138290 79840
rect 138630 79620 138658 79988
rect 138998 79960 139026 79988
rect 140470 79960 140498 80056
rect 141436 80016 141464 80464
rect 141528 80084 141556 80532
rect 141620 80152 141648 80600
rect 142126 80260 144730 80288
rect 142126 80152 142154 80260
rect 141620 80124 142154 80152
rect 143414 80192 144362 80220
rect 143414 80084 143442 80192
rect 141528 80056 143442 80084
rect 141436 79988 143626 80016
rect 138888 79948 138894 79960
rect 138566 79568 138572 79620
rect 138624 79580 138658 79620
rect 138768 79920 138894 79948
rect 138624 79568 138630 79580
rect 137888 79512 138290 79540
rect 137888 79500 137894 79512
rect 136508 79444 136634 79472
rect 136508 79432 136514 79444
rect 138382 79432 138388 79484
rect 138440 79472 138446 79484
rect 138768 79472 138796 79920
rect 138888 79908 138894 79920
rect 138946 79908 138952 79960
rect 138980 79908 138986 79960
rect 139038 79908 139044 79960
rect 139164 79908 139170 79960
rect 139222 79908 139228 79960
rect 139256 79908 139262 79960
rect 139314 79908 139320 79960
rect 139716 79948 139722 79960
rect 139458 79920 139722 79948
rect 139182 79812 139210 79908
rect 138998 79784 139210 79812
rect 138998 79552 139026 79784
rect 139274 79744 139302 79908
rect 139136 79716 139302 79744
rect 139136 79688 139164 79716
rect 139118 79636 139124 79688
rect 139176 79636 139182 79688
rect 139458 79676 139486 79920
rect 139716 79908 139722 79920
rect 139774 79908 139780 79960
rect 139808 79908 139814 79960
rect 139866 79948 139872 79960
rect 139866 79920 139946 79948
rect 139866 79908 139872 79920
rect 139762 79704 139768 79756
rect 139820 79744 139826 79756
rect 139918 79744 139946 79920
rect 139992 79908 139998 79960
rect 140050 79948 140056 79960
rect 140050 79920 140406 79948
rect 140050 79908 140056 79920
rect 140084 79840 140090 79892
rect 140142 79840 140148 79892
rect 140268 79880 140274 79892
rect 140240 79840 140274 79880
rect 140326 79840 140332 79892
rect 139820 79716 139946 79744
rect 139820 79704 139826 79716
rect 139274 79648 139486 79676
rect 138998 79512 139032 79552
rect 139026 79500 139032 79512
rect 139084 79500 139090 79552
rect 138440 79444 138796 79472
rect 139274 79484 139302 79648
rect 139946 79636 139952 79688
rect 140004 79676 140010 79688
rect 140102 79676 140130 79840
rect 140004 79648 140130 79676
rect 140004 79636 140010 79648
rect 139394 79568 139400 79620
rect 139452 79568 139458 79620
rect 139274 79444 139308 79484
rect 138440 79432 138446 79444
rect 139302 79432 139308 79444
rect 139360 79432 139366 79484
rect 139412 79472 139440 79568
rect 139670 79500 139676 79552
rect 139728 79540 139734 79552
rect 140240 79540 140268 79840
rect 140378 79812 140406 79920
rect 140452 79908 140458 79960
rect 140510 79908 140516 79960
rect 140544 79908 140550 79960
rect 140602 79908 140608 79960
rect 140636 79908 140642 79960
rect 140694 79908 140700 79960
rect 140820 79948 140826 79960
rect 140792 79908 140826 79948
rect 140878 79908 140884 79960
rect 141556 79948 141562 79960
rect 141160 79920 141562 79948
rect 140332 79784 140406 79812
rect 140332 79756 140360 79784
rect 140314 79704 140320 79756
rect 140372 79704 140378 79756
rect 140406 79704 140412 79756
rect 140464 79744 140470 79756
rect 140562 79744 140590 79908
rect 140464 79716 140590 79744
rect 140464 79704 140470 79716
rect 140654 79688 140682 79908
rect 140654 79648 140688 79688
rect 140682 79636 140688 79648
rect 140740 79636 140746 79688
rect 140792 79608 140820 79908
rect 141004 79880 141010 79892
rect 140884 79852 141010 79880
rect 140884 79620 140912 79852
rect 141004 79840 141010 79852
rect 141062 79840 141068 79892
rect 139728 79512 139992 79540
rect 139728 79500 139734 79512
rect 139854 79472 139860 79484
rect 139412 79444 139860 79472
rect 139854 79432 139860 79444
rect 139912 79432 139918 79484
rect 139964 79472 139992 79512
rect 140102 79512 140268 79540
rect 140332 79580 140820 79608
rect 140102 79472 140130 79512
rect 139964 79444 140130 79472
rect 140222 79432 140228 79484
rect 140280 79472 140286 79484
rect 140332 79472 140360 79580
rect 140866 79568 140872 79620
rect 140924 79568 140930 79620
rect 141160 79552 141188 79920
rect 141556 79908 141562 79920
rect 141614 79908 141620 79960
rect 141740 79908 141746 79960
rect 141798 79908 141804 79960
rect 141832 79908 141838 79960
rect 141890 79908 141896 79960
rect 141924 79908 141930 79960
rect 141982 79908 141988 79960
rect 142200 79908 142206 79960
rect 142258 79908 142264 79960
rect 143120 79948 143126 79960
rect 142954 79920 143126 79948
rect 141280 79880 141286 79892
rect 141252 79840 141286 79880
rect 141338 79840 141344 79892
rect 141252 79552 141280 79840
rect 141758 79812 141786 79908
rect 141620 79784 141786 79812
rect 141620 79688 141648 79784
rect 141850 79744 141878 79908
rect 141712 79716 141878 79744
rect 141602 79636 141608 79688
rect 141660 79636 141666 79688
rect 141712 79620 141740 79716
rect 141942 79676 141970 79908
rect 142108 79840 142114 79892
rect 142166 79840 142172 79892
rect 142126 79744 142154 79840
rect 142218 79812 142246 79908
rect 142476 79840 142482 79892
rect 142534 79840 142540 79892
rect 142568 79840 142574 79892
rect 142626 79840 142632 79892
rect 142218 79784 142384 79812
rect 142126 79716 142292 79744
rect 142264 79688 142292 79716
rect 141804 79648 141970 79676
rect 141694 79568 141700 79620
rect 141752 79568 141758 79620
rect 141804 79552 141832 79648
rect 142246 79636 142252 79688
rect 142304 79636 142310 79688
rect 142154 79568 142160 79620
rect 142212 79608 142218 79620
rect 142356 79608 142384 79784
rect 142494 79676 142522 79840
rect 142586 79756 142614 79840
rect 142586 79716 142620 79756
rect 142614 79704 142620 79716
rect 142672 79704 142678 79756
rect 142494 79648 142752 79676
rect 142212 79580 142384 79608
rect 142212 79568 142218 79580
rect 141142 79500 141148 79552
rect 141200 79500 141206 79552
rect 141234 79500 141240 79552
rect 141292 79500 141298 79552
rect 141786 79500 141792 79552
rect 141844 79500 141850 79552
rect 142724 79540 142752 79648
rect 142724 79512 142844 79540
rect 140280 79444 140360 79472
rect 140280 79432 140286 79444
rect 140590 79432 140596 79484
rect 140648 79472 140654 79484
rect 141418 79472 141424 79484
rect 140648 79444 141424 79472
rect 140648 79432 140654 79444
rect 141418 79432 141424 79444
rect 141476 79432 141482 79484
rect 141510 79432 141516 79484
rect 141568 79472 141574 79484
rect 142522 79472 142528 79484
rect 141568 79444 142528 79472
rect 141568 79432 141574 79444
rect 142522 79432 142528 79444
rect 142580 79432 142586 79484
rect 142816 79416 142844 79512
rect 142954 79416 142982 79920
rect 143120 79908 143126 79920
rect 143178 79908 143184 79960
rect 143212 79908 143218 79960
rect 143270 79908 143276 79960
rect 143396 79908 143402 79960
rect 143454 79908 143460 79960
rect 143488 79908 143494 79960
rect 143546 79908 143552 79960
rect 143230 79880 143258 79908
rect 143092 79852 143258 79880
rect 143092 79620 143120 79852
rect 143414 79812 143442 79908
rect 143184 79784 143442 79812
rect 143184 79676 143212 79784
rect 143258 79704 143264 79756
rect 143316 79744 143322 79756
rect 143506 79744 143534 79908
rect 143598 79812 143626 79988
rect 143736 79920 143994 79948
rect 143598 79784 143672 79812
rect 143316 79716 143534 79744
rect 143316 79704 143322 79716
rect 143350 79676 143356 79688
rect 143184 79648 143356 79676
rect 143350 79636 143356 79648
rect 143408 79636 143414 79688
rect 143074 79568 143080 79620
rect 143132 79568 143138 79620
rect 143644 79552 143672 79784
rect 143626 79500 143632 79552
rect 143684 79500 143690 79552
rect 143736 79540 143764 79920
rect 143966 79892 143994 79920
rect 144334 79892 144362 80192
rect 144408 79908 144414 79960
rect 144466 79908 144472 79960
rect 144500 79908 144506 79960
rect 144558 79908 144564 79960
rect 143856 79840 143862 79892
rect 143914 79840 143920 79892
rect 143948 79840 143954 79892
rect 144006 79840 144012 79892
rect 144132 79880 144138 79892
rect 144104 79840 144138 79880
rect 144190 79840 144196 79892
rect 144316 79840 144322 79892
rect 144374 79840 144380 79892
rect 143874 79676 143902 79840
rect 144104 79756 144132 79840
rect 144086 79704 144092 79756
rect 144144 79704 144150 79756
rect 144178 79676 144184 79688
rect 143874 79648 144184 79676
rect 144178 79636 144184 79648
rect 144236 79636 144242 79688
rect 143810 79568 143816 79620
rect 143868 79608 143874 79620
rect 144334 79608 144362 79840
rect 144426 79824 144454 79908
rect 144408 79772 144414 79824
rect 144466 79772 144472 79824
rect 144518 79688 144546 79908
rect 144702 79892 144730 80260
rect 144868 79908 144874 79960
rect 144926 79908 144932 79960
rect 145144 79948 145150 79960
rect 145116 79908 145150 79948
rect 145202 79908 145208 79960
rect 145236 79908 145242 79960
rect 145294 79908 145300 79960
rect 145328 79908 145334 79960
rect 145386 79948 145392 79960
rect 145386 79908 145420 79948
rect 144592 79840 144598 79892
rect 144650 79840 144656 79892
rect 144684 79840 144690 79892
rect 144742 79840 144748 79892
rect 144454 79636 144460 79688
rect 144512 79648 144546 79688
rect 144512 79636 144518 79648
rect 143868 79580 144362 79608
rect 143868 79568 143874 79580
rect 143902 79540 143908 79552
rect 143736 79512 143908 79540
rect 143902 79500 143908 79512
rect 143960 79500 143966 79552
rect 143644 79472 143672 79500
rect 144610 79472 144638 79840
rect 143644 79444 144638 79472
rect 135496 79376 135714 79404
rect 135496 79364 135502 79376
rect 136910 79364 136916 79416
rect 136968 79404 136974 79416
rect 142706 79404 142712 79416
rect 136968 79376 142712 79404
rect 136968 79364 136974 79376
rect 142706 79364 142712 79376
rect 142764 79364 142770 79416
rect 142798 79364 142804 79416
rect 142856 79364 142862 79416
rect 142890 79364 142896 79416
rect 142948 79376 142982 79416
rect 142948 79364 142954 79376
rect 144546 79364 144552 79416
rect 144604 79404 144610 79416
rect 144886 79404 144914 79908
rect 144604 79376 144914 79404
rect 145116 79404 145144 79908
rect 145254 79880 145282 79908
rect 145208 79852 145282 79880
rect 145208 79756 145236 79852
rect 145190 79704 145196 79756
rect 145248 79704 145254 79756
rect 145392 79688 145420 79908
rect 145374 79636 145380 79688
rect 145432 79636 145438 79688
rect 145484 79484 145512 80668
rect 145622 79960 145650 80736
rect 146634 80016 146662 80804
rect 161446 80804 174722 80832
rect 161446 80560 161474 80804
rect 174694 80764 174722 80804
rect 178236 80804 205088 80832
rect 174694 80736 178172 80764
rect 155926 80532 161474 80560
rect 161722 80668 173204 80696
rect 146634 79988 147352 80016
rect 146634 79960 146662 79988
rect 145604 79908 145610 79960
rect 145662 79948 145668 79960
rect 145662 79908 145696 79948
rect 145880 79908 145886 79960
rect 145938 79908 145944 79960
rect 145972 79908 145978 79960
rect 146030 79908 146036 79960
rect 146340 79948 146346 79960
rect 146312 79908 146346 79948
rect 146398 79908 146404 79960
rect 146432 79908 146438 79960
rect 146490 79908 146496 79960
rect 146616 79908 146622 79960
rect 146674 79908 146680 79960
rect 146708 79908 146714 79960
rect 146766 79908 146772 79960
rect 146800 79908 146806 79960
rect 146858 79908 146864 79960
rect 146984 79908 146990 79960
rect 147042 79908 147048 79960
rect 147076 79908 147082 79960
rect 147134 79908 147140 79960
rect 147168 79908 147174 79960
rect 147226 79948 147232 79960
rect 147226 79908 147260 79948
rect 145668 79552 145696 79908
rect 145788 79880 145794 79892
rect 145760 79840 145794 79880
rect 145846 79840 145852 79892
rect 145650 79500 145656 79552
rect 145708 79500 145714 79552
rect 145466 79432 145472 79484
rect 145524 79472 145530 79484
rect 145760 79472 145788 79840
rect 145898 79756 145926 79908
rect 145834 79704 145840 79756
rect 145892 79716 145926 79756
rect 145892 79704 145898 79716
rect 145990 79688 146018 79908
rect 146064 79840 146070 79892
rect 146122 79840 146128 79892
rect 146156 79840 146162 79892
rect 146214 79880 146220 79892
rect 146214 79840 146248 79880
rect 146082 79812 146110 79840
rect 146082 79784 146156 79812
rect 146128 79756 146156 79784
rect 146110 79704 146116 79756
rect 146168 79704 146174 79756
rect 146220 79688 146248 79840
rect 145926 79636 145932 79688
rect 145984 79648 146018 79688
rect 145984 79636 145990 79648
rect 146202 79636 146208 79688
rect 146260 79636 146266 79688
rect 146312 79620 146340 79908
rect 146450 79620 146478 79908
rect 146524 79840 146530 79892
rect 146582 79840 146588 79892
rect 146542 79688 146570 79840
rect 146726 79688 146754 79908
rect 146542 79648 146576 79688
rect 146570 79636 146576 79648
rect 146628 79636 146634 79688
rect 146662 79636 146668 79688
rect 146720 79648 146754 79688
rect 146720 79636 146726 79648
rect 146294 79568 146300 79620
rect 146352 79568 146358 79620
rect 146386 79568 146392 79620
rect 146444 79580 146478 79620
rect 146444 79568 146450 79580
rect 146818 79552 146846 79908
rect 146892 79772 146898 79824
rect 146950 79772 146956 79824
rect 146754 79500 146760 79552
rect 146812 79512 146846 79552
rect 146812 79500 146818 79512
rect 146910 79484 146938 79772
rect 145524 79444 145788 79472
rect 145524 79432 145530 79444
rect 146846 79432 146852 79484
rect 146904 79444 146938 79484
rect 146904 79432 146910 79444
rect 147002 79416 147030 79908
rect 147094 79744 147122 79908
rect 147094 79716 147168 79744
rect 147140 79540 147168 79716
rect 147232 79620 147260 79908
rect 147324 79676 147352 79988
rect 152154 79988 154528 80016
rect 152154 79960 152182 79988
rect 148088 79948 148094 79960
rect 148060 79908 148094 79948
rect 148146 79908 148152 79960
rect 149100 79908 149106 79960
rect 149158 79908 149164 79960
rect 149284 79908 149290 79960
rect 149342 79908 149348 79960
rect 149468 79908 149474 79960
rect 149526 79908 149532 79960
rect 149560 79908 149566 79960
rect 149618 79908 149624 79960
rect 149836 79908 149842 79960
rect 149894 79908 149900 79960
rect 150020 79908 150026 79960
rect 150078 79908 150084 79960
rect 150112 79908 150118 79960
rect 150170 79908 150176 79960
rect 150664 79908 150670 79960
rect 150722 79908 150728 79960
rect 150756 79908 150762 79960
rect 150814 79948 150820 79960
rect 151400 79948 151406 79960
rect 150814 79920 151032 79948
rect 150814 79908 150820 79920
rect 147536 79772 147542 79824
rect 147594 79812 147600 79824
rect 147594 79772 147628 79812
rect 147600 79688 147628 79772
rect 148060 79688 148088 79908
rect 148456 79840 148462 79892
rect 148514 79840 148520 79892
rect 148824 79840 148830 79892
rect 148882 79880 148888 79892
rect 148882 79852 149008 79880
rect 148882 79840 148888 79852
rect 148272 79772 148278 79824
rect 148330 79772 148336 79824
rect 147490 79676 147496 79688
rect 147324 79648 147496 79676
rect 147490 79636 147496 79648
rect 147548 79636 147554 79688
rect 147582 79636 147588 79688
rect 147640 79636 147646 79688
rect 148042 79636 148048 79688
rect 148100 79636 148106 79688
rect 148290 79620 148318 79772
rect 147214 79568 147220 79620
rect 147272 79568 147278 79620
rect 147858 79568 147864 79620
rect 147916 79568 147922 79620
rect 148226 79568 148232 79620
rect 148284 79580 148318 79620
rect 148284 79568 148290 79580
rect 147398 79540 147404 79552
rect 147140 79512 147404 79540
rect 147398 79500 147404 79512
rect 147456 79500 147462 79552
rect 147876 79540 147904 79568
rect 147876 79512 148410 79540
rect 145742 79404 145748 79416
rect 145116 79376 145748 79404
rect 144604 79364 144610 79376
rect 145742 79364 145748 79376
rect 145800 79364 145806 79416
rect 147002 79376 147036 79416
rect 147030 79364 147036 79376
rect 147088 79364 147094 79416
rect 148382 79404 148410 79512
rect 148474 79484 148502 79840
rect 148980 79620 149008 79852
rect 149118 79620 149146 79908
rect 149302 79880 149330 79908
rect 149302 79852 149376 79880
rect 149192 79772 149198 79824
rect 149250 79812 149256 79824
rect 149250 79772 149284 79812
rect 148962 79568 148968 79620
rect 149020 79568 149026 79620
rect 149118 79580 149152 79620
rect 149146 79568 149152 79580
rect 149204 79568 149210 79620
rect 149256 79552 149284 79772
rect 149238 79500 149244 79552
rect 149296 79500 149302 79552
rect 149348 79484 149376 79852
rect 149486 79824 149514 79908
rect 149578 79880 149606 79908
rect 149578 79852 149652 79880
rect 149486 79784 149520 79824
rect 149514 79772 149520 79784
rect 149572 79772 149578 79824
rect 149624 79484 149652 79852
rect 149854 79552 149882 79908
rect 150038 79756 150066 79908
rect 150130 79880 150158 79908
rect 150572 79880 150578 79892
rect 150130 79852 150204 79880
rect 150038 79716 150072 79756
rect 150066 79704 150072 79716
rect 150124 79704 150130 79756
rect 149790 79500 149796 79552
rect 149848 79512 149882 79552
rect 149848 79500 149854 79512
rect 148474 79444 148508 79484
rect 148502 79432 148508 79444
rect 148560 79432 148566 79484
rect 149330 79432 149336 79484
rect 149388 79432 149394 79484
rect 149606 79432 149612 79484
rect 149664 79432 149670 79484
rect 148870 79404 148876 79416
rect 148382 79376 148876 79404
rect 148870 79364 148876 79376
rect 148928 79364 148934 79416
rect 149422 79364 149428 79416
rect 149480 79404 149486 79416
rect 150176 79404 150204 79852
rect 150452 79852 150578 79880
rect 150452 79608 150480 79852
rect 150572 79840 150578 79852
rect 150630 79840 150636 79892
rect 150682 79812 150710 79908
rect 150544 79784 150710 79812
rect 150544 79688 150572 79784
rect 150526 79636 150532 79688
rect 150584 79636 150590 79688
rect 150802 79608 150808 79620
rect 150452 79580 150808 79608
rect 150802 79568 150808 79580
rect 150860 79568 150866 79620
rect 151004 79472 151032 79920
rect 151188 79920 151406 79948
rect 151078 79500 151084 79552
rect 151136 79540 151142 79552
rect 151188 79540 151216 79920
rect 151400 79908 151406 79920
rect 151458 79908 151464 79960
rect 152136 79908 152142 79960
rect 152194 79908 152200 79960
rect 152412 79908 152418 79960
rect 152470 79908 152476 79960
rect 152504 79908 152510 79960
rect 152562 79908 152568 79960
rect 153332 79908 153338 79960
rect 153390 79908 153396 79960
rect 153424 79908 153430 79960
rect 153482 79908 153488 79960
rect 153516 79908 153522 79960
rect 153574 79908 153580 79960
rect 153792 79908 153798 79960
rect 153850 79908 153856 79960
rect 154068 79908 154074 79960
rect 154126 79908 154132 79960
rect 154160 79908 154166 79960
rect 154218 79908 154224 79960
rect 154344 79908 154350 79960
rect 154402 79908 154408 79960
rect 151584 79880 151590 79892
rect 151464 79852 151590 79880
rect 151464 79552 151492 79852
rect 151584 79840 151590 79852
rect 151642 79840 151648 79892
rect 151952 79880 151958 79892
rect 151924 79840 151958 79880
rect 152010 79840 152016 79892
rect 152228 79840 152234 79892
rect 152286 79840 152292 79892
rect 151630 79744 151636 79756
rect 151556 79716 151636 79744
rect 151556 79620 151584 79716
rect 151630 79704 151636 79716
rect 151688 79704 151694 79756
rect 151538 79568 151544 79620
rect 151596 79568 151602 79620
rect 151924 79608 151952 79840
rect 152246 79688 152274 79840
rect 152430 79756 152458 79908
rect 152366 79704 152372 79756
rect 152424 79716 152458 79756
rect 152424 79704 152430 79716
rect 152522 79688 152550 79908
rect 152964 79840 152970 79892
rect 153022 79840 153028 79892
rect 153148 79840 153154 79892
rect 153206 79840 153212 79892
rect 153240 79840 153246 79892
rect 153298 79840 153304 79892
rect 152688 79772 152694 79824
rect 152746 79772 152752 79824
rect 152706 79688 152734 79772
rect 152182 79636 152188 79688
rect 152240 79648 152274 79688
rect 152240 79636 152246 79648
rect 152458 79636 152464 79688
rect 152516 79648 152550 79688
rect 152516 79636 152522 79648
rect 152642 79636 152648 79688
rect 152700 79648 152734 79688
rect 152700 79636 152706 79648
rect 151998 79608 152004 79620
rect 151924 79580 152004 79608
rect 151998 79568 152004 79580
rect 152056 79568 152062 79620
rect 152826 79568 152832 79620
rect 152884 79608 152890 79620
rect 152982 79608 153010 79840
rect 153166 79676 153194 79840
rect 152884 79580 153010 79608
rect 153120 79648 153194 79676
rect 152884 79568 152890 79580
rect 151136 79512 151216 79540
rect 151136 79500 151142 79512
rect 151446 79500 151452 79552
rect 151504 79500 151510 79552
rect 151354 79472 151360 79484
rect 151004 79444 151360 79472
rect 151354 79432 151360 79444
rect 151412 79432 151418 79484
rect 151814 79432 151820 79484
rect 151872 79472 151878 79484
rect 153120 79472 153148 79648
rect 153258 79608 153286 79840
rect 153350 79756 153378 79908
rect 153442 79812 153470 79908
rect 153534 79880 153562 79908
rect 153534 79852 153608 79880
rect 153442 79784 153516 79812
rect 153350 79716 153384 79756
rect 153378 79704 153384 79716
rect 153436 79704 153442 79756
rect 153488 79688 153516 79784
rect 153580 79688 153608 79852
rect 153810 79756 153838 79908
rect 153810 79716 153844 79756
rect 153838 79704 153844 79716
rect 153896 79704 153902 79756
rect 153470 79636 153476 79688
rect 153528 79636 153534 79688
rect 153562 79636 153568 79688
rect 153620 79636 153626 79688
rect 151872 79444 153148 79472
rect 153212 79580 153286 79608
rect 153212 79472 153240 79580
rect 153930 79568 153936 79620
rect 153988 79608 153994 79620
rect 154086 79608 154114 79908
rect 153988 79580 154114 79608
rect 153988 79568 153994 79580
rect 153746 79500 153752 79552
rect 153804 79540 153810 79552
rect 154178 79540 154206 79908
rect 154362 79756 154390 79908
rect 154298 79704 154304 79756
rect 154356 79716 154390 79756
rect 154356 79704 154362 79716
rect 154500 79688 154528 79988
rect 155926 79960 155954 80532
rect 161722 80152 161750 80668
rect 159606 80124 161750 80152
rect 161814 80600 168374 80628
rect 159606 79960 159634 80124
rect 161814 80084 161842 80600
rect 168346 80356 168374 80600
rect 173176 80424 173204 80668
rect 178144 80560 178172 80736
rect 178236 80640 178264 80804
rect 205082 80792 205088 80804
rect 205140 80792 205146 80844
rect 213178 80764 213184 80776
rect 178880 80736 213184 80764
rect 178218 80588 178224 80640
rect 178276 80588 178282 80640
rect 178880 80560 178908 80736
rect 213178 80724 213184 80736
rect 213236 80764 213242 80776
rect 302234 80764 302240 80776
rect 213236 80736 302240 80764
rect 213236 80724 213242 80736
rect 302234 80724 302240 80736
rect 302292 80724 302298 80776
rect 196710 80696 196716 80708
rect 178144 80532 178908 80560
rect 183296 80668 196716 80696
rect 177758 80452 177764 80504
rect 177816 80492 177822 80504
rect 183296 80492 183324 80668
rect 196710 80656 196716 80668
rect 196768 80696 196774 80708
rect 380894 80696 380900 80708
rect 196768 80668 380900 80696
rect 196768 80656 196774 80668
rect 380894 80656 380900 80668
rect 380952 80656 380958 80708
rect 192478 80628 192484 80640
rect 177816 80464 183324 80492
rect 183388 80600 192484 80628
rect 177816 80452 177822 80464
rect 183388 80424 183416 80600
rect 192478 80588 192484 80600
rect 192536 80588 192542 80640
rect 191006 80560 191012 80572
rect 173176 80396 183416 80424
rect 183526 80532 191012 80560
rect 177758 80356 177764 80368
rect 168346 80328 177764 80356
rect 177758 80316 177764 80328
rect 177816 80316 177822 80368
rect 178310 80316 178316 80368
rect 178368 80356 178374 80368
rect 183526 80356 183554 80532
rect 191006 80520 191012 80532
rect 191064 80520 191070 80572
rect 188338 80452 188344 80504
rect 188396 80492 188402 80504
rect 192386 80492 192392 80504
rect 188396 80464 192392 80492
rect 188396 80452 188402 80464
rect 192386 80452 192392 80464
rect 192444 80452 192450 80504
rect 188430 80384 188436 80436
rect 188488 80424 188494 80436
rect 195330 80424 195336 80436
rect 188488 80396 195336 80424
rect 188488 80384 188494 80396
rect 195330 80384 195336 80396
rect 195388 80384 195394 80436
rect 178368 80328 183554 80356
rect 178368 80316 178374 80328
rect 187050 80316 187056 80368
rect 187108 80356 187114 80368
rect 195146 80356 195152 80368
rect 187108 80328 195152 80356
rect 187108 80316 187114 80328
rect 195146 80316 195152 80328
rect 195204 80316 195210 80368
rect 178402 80288 178408 80300
rect 172578 80260 178408 80288
rect 172578 80220 172606 80260
rect 178402 80248 178408 80260
rect 178460 80248 178466 80300
rect 178126 80220 178132 80232
rect 170922 80192 172606 80220
rect 172762 80192 178132 80220
rect 161814 80056 162026 80084
rect 159974 79988 161520 80016
rect 159974 79960 160002 79988
rect 154620 79908 154626 79960
rect 154678 79908 154684 79960
rect 154988 79948 154994 79960
rect 154822 79920 154994 79948
rect 154482 79636 154488 79688
rect 154540 79636 154546 79688
rect 154638 79620 154666 79908
rect 154574 79568 154580 79620
rect 154632 79580 154666 79620
rect 154632 79568 154638 79580
rect 153804 79512 154206 79540
rect 153804 79500 153810 79512
rect 154206 79472 154212 79484
rect 153212 79444 154212 79472
rect 151872 79432 151878 79444
rect 154206 79432 154212 79444
rect 154264 79432 154270 79484
rect 149480 79376 150204 79404
rect 154822 79416 154850 79920
rect 154988 79908 154994 79920
rect 155046 79908 155052 79960
rect 155080 79908 155086 79960
rect 155138 79908 155144 79960
rect 155172 79908 155178 79960
rect 155230 79908 155236 79960
rect 155448 79908 155454 79960
rect 155506 79908 155512 79960
rect 155540 79908 155546 79960
rect 155598 79908 155604 79960
rect 155724 79908 155730 79960
rect 155782 79908 155788 79960
rect 155816 79908 155822 79960
rect 155874 79908 155880 79960
rect 155908 79908 155914 79960
rect 155966 79908 155972 79960
rect 158024 79908 158030 79960
rect 158082 79908 158088 79960
rect 158208 79948 158214 79960
rect 158134 79920 158214 79948
rect 154896 79840 154902 79892
rect 154954 79840 154960 79892
rect 154914 79472 154942 79840
rect 155098 79552 155126 79908
rect 155034 79500 155040 79552
rect 155092 79512 155126 79552
rect 155190 79552 155218 79908
rect 155466 79620 155494 79908
rect 155402 79568 155408 79620
rect 155460 79580 155494 79620
rect 155460 79568 155466 79580
rect 155558 79552 155586 79908
rect 155632 79772 155638 79824
rect 155690 79772 155696 79824
rect 155190 79512 155224 79552
rect 155092 79500 155098 79512
rect 155218 79500 155224 79512
rect 155276 79500 155282 79552
rect 155494 79500 155500 79552
rect 155552 79512 155586 79552
rect 155552 79500 155558 79512
rect 154914 79444 155172 79472
rect 155144 79416 155172 79444
rect 155310 79432 155316 79484
rect 155368 79472 155374 79484
rect 155650 79472 155678 79772
rect 155742 79608 155770 79908
rect 155834 79744 155862 79908
rect 156828 79840 156834 79892
rect 156886 79840 156892 79892
rect 156920 79840 156926 79892
rect 156978 79840 156984 79892
rect 157472 79840 157478 79892
rect 157530 79840 157536 79892
rect 157840 79840 157846 79892
rect 157898 79840 157904 79892
rect 156276 79772 156282 79824
rect 156334 79772 156340 79824
rect 155834 79716 156000 79744
rect 155742 79580 155908 79608
rect 155880 79552 155908 79580
rect 155862 79500 155868 79552
rect 155920 79500 155926 79552
rect 155368 79444 155678 79472
rect 155368 79432 155374 79444
rect 155770 79432 155776 79484
rect 155828 79472 155834 79484
rect 155972 79472 156000 79716
rect 156294 79540 156322 79772
rect 156846 79620 156874 79840
rect 156938 79756 156966 79840
rect 156938 79716 156972 79756
rect 156966 79704 156972 79716
rect 157024 79704 157030 79756
rect 156782 79568 156788 79620
rect 156840 79580 156874 79620
rect 156840 79568 156846 79580
rect 157490 79552 157518 79840
rect 157610 79568 157616 79620
rect 157668 79608 157674 79620
rect 157858 79608 157886 79840
rect 157668 79580 157886 79608
rect 157668 79568 157674 79580
rect 156690 79540 156696 79552
rect 156294 79512 156696 79540
rect 156690 79500 156696 79512
rect 156748 79500 156754 79552
rect 157426 79500 157432 79552
rect 157484 79512 157518 79552
rect 157484 79500 157490 79512
rect 155828 79444 156000 79472
rect 158042 79484 158070 79908
rect 158134 79620 158162 79920
rect 158208 79908 158214 79920
rect 158266 79908 158272 79960
rect 158300 79908 158306 79960
rect 158358 79908 158364 79960
rect 158484 79948 158490 79960
rect 158410 79920 158490 79948
rect 158318 79824 158346 79908
rect 158300 79772 158306 79824
rect 158358 79772 158364 79824
rect 158254 79636 158260 79688
rect 158312 79676 158318 79688
rect 158410 79676 158438 79920
rect 158484 79908 158490 79920
rect 158542 79908 158548 79960
rect 158576 79908 158582 79960
rect 158634 79908 158640 79960
rect 158668 79908 158674 79960
rect 158726 79908 158732 79960
rect 159128 79948 159134 79960
rect 158824 79920 159134 79948
rect 158594 79880 158622 79908
rect 158312 79648 158438 79676
rect 158548 79852 158622 79880
rect 158312 79636 158318 79648
rect 158548 79620 158576 79852
rect 158686 79824 158714 79908
rect 158622 79772 158628 79824
rect 158680 79784 158714 79824
rect 158680 79772 158686 79784
rect 158824 79688 158852 79920
rect 159128 79908 159134 79920
rect 159186 79908 159192 79960
rect 159220 79908 159226 79960
rect 159278 79908 159284 79960
rect 159312 79908 159318 79960
rect 159370 79908 159376 79960
rect 159496 79908 159502 79960
rect 159554 79908 159560 79960
rect 159588 79908 159594 79960
rect 159646 79908 159652 79960
rect 159956 79908 159962 79960
rect 160014 79908 160020 79960
rect 160140 79908 160146 79960
rect 160198 79908 160204 79960
rect 160508 79948 160514 79960
rect 160480 79908 160514 79948
rect 160566 79908 160572 79960
rect 159238 79824 159266 79908
rect 158944 79772 158950 79824
rect 159002 79772 159008 79824
rect 159036 79772 159042 79824
rect 159094 79772 159100 79824
rect 159174 79772 159180 79824
rect 159232 79784 159266 79824
rect 159232 79772 159238 79784
rect 158714 79636 158720 79688
rect 158772 79636 158778 79688
rect 158806 79636 158812 79688
rect 158864 79636 158870 79688
rect 158134 79580 158168 79620
rect 158162 79568 158168 79580
rect 158220 79568 158226 79620
rect 158530 79568 158536 79620
rect 158588 79568 158594 79620
rect 158732 79608 158760 79636
rect 158962 79620 158990 79772
rect 158640 79580 158760 79608
rect 158042 79444 158076 79484
rect 155828 79432 155834 79444
rect 158070 79432 158076 79444
rect 158128 79432 158134 79484
rect 158640 79472 158668 79580
rect 158898 79568 158904 79620
rect 158956 79580 158990 79620
rect 158956 79568 158962 79580
rect 158898 79472 158904 79484
rect 158640 79444 158904 79472
rect 158898 79432 158904 79444
rect 158956 79432 158962 79484
rect 154822 79376 154856 79416
rect 149480 79364 149486 79376
rect 154850 79364 154856 79376
rect 154908 79364 154914 79416
rect 155126 79364 155132 79416
rect 155184 79364 155190 79416
rect 159054 79404 159082 79772
rect 159330 79756 159358 79908
rect 159266 79704 159272 79756
rect 159324 79716 159358 79756
rect 159514 79756 159542 79908
rect 159772 79772 159778 79824
rect 159830 79772 159836 79824
rect 159514 79716 159548 79756
rect 159324 79704 159330 79716
rect 159542 79704 159548 79716
rect 159600 79704 159606 79756
rect 159790 79688 159818 79772
rect 160158 79688 160186 79908
rect 160480 79824 160508 79908
rect 160600 79880 160606 79892
rect 160572 79840 160606 79880
rect 160658 79840 160664 79892
rect 160784 79840 160790 79892
rect 160842 79840 160848 79892
rect 161060 79880 161066 79892
rect 161032 79840 161066 79880
rect 161118 79840 161124 79892
rect 161336 79880 161342 79892
rect 161216 79852 161342 79880
rect 160462 79772 160468 79824
rect 160520 79772 160526 79824
rect 160572 79756 160600 79840
rect 160554 79704 160560 79756
rect 160612 79704 160618 79756
rect 159790 79648 159824 79688
rect 159818 79636 159824 79648
rect 159876 79636 159882 79688
rect 160094 79636 160100 79688
rect 160152 79648 160186 79688
rect 160152 79636 160158 79648
rect 160802 79416 160830 79840
rect 161032 79620 161060 79840
rect 161216 79620 161244 79852
rect 161336 79840 161342 79852
rect 161394 79840 161400 79892
rect 161492 79620 161520 79988
rect 161998 79960 162026 80056
rect 166184 79988 166534 80016
rect 161980 79908 161986 79960
rect 162038 79908 162044 79960
rect 162072 79908 162078 79960
rect 162130 79908 162136 79960
rect 162164 79908 162170 79960
rect 162222 79908 162228 79960
rect 162348 79908 162354 79960
rect 162406 79908 162412 79960
rect 162440 79908 162446 79960
rect 162498 79908 162504 79960
rect 162532 79908 162538 79960
rect 162590 79908 162596 79960
rect 162716 79908 162722 79960
rect 162774 79908 162780 79960
rect 163084 79908 163090 79960
rect 163142 79908 163148 79960
rect 163268 79908 163274 79960
rect 163326 79908 163332 79960
rect 163360 79908 163366 79960
rect 163418 79908 163424 79960
rect 163452 79908 163458 79960
rect 163510 79948 163516 79960
rect 163510 79920 163636 79948
rect 163510 79908 163516 79920
rect 161612 79840 161618 79892
rect 161670 79840 161676 79892
rect 161704 79840 161710 79892
rect 161762 79880 161768 79892
rect 161762 79852 161980 79880
rect 161762 79840 161768 79852
rect 161630 79812 161658 79840
rect 161630 79784 161888 79812
rect 161014 79568 161020 79620
rect 161072 79568 161078 79620
rect 161198 79568 161204 79620
rect 161256 79568 161262 79620
rect 161474 79568 161480 79620
rect 161532 79568 161538 79620
rect 161860 79552 161888 79784
rect 161842 79500 161848 79552
rect 161900 79500 161906 79552
rect 161952 79540 161980 79852
rect 162090 79824 162118 79908
rect 162026 79772 162032 79824
rect 162084 79784 162118 79824
rect 162084 79772 162090 79784
rect 162182 79756 162210 79908
rect 162366 79824 162394 79908
rect 162458 79824 162486 79908
rect 162302 79772 162308 79824
rect 162360 79784 162394 79824
rect 162360 79772 162366 79784
rect 162440 79772 162446 79824
rect 162498 79772 162504 79824
rect 162118 79704 162124 79756
rect 162176 79716 162210 79756
rect 162550 79744 162578 79908
rect 162504 79716 162578 79744
rect 162176 79704 162182 79716
rect 162504 79688 162532 79716
rect 162486 79636 162492 79688
rect 162544 79636 162550 79688
rect 162734 79620 162762 79908
rect 162992 79772 162998 79824
rect 163050 79772 163056 79824
rect 162670 79568 162676 79620
rect 162728 79580 162762 79620
rect 163010 79620 163038 79772
rect 163102 79688 163130 79908
rect 163286 79744 163314 79908
rect 163240 79716 163314 79744
rect 163240 79688 163268 79716
rect 163378 79688 163406 79908
rect 163102 79648 163136 79688
rect 163130 79636 163136 79648
rect 163188 79636 163194 79688
rect 163222 79636 163228 79688
rect 163280 79636 163286 79688
rect 163314 79636 163320 79688
rect 163372 79648 163406 79688
rect 163372 79636 163378 79648
rect 163010 79580 163044 79620
rect 162728 79568 162734 79580
rect 163038 79568 163044 79580
rect 163096 79568 163102 79620
rect 162486 79540 162492 79552
rect 161952 79512 162492 79540
rect 162486 79500 162492 79512
rect 162544 79500 162550 79552
rect 162854 79500 162860 79552
rect 162912 79540 162918 79552
rect 163608 79540 163636 79920
rect 164372 79908 164378 79960
rect 164430 79908 164436 79960
rect 164556 79908 164562 79960
rect 164614 79908 164620 79960
rect 165016 79908 165022 79960
rect 165074 79908 165080 79960
rect 165568 79948 165574 79960
rect 165540 79908 165574 79948
rect 165626 79908 165632 79960
rect 165752 79908 165758 79960
rect 165810 79908 165816 79960
rect 165936 79908 165942 79960
rect 165994 79908 166000 79960
rect 166028 79908 166034 79960
rect 166086 79908 166092 79960
rect 163728 79840 163734 79892
rect 163786 79840 163792 79892
rect 163746 79608 163774 79840
rect 164096 79772 164102 79824
rect 164154 79772 164160 79824
rect 164114 79676 164142 79772
rect 164390 79744 164418 79908
rect 164574 79812 164602 79908
rect 164648 79840 164654 79892
rect 164706 79880 164712 79892
rect 164706 79852 164924 79880
rect 164706 79840 164712 79852
rect 164574 79784 164648 79812
rect 164620 79756 164648 79784
rect 164510 79744 164516 79756
rect 164390 79716 164516 79744
rect 164510 79704 164516 79716
rect 164568 79704 164574 79756
rect 164602 79704 164608 79756
rect 164660 79704 164666 79756
rect 164896 79688 164924 79852
rect 164326 79676 164332 79688
rect 164114 79648 164332 79676
rect 164326 79636 164332 79648
rect 164384 79636 164390 79688
rect 164878 79636 164884 79688
rect 164936 79636 164942 79688
rect 164050 79608 164056 79620
rect 163746 79580 164056 79608
rect 164050 79568 164056 79580
rect 164108 79568 164114 79620
rect 162912 79512 163636 79540
rect 162912 79500 162918 79512
rect 161934 79432 161940 79484
rect 161992 79472 161998 79484
rect 161992 79444 162854 79472
rect 161992 79432 161998 79444
rect 159542 79404 159548 79416
rect 159054 79376 159548 79404
rect 159542 79364 159548 79376
rect 159600 79364 159606 79416
rect 160738 79364 160744 79416
rect 160796 79376 160830 79416
rect 160796 79364 160802 79376
rect 143166 79336 143172 79348
rect 132420 79308 143172 79336
rect 143166 79296 143172 79308
rect 143224 79296 143230 79348
rect 162826 79336 162854 79444
rect 164418 79364 164424 79416
rect 164476 79404 164482 79416
rect 165034 79404 165062 79908
rect 165200 79840 165206 79892
rect 165258 79840 165264 79892
rect 165218 79540 165246 79840
rect 165292 79772 165298 79824
rect 165350 79772 165356 79824
rect 165384 79772 165390 79824
rect 165442 79812 165448 79824
rect 165442 79772 165476 79812
rect 165310 79620 165338 79772
rect 165448 79688 165476 79772
rect 165540 79688 165568 79908
rect 165770 79756 165798 79908
rect 165770 79716 165804 79756
rect 165798 79704 165804 79716
rect 165856 79704 165862 79756
rect 165430 79636 165436 79688
rect 165488 79636 165494 79688
rect 165522 79636 165528 79688
rect 165580 79636 165586 79688
rect 165310 79580 165344 79620
rect 165338 79568 165344 79580
rect 165396 79568 165402 79620
rect 165954 79608 165982 79908
rect 166046 79824 166074 79908
rect 166028 79772 166034 79824
rect 166086 79772 166092 79824
rect 166184 79620 166212 79988
rect 166506 79960 166534 79988
rect 166966 79988 167546 80016
rect 166304 79908 166310 79960
rect 166362 79908 166368 79960
rect 166396 79908 166402 79960
rect 166454 79908 166460 79960
rect 166488 79908 166494 79960
rect 166546 79908 166552 79960
rect 166856 79908 166862 79960
rect 166914 79908 166920 79960
rect 166322 79744 166350 79908
rect 166414 79880 166442 79908
rect 166414 79852 166672 79880
rect 166322 79716 166488 79744
rect 166460 79688 166488 79716
rect 166442 79636 166448 79688
rect 166500 79636 166506 79688
rect 166644 79620 166672 79852
rect 166874 79620 166902 79908
rect 166966 79688 166994 79988
rect 167518 79960 167546 79988
rect 170922 79960 170950 80192
rect 172762 80016 172790 80192
rect 178126 80180 178132 80192
rect 178184 80180 178190 80232
rect 191282 80180 191288 80232
rect 191340 80220 191346 80232
rect 191926 80220 191932 80232
rect 191340 80192 191932 80220
rect 191340 80180 191346 80192
rect 191926 80180 191932 80192
rect 191984 80180 191990 80232
rect 178034 80152 178040 80164
rect 175614 80124 178040 80152
rect 175614 80084 175642 80124
rect 178034 80112 178040 80124
rect 178092 80112 178098 80164
rect 178218 80084 178224 80096
rect 171290 79988 172790 80016
rect 172854 80056 175642 80084
rect 175706 80056 178224 80084
rect 171290 79960 171318 79988
rect 167040 79908 167046 79960
rect 167098 79948 167104 79960
rect 167098 79920 167316 79948
rect 167098 79908 167104 79920
rect 166966 79648 167000 79688
rect 166994 79636 167000 79648
rect 167052 79636 167058 79688
rect 166074 79608 166080 79620
rect 165954 79580 166080 79608
rect 166074 79568 166080 79580
rect 166132 79568 166138 79620
rect 166166 79568 166172 79620
rect 166224 79568 166230 79620
rect 166626 79568 166632 79620
rect 166684 79568 166690 79620
rect 166874 79580 166908 79620
rect 166902 79568 166908 79580
rect 166960 79568 166966 79620
rect 166350 79540 166356 79552
rect 165218 79512 166356 79540
rect 166350 79500 166356 79512
rect 166408 79500 166414 79552
rect 167086 79500 167092 79552
rect 167144 79500 167150 79552
rect 167288 79540 167316 79920
rect 167408 79908 167414 79960
rect 167466 79908 167472 79960
rect 167500 79908 167506 79960
rect 167558 79908 167564 79960
rect 168328 79908 168334 79960
rect 168386 79908 168392 79960
rect 168420 79908 168426 79960
rect 168478 79908 168484 79960
rect 168696 79908 168702 79960
rect 168754 79948 168760 79960
rect 168754 79908 168788 79948
rect 168972 79908 168978 79960
rect 169030 79908 169036 79960
rect 169064 79908 169070 79960
rect 169122 79908 169128 79960
rect 169156 79908 169162 79960
rect 169214 79948 169220 79960
rect 169524 79948 169530 79960
rect 169214 79920 169432 79948
rect 169214 79908 169220 79920
rect 167426 79676 167454 79908
rect 167960 79840 167966 79892
rect 168018 79840 168024 79892
rect 168144 79840 168150 79892
rect 168202 79880 168208 79892
rect 168202 79840 168236 79880
rect 167978 79744 168006 79840
rect 168098 79744 168104 79756
rect 167978 79716 168104 79744
rect 168098 79704 168104 79716
rect 168156 79704 168162 79756
rect 168208 79688 168236 79840
rect 168006 79676 168012 79688
rect 167426 79648 168012 79676
rect 168006 79636 168012 79648
rect 168064 79636 168070 79688
rect 168190 79636 168196 79688
rect 168248 79636 168254 79688
rect 167914 79540 167920 79552
rect 167288 79512 167920 79540
rect 167914 79500 167920 79512
rect 167972 79500 167978 79552
rect 167104 79472 167132 79500
rect 167546 79472 167552 79484
rect 167104 79444 167552 79472
rect 167546 79432 167552 79444
rect 167604 79432 167610 79484
rect 168346 79472 168374 79908
rect 168438 79620 168466 79908
rect 168512 79840 168518 79892
rect 168570 79840 168576 79892
rect 168530 79812 168558 79840
rect 168760 79824 168788 79908
rect 168880 79840 168886 79892
rect 168938 79840 168944 79892
rect 168650 79812 168656 79824
rect 168530 79784 168656 79812
rect 168650 79772 168656 79784
rect 168708 79772 168714 79824
rect 168742 79772 168748 79824
rect 168800 79772 168806 79824
rect 168898 79756 168926 79840
rect 168834 79704 168840 79756
rect 168892 79716 168926 79756
rect 168892 79704 168898 79716
rect 168438 79580 168472 79620
rect 168466 79568 168472 79580
rect 168524 79568 168530 79620
rect 168990 79608 169018 79908
rect 169082 79756 169110 79908
rect 169248 79880 169254 79892
rect 169220 79840 169254 79880
rect 169306 79840 169312 79892
rect 169220 79756 169248 79840
rect 169082 79716 169116 79756
rect 169110 79704 169116 79716
rect 169168 79704 169174 79756
rect 169202 79704 169208 79756
rect 169260 79704 169266 79756
rect 169404 79688 169432 79920
rect 169496 79908 169530 79948
rect 169582 79908 169588 79960
rect 170904 79948 170910 79960
rect 170370 79920 170910 79948
rect 169496 79756 169524 79908
rect 169708 79840 169714 79892
rect 169766 79840 169772 79892
rect 169478 79704 169484 79756
rect 169536 79704 169542 79756
rect 169386 79636 169392 79688
rect 169444 79636 169450 79688
rect 168990 79580 169064 79608
rect 168926 79472 168932 79484
rect 168346 79444 168932 79472
rect 164476 79376 165062 79404
rect 164476 79364 164482 79376
rect 167086 79364 167092 79416
rect 167144 79404 167150 79416
rect 168346 79404 168374 79444
rect 168926 79432 168932 79444
rect 168984 79432 168990 79484
rect 167144 79376 168374 79404
rect 169036 79404 169064 79580
rect 169570 79500 169576 79552
rect 169628 79540 169634 79552
rect 169726 79540 169754 79840
rect 169892 79812 169898 79824
rect 169818 79784 169898 79812
rect 169818 79620 169846 79784
rect 169892 79772 169898 79784
rect 169950 79772 169956 79824
rect 169984 79772 169990 79824
rect 170042 79772 170048 79824
rect 170168 79812 170174 79824
rect 170140 79772 170174 79812
rect 170226 79772 170232 79824
rect 170260 79772 170266 79824
rect 170318 79772 170324 79824
rect 170002 79744 170030 79772
rect 170140 79744 170168 79772
rect 169956 79716 170030 79744
rect 170094 79716 170168 79744
rect 169956 79620 169984 79716
rect 170094 79688 170122 79716
rect 170030 79636 170036 79688
rect 170088 79648 170122 79688
rect 170088 79636 170094 79648
rect 169818 79580 169852 79620
rect 169846 79568 169852 79580
rect 169904 79568 169910 79620
rect 169938 79568 169944 79620
rect 169996 79568 170002 79620
rect 170122 79568 170128 79620
rect 170180 79608 170186 79620
rect 170278 79608 170306 79772
rect 170180 79580 170306 79608
rect 170180 79568 170186 79580
rect 169628 79512 169754 79540
rect 169628 79500 169634 79512
rect 169754 79432 169760 79484
rect 169812 79472 169818 79484
rect 170370 79472 170398 79920
rect 170904 79908 170910 79920
rect 170962 79908 170968 79960
rect 171272 79908 171278 79960
rect 171330 79908 171336 79960
rect 171364 79908 171370 79960
rect 171422 79908 171428 79960
rect 171548 79908 171554 79960
rect 171606 79908 171612 79960
rect 171640 79908 171646 79960
rect 171698 79908 171704 79960
rect 171824 79908 171830 79960
rect 171882 79908 171888 79960
rect 171916 79908 171922 79960
rect 171974 79948 171980 79960
rect 172100 79948 172106 79960
rect 171974 79908 172008 79948
rect 170720 79840 170726 79892
rect 170778 79840 170784 79892
rect 170812 79840 170818 79892
rect 170870 79840 170876 79892
rect 170738 79676 170766 79840
rect 170830 79744 170858 79840
rect 171382 79756 171410 79908
rect 171566 79756 171594 79908
rect 170830 79716 170996 79744
rect 171382 79716 171416 79756
rect 170858 79676 170864 79688
rect 170738 79648 170864 79676
rect 170858 79636 170864 79648
rect 170916 79636 170922 79688
rect 170674 79568 170680 79620
rect 170732 79608 170738 79620
rect 170968 79608 170996 79716
rect 171410 79704 171416 79716
rect 171468 79704 171474 79756
rect 171502 79704 171508 79756
rect 171560 79716 171594 79756
rect 171560 79704 171566 79716
rect 171658 79688 171686 79908
rect 171732 79840 171738 79892
rect 171790 79840 171796 79892
rect 171594 79636 171600 79688
rect 171652 79648 171686 79688
rect 171652 79636 171658 79648
rect 170732 79580 170996 79608
rect 170732 79568 170738 79580
rect 171226 79568 171232 79620
rect 171284 79608 171290 79620
rect 171750 79608 171778 79840
rect 171284 79580 171778 79608
rect 171842 79620 171870 79908
rect 171980 79688 172008 79908
rect 172072 79908 172106 79948
rect 172158 79908 172164 79960
rect 172284 79908 172290 79960
rect 172342 79908 172348 79960
rect 172652 79908 172658 79960
rect 172710 79948 172716 79960
rect 172854 79948 172882 80056
rect 173958 79988 174446 80016
rect 173958 79948 173986 79988
rect 172710 79920 172882 79948
rect 172946 79920 173986 79948
rect 172710 79908 172716 79920
rect 171962 79636 171968 79688
rect 172020 79636 172026 79688
rect 172072 79620 172100 79908
rect 172192 79880 172198 79892
rect 172164 79840 172198 79880
rect 172250 79840 172256 79892
rect 172164 79620 172192 79840
rect 172302 79756 172330 79908
rect 172744 79840 172750 79892
rect 172802 79880 172808 79892
rect 172946 79880 172974 79920
rect 174032 79908 174038 79960
rect 174090 79908 174096 79960
rect 172802 79852 172974 79880
rect 172802 79840 172808 79852
rect 173020 79840 173026 79892
rect 173078 79880 173084 79892
rect 173078 79852 173480 79880
rect 173078 79840 173084 79852
rect 172376 79772 172382 79824
rect 172434 79772 172440 79824
rect 172560 79772 172566 79824
rect 172618 79772 172624 79824
rect 173296 79772 173302 79824
rect 173354 79772 173360 79824
rect 172238 79704 172244 79756
rect 172296 79716 172330 79756
rect 172296 79704 172302 79716
rect 171842 79580 171876 79620
rect 171284 79568 171290 79580
rect 169812 79444 170398 79472
rect 171750 79472 171778 79580
rect 171870 79568 171876 79580
rect 171928 79568 171934 79620
rect 172054 79568 172060 79620
rect 172112 79568 172118 79620
rect 172146 79568 172152 79620
rect 172204 79568 172210 79620
rect 172394 79552 172422 79772
rect 172578 79688 172606 79772
rect 173314 79688 173342 79772
rect 172578 79648 172612 79688
rect 172606 79636 172612 79648
rect 172664 79636 172670 79688
rect 173314 79648 173348 79688
rect 173342 79636 173348 79648
rect 173400 79636 173406 79688
rect 172394 79512 172428 79552
rect 172422 79500 172428 79512
rect 172480 79500 172486 79552
rect 171750 79444 172514 79472
rect 169812 79432 169818 79444
rect 169294 79404 169300 79416
rect 169036 79376 169300 79404
rect 167144 79364 167150 79376
rect 169294 79364 169300 79376
rect 169352 79364 169358 79416
rect 171134 79364 171140 79416
rect 171192 79404 171198 79416
rect 171778 79404 171784 79416
rect 171192 79376 171784 79404
rect 171192 79364 171198 79376
rect 171778 79364 171784 79376
rect 171836 79364 171842 79416
rect 172486 79404 172514 79444
rect 172882 79404 172888 79416
rect 172486 79376 172888 79404
rect 172882 79364 172888 79376
rect 172940 79364 172946 79416
rect 172974 79364 172980 79416
rect 173032 79404 173038 79416
rect 173250 79404 173256 79416
rect 173032 79376 173256 79404
rect 173032 79364 173038 79376
rect 173250 79364 173256 79376
rect 173308 79364 173314 79416
rect 173066 79336 173072 79348
rect 162826 79308 173072 79336
rect 173066 79296 173072 79308
rect 173124 79296 173130 79348
rect 96080 79132 96108 79296
rect 111334 79228 111340 79280
rect 111392 79268 111398 79280
rect 145006 79268 145012 79280
rect 111392 79240 145012 79268
rect 111392 79228 111398 79240
rect 145006 79228 145012 79240
rect 145064 79228 145070 79280
rect 147858 79228 147864 79280
rect 147916 79268 147922 79280
rect 172974 79268 172980 79280
rect 147916 79240 172980 79268
rect 147916 79228 147922 79240
rect 172974 79228 172980 79240
rect 173032 79228 173038 79280
rect 173452 79268 173480 79852
rect 173940 79772 173946 79824
rect 173998 79772 174004 79824
rect 173958 79688 173986 79772
rect 173894 79636 173900 79688
rect 173952 79648 173986 79688
rect 173952 79636 173958 79648
rect 174050 79608 174078 79908
rect 174216 79840 174222 79892
rect 174274 79880 174280 79892
rect 174274 79840 174308 79880
rect 174280 79688 174308 79840
rect 174262 79636 174268 79688
rect 174320 79636 174326 79688
rect 173866 79580 174078 79608
rect 174418 79608 174446 79988
rect 174492 79908 174498 79960
rect 174550 79908 174556 79960
rect 174584 79908 174590 79960
rect 174642 79908 174648 79960
rect 174676 79908 174682 79960
rect 174734 79948 174740 79960
rect 174734 79920 174906 79948
rect 174734 79908 174740 79920
rect 174510 79824 174538 79908
rect 174602 79880 174630 79908
rect 174602 79852 174768 79880
rect 174510 79784 174544 79824
rect 174538 79772 174544 79784
rect 174596 79772 174602 79824
rect 174740 79688 174768 79852
rect 174878 79744 174906 79920
rect 175320 79908 175326 79960
rect 175378 79948 175384 79960
rect 175706 79948 175734 80056
rect 178218 80044 178224 80056
rect 178276 80044 178282 80096
rect 186958 80044 186964 80096
rect 187016 80084 187022 80096
rect 190086 80084 190092 80096
rect 187016 80056 190092 80084
rect 187016 80044 187022 80056
rect 190086 80044 190092 80056
rect 190144 80044 190150 80096
rect 215846 80044 215852 80096
rect 215904 80084 215910 80096
rect 288434 80084 288440 80096
rect 215904 80056 288440 80084
rect 215904 80044 215910 80056
rect 288434 80044 288440 80056
rect 288492 80044 288498 80096
rect 178770 80016 178776 80028
rect 176350 79988 178776 80016
rect 176350 79960 176378 79988
rect 178770 79976 178776 79988
rect 178828 79976 178834 80028
rect 175378 79920 175734 79948
rect 175378 79908 175384 79920
rect 175872 79908 175878 79960
rect 175930 79908 175936 79960
rect 175964 79908 175970 79960
rect 176022 79908 176028 79960
rect 176148 79908 176154 79960
rect 176206 79908 176212 79960
rect 176332 79908 176338 79960
rect 176390 79908 176396 79960
rect 176424 79908 176430 79960
rect 176482 79908 176488 79960
rect 176884 79908 176890 79960
rect 176942 79908 176948 79960
rect 177068 79908 177074 79960
rect 177126 79948 177132 79960
rect 177758 79948 177764 79960
rect 177126 79920 177764 79948
rect 177126 79908 177132 79920
rect 177758 79908 177764 79920
rect 177816 79908 177822 79960
rect 174878 79716 175228 79744
rect 175200 79688 175228 79716
rect 175338 79688 175366 79908
rect 175688 79840 175694 79892
rect 175746 79840 175752 79892
rect 175504 79772 175510 79824
rect 175562 79772 175568 79824
rect 175522 79688 175550 79772
rect 174722 79636 174728 79688
rect 174780 79636 174786 79688
rect 175182 79636 175188 79688
rect 175240 79636 175246 79688
rect 175274 79636 175280 79688
rect 175332 79648 175366 79688
rect 175332 79636 175338 79648
rect 175458 79636 175464 79688
rect 175516 79648 175550 79688
rect 175706 79676 175734 79840
rect 175890 79756 175918 79908
rect 175826 79704 175832 79756
rect 175884 79716 175918 79756
rect 175982 79756 176010 79908
rect 176166 79756 176194 79908
rect 176442 79756 176470 79908
rect 176608 79840 176614 79892
rect 176666 79880 176672 79892
rect 176666 79840 176700 79880
rect 176792 79840 176798 79892
rect 176850 79840 176856 79892
rect 175982 79716 176016 79756
rect 175884 79704 175890 79716
rect 176010 79704 176016 79716
rect 176068 79704 176074 79756
rect 176166 79716 176200 79756
rect 176194 79704 176200 79716
rect 176252 79704 176258 79756
rect 176378 79704 176384 79756
rect 176436 79716 176470 79756
rect 176436 79704 176442 79716
rect 176286 79676 176292 79688
rect 175706 79648 176292 79676
rect 175516 79636 175522 79648
rect 176286 79636 176292 79648
rect 176344 79636 176350 79688
rect 175918 79608 175924 79620
rect 174418 79580 175924 79608
rect 173526 79500 173532 79552
rect 173584 79540 173590 79552
rect 173866 79540 173894 79580
rect 175918 79568 175924 79580
rect 175976 79568 175982 79620
rect 176102 79568 176108 79620
rect 176160 79608 176166 79620
rect 176672 79608 176700 79840
rect 176160 79580 176700 79608
rect 176810 79608 176838 79840
rect 176902 79744 176930 79908
rect 177160 79880 177166 79892
rect 177132 79840 177166 79880
rect 177218 79840 177224 79892
rect 213086 79840 213092 79892
rect 213144 79880 213150 79892
rect 238754 79880 238760 79892
rect 213144 79852 238760 79880
rect 213144 79840 213150 79852
rect 238754 79840 238760 79852
rect 238812 79840 238818 79892
rect 177132 79756 177160 79840
rect 216766 79772 216772 79824
rect 216824 79812 216830 79824
rect 217410 79812 217416 79824
rect 216824 79784 217416 79812
rect 216824 79772 216830 79784
rect 217410 79772 217416 79784
rect 217468 79812 217474 79824
rect 252554 79812 252560 79824
rect 217468 79784 252560 79812
rect 217468 79772 217474 79784
rect 252554 79772 252560 79784
rect 252612 79772 252618 79824
rect 176902 79716 177068 79744
rect 177040 79620 177068 79716
rect 177114 79704 177120 79756
rect 177172 79704 177178 79756
rect 183738 79704 183744 79756
rect 183796 79744 183802 79756
rect 219986 79744 219992 79756
rect 183796 79716 219992 79744
rect 183796 79704 183802 79716
rect 219986 79704 219992 79716
rect 220044 79704 220050 79756
rect 180426 79636 180432 79688
rect 180484 79676 180490 79688
rect 217502 79676 217508 79688
rect 180484 79648 217508 79676
rect 180484 79636 180490 79648
rect 217502 79636 217508 79648
rect 217560 79636 217566 79688
rect 176930 79608 176936 79620
rect 176810 79580 176936 79608
rect 176160 79568 176166 79580
rect 176930 79568 176936 79580
rect 176988 79568 176994 79620
rect 177022 79568 177028 79620
rect 177080 79568 177086 79620
rect 178954 79568 178960 79620
rect 179012 79608 179018 79620
rect 216030 79608 216036 79620
rect 179012 79580 216036 79608
rect 179012 79568 179018 79580
rect 216030 79568 216036 79580
rect 216088 79608 216094 79620
rect 376754 79608 376760 79620
rect 216088 79580 376760 79608
rect 216088 79568 216094 79580
rect 376754 79568 376760 79580
rect 376812 79568 376818 79620
rect 173584 79512 173894 79540
rect 173584 79500 173590 79512
rect 176654 79500 176660 79552
rect 176712 79540 176718 79552
rect 176838 79540 176844 79552
rect 176712 79512 176844 79540
rect 176712 79500 176718 79512
rect 176838 79500 176844 79512
rect 176896 79500 176902 79552
rect 212166 79500 212172 79552
rect 212224 79540 212230 79552
rect 480254 79540 480260 79552
rect 212224 79512 480260 79540
rect 212224 79500 212230 79512
rect 480254 79500 480260 79512
rect 480312 79500 480318 79552
rect 173986 79432 173992 79484
rect 174044 79472 174050 79484
rect 179414 79472 179420 79484
rect 174044 79444 179420 79472
rect 174044 79432 174050 79444
rect 179414 79432 179420 79444
rect 179472 79432 179478 79484
rect 201402 79432 201408 79484
rect 201460 79472 201466 79484
rect 212902 79472 212908 79484
rect 201460 79444 212908 79472
rect 201460 79432 201466 79444
rect 212902 79432 212908 79444
rect 212960 79472 212966 79484
rect 500954 79472 500960 79484
rect 212960 79444 500960 79472
rect 212960 79432 212966 79444
rect 500954 79432 500960 79444
rect 501012 79432 501018 79484
rect 174906 79364 174912 79416
rect 174964 79404 174970 79416
rect 197262 79404 197268 79416
rect 174964 79376 197268 79404
rect 174964 79364 174970 79376
rect 197262 79364 197268 79376
rect 197320 79364 197326 79416
rect 197354 79364 197360 79416
rect 197412 79404 197418 79416
rect 211982 79404 211988 79416
rect 197412 79376 211988 79404
rect 197412 79364 197418 79376
rect 211982 79364 211988 79376
rect 212040 79404 212046 79416
rect 212166 79404 212172 79416
rect 212040 79376 212172 79404
rect 212040 79364 212046 79376
rect 212166 79364 212172 79376
rect 212224 79364 212230 79416
rect 213730 79364 213736 79416
rect 213788 79404 213794 79416
rect 525794 79404 525800 79416
rect 213788 79376 525800 79404
rect 213788 79364 213794 79376
rect 525794 79364 525800 79376
rect 525852 79364 525858 79416
rect 174446 79296 174452 79348
rect 174504 79336 174510 79348
rect 179506 79336 179512 79348
rect 174504 79308 179512 79336
rect 174504 79296 174510 79308
rect 179506 79296 179512 79308
rect 179564 79296 179570 79348
rect 191282 79296 191288 79348
rect 191340 79336 191346 79348
rect 198182 79336 198188 79348
rect 191340 79308 198188 79336
rect 191340 79296 191346 79308
rect 198182 79296 198188 79308
rect 198240 79296 198246 79348
rect 523126 79336 523132 79348
rect 200086 79308 523132 79336
rect 200086 79280 200114 79308
rect 523126 79296 523132 79308
rect 523184 79296 523190 79348
rect 200022 79268 200028 79280
rect 173452 79240 200028 79268
rect 200022 79228 200028 79240
rect 200080 79240 200114 79280
rect 200080 79228 200086 79240
rect 221182 79228 221188 79280
rect 221240 79268 221246 79280
rect 221366 79268 221372 79280
rect 221240 79240 221372 79268
rect 221240 79228 221246 79240
rect 221366 79228 221372 79240
rect 221424 79228 221430 79280
rect 116394 79160 116400 79212
rect 116452 79200 116458 79212
rect 146846 79200 146852 79212
rect 116452 79172 146852 79200
rect 116452 79160 116458 79172
rect 146846 79160 146852 79172
rect 146904 79160 146910 79212
rect 157306 79172 173020 79200
rect 96154 79132 96160 79144
rect 96080 79104 96160 79132
rect 96154 79092 96160 79104
rect 96212 79092 96218 79144
rect 119798 79092 119804 79144
rect 119856 79132 119862 79144
rect 147214 79132 147220 79144
rect 119856 79104 147220 79132
rect 119856 79092 119862 79104
rect 147214 79092 147220 79104
rect 147272 79092 147278 79144
rect 157306 79132 157334 79172
rect 148520 79104 157334 79132
rect 112530 79024 112536 79076
rect 112588 79064 112594 79076
rect 146110 79064 146116 79076
rect 112588 79036 146116 79064
rect 112588 79024 112594 79036
rect 146110 79024 146116 79036
rect 146168 79064 146174 79076
rect 148520 79064 148548 79104
rect 161934 79092 161940 79144
rect 161992 79092 161998 79144
rect 164878 79092 164884 79144
rect 164936 79132 164942 79144
rect 172514 79132 172520 79144
rect 164936 79104 172520 79132
rect 164936 79092 164942 79104
rect 172514 79092 172520 79104
rect 172572 79092 172578 79144
rect 172992 79132 173020 79172
rect 173066 79160 173072 79212
rect 173124 79200 173130 79212
rect 173986 79200 173992 79212
rect 173124 79172 173992 79200
rect 173124 79160 173130 79172
rect 173986 79160 173992 79172
rect 174044 79160 174050 79212
rect 174078 79160 174084 79212
rect 174136 79200 174142 79212
rect 174538 79200 174544 79212
rect 174136 79172 174544 79200
rect 174136 79160 174142 79172
rect 174538 79160 174544 79172
rect 174596 79200 174602 79212
rect 207658 79200 207664 79212
rect 174596 79172 207664 79200
rect 174596 79160 174602 79172
rect 207658 79160 207664 79172
rect 207716 79160 207722 79212
rect 174446 79132 174452 79144
rect 172992 79104 174452 79132
rect 174446 79092 174452 79104
rect 174504 79092 174510 79144
rect 174630 79092 174636 79144
rect 174688 79132 174694 79144
rect 201310 79132 201316 79144
rect 174688 79104 201316 79132
rect 174688 79092 174694 79104
rect 201310 79092 201316 79104
rect 201368 79092 201374 79144
rect 161952 79064 161980 79092
rect 146168 79036 148548 79064
rect 154546 79036 161980 79064
rect 146168 79024 146174 79036
rect 115106 78956 115112 79008
rect 115164 78996 115170 79008
rect 146294 78996 146300 79008
rect 115164 78968 146300 78996
rect 115164 78956 115170 78968
rect 146294 78956 146300 78968
rect 146352 78996 146358 79008
rect 154546 78996 154574 79036
rect 162854 79024 162860 79076
rect 162912 79064 162918 79076
rect 197906 79064 197912 79076
rect 162912 79036 197912 79064
rect 162912 79024 162918 79036
rect 197906 79024 197912 79036
rect 197964 79024 197970 79076
rect 146352 78968 154574 78996
rect 146352 78956 146358 78968
rect 163406 78956 163412 79008
rect 163464 78996 163470 79008
rect 165246 78996 165252 79008
rect 163464 78968 165252 78996
rect 163464 78956 163470 78968
rect 165246 78956 165252 78968
rect 165304 78956 165310 79008
rect 170490 78956 170496 79008
rect 170548 78996 170554 79008
rect 170766 78996 170772 79008
rect 170548 78968 170772 78996
rect 170548 78956 170554 78968
rect 170766 78956 170772 78968
rect 170824 78956 170830 79008
rect 173342 78956 173348 79008
rect 173400 78996 173406 79008
rect 212810 78996 212816 79008
rect 173400 78968 212816 78996
rect 173400 78956 173406 78968
rect 212810 78956 212816 78968
rect 212868 78996 212874 79008
rect 213730 78996 213736 79008
rect 212868 78968 213736 78996
rect 212868 78956 212874 78968
rect 213730 78956 213736 78968
rect 213788 78956 213794 79008
rect 111242 78888 111248 78940
rect 111300 78928 111306 78940
rect 145834 78928 145840 78940
rect 111300 78900 145840 78928
rect 111300 78888 111306 78900
rect 145834 78888 145840 78900
rect 145892 78928 145898 78940
rect 146018 78928 146024 78940
rect 145892 78900 146024 78928
rect 145892 78888 145898 78900
rect 146018 78888 146024 78900
rect 146076 78888 146082 78940
rect 156046 78888 156052 78940
rect 156104 78928 156110 78940
rect 157058 78928 157064 78940
rect 156104 78900 157064 78928
rect 156104 78888 156110 78900
rect 157058 78888 157064 78900
rect 157116 78888 157122 78940
rect 157518 78888 157524 78940
rect 157576 78928 157582 78940
rect 157886 78928 157892 78940
rect 157576 78900 157892 78928
rect 157576 78888 157582 78900
rect 157886 78888 157892 78900
rect 157944 78888 157950 78940
rect 161198 78888 161204 78940
rect 161256 78928 161262 78940
rect 208946 78928 208952 78940
rect 161256 78900 208952 78928
rect 161256 78888 161262 78900
rect 208946 78888 208952 78900
rect 209004 78888 209010 78940
rect 124122 78820 124128 78872
rect 124180 78860 124186 78872
rect 140590 78860 140596 78872
rect 124180 78832 128354 78860
rect 124180 78820 124186 78832
rect 128326 78792 128354 78832
rect 133846 78832 140596 78860
rect 133846 78792 133874 78832
rect 140590 78820 140596 78832
rect 140648 78820 140654 78872
rect 150710 78820 150716 78872
rect 150768 78860 150774 78872
rect 213086 78860 213092 78872
rect 150768 78832 213092 78860
rect 150768 78820 150774 78832
rect 213086 78820 213092 78832
rect 213144 78820 213150 78872
rect 128326 78764 133874 78792
rect 134242 78752 134248 78804
rect 134300 78792 134306 78804
rect 147858 78792 147864 78804
rect 134300 78764 147864 78792
rect 134300 78752 134306 78764
rect 147858 78752 147864 78764
rect 147916 78752 147922 78804
rect 152090 78752 152096 78804
rect 152148 78792 152154 78804
rect 216766 78792 216772 78804
rect 152148 78764 216772 78792
rect 152148 78752 152154 78764
rect 216766 78752 216772 78764
rect 216824 78752 216830 78804
rect 130838 78684 130844 78736
rect 130896 78724 130902 78736
rect 137002 78724 137008 78736
rect 130896 78696 137008 78724
rect 130896 78684 130902 78696
rect 137002 78684 137008 78696
rect 137060 78684 137066 78736
rect 142430 78724 142436 78736
rect 137112 78696 142436 78724
rect 99926 78616 99932 78668
rect 99984 78656 99990 78668
rect 99984 78628 122834 78656
rect 99984 78616 99990 78628
rect 122806 78588 122834 78628
rect 125502 78616 125508 78668
rect 125560 78656 125566 78668
rect 134058 78656 134064 78668
rect 125560 78628 134064 78656
rect 125560 78616 125566 78628
rect 134058 78616 134064 78628
rect 134116 78616 134122 78668
rect 130286 78588 130292 78600
rect 122806 78560 130292 78588
rect 130286 78548 130292 78560
rect 130344 78548 130350 78600
rect 132310 78548 132316 78600
rect 132368 78588 132374 78600
rect 137112 78588 137140 78696
rect 142430 78684 142436 78696
rect 142488 78684 142494 78736
rect 155954 78684 155960 78736
rect 156012 78724 156018 78736
rect 157242 78724 157248 78736
rect 156012 78696 157248 78724
rect 156012 78684 156018 78696
rect 157242 78684 157248 78696
rect 157300 78684 157306 78736
rect 159082 78684 159088 78736
rect 159140 78724 159146 78736
rect 160094 78724 160100 78736
rect 159140 78696 160100 78724
rect 159140 78684 159146 78696
rect 160094 78684 160100 78696
rect 160152 78684 160158 78736
rect 162578 78684 162584 78736
rect 162636 78724 162642 78736
rect 162636 78696 166856 78724
rect 162636 78684 162642 78696
rect 138474 78616 138480 78668
rect 138532 78656 138538 78668
rect 138750 78656 138756 78668
rect 138532 78628 138756 78656
rect 138532 78616 138538 78628
rect 138750 78616 138756 78628
rect 138808 78616 138814 78668
rect 140222 78616 140228 78668
rect 140280 78656 140286 78668
rect 140682 78656 140688 78668
rect 140280 78628 140688 78656
rect 140280 78616 140286 78628
rect 140682 78616 140688 78628
rect 140740 78616 140746 78668
rect 141234 78616 141240 78668
rect 141292 78656 141298 78668
rect 141602 78656 141608 78668
rect 141292 78628 141608 78656
rect 141292 78616 141298 78628
rect 141602 78616 141608 78628
rect 141660 78616 141666 78668
rect 147030 78616 147036 78668
rect 147088 78656 147094 78668
rect 147398 78656 147404 78668
rect 147088 78628 147404 78656
rect 147088 78616 147094 78628
rect 147398 78616 147404 78628
rect 147456 78616 147462 78668
rect 156046 78616 156052 78668
rect 156104 78656 156110 78668
rect 156874 78656 156880 78668
rect 156104 78628 156880 78656
rect 156104 78616 156110 78628
rect 156874 78616 156880 78628
rect 156932 78616 156938 78668
rect 165982 78616 165988 78668
rect 166040 78656 166046 78668
rect 166718 78656 166724 78668
rect 166040 78628 166724 78656
rect 166040 78616 166046 78628
rect 166718 78616 166724 78628
rect 166776 78616 166782 78668
rect 166828 78656 166856 78696
rect 168006 78684 168012 78736
rect 168064 78724 168070 78736
rect 179322 78724 179328 78736
rect 168064 78696 179328 78724
rect 168064 78684 168070 78696
rect 179322 78684 179328 78696
rect 179380 78684 179386 78736
rect 201310 78684 201316 78736
rect 201368 78724 201374 78736
rect 539686 78724 539692 78736
rect 201368 78696 539692 78724
rect 201368 78684 201374 78696
rect 539686 78684 539692 78696
rect 539744 78684 539750 78736
rect 171870 78656 171876 78668
rect 166828 78628 171876 78656
rect 171870 78616 171876 78628
rect 171928 78616 171934 78668
rect 172698 78616 172704 78668
rect 172756 78656 172762 78668
rect 172882 78656 172888 78668
rect 172756 78628 172888 78656
rect 172756 78616 172762 78628
rect 172882 78616 172888 78628
rect 172940 78616 172946 78668
rect 172974 78616 172980 78668
rect 173032 78656 173038 78668
rect 174906 78656 174912 78668
rect 173032 78628 174912 78656
rect 173032 78616 173038 78628
rect 174906 78616 174912 78628
rect 174964 78616 174970 78668
rect 176654 78616 176660 78668
rect 176712 78656 176718 78668
rect 177206 78656 177212 78668
rect 176712 78628 177212 78656
rect 176712 78616 176718 78628
rect 177206 78616 177212 78628
rect 177264 78616 177270 78668
rect 132368 78560 137140 78588
rect 132368 78548 132374 78560
rect 156230 78548 156236 78600
rect 156288 78588 156294 78600
rect 156288 78560 164234 78588
rect 156288 78548 156294 78560
rect 119430 78480 119436 78532
rect 119488 78520 119494 78532
rect 145374 78520 145380 78532
rect 119488 78492 145380 78520
rect 119488 78480 119494 78492
rect 145374 78480 145380 78492
rect 145432 78480 145438 78532
rect 158898 78480 158904 78532
rect 158956 78520 158962 78532
rect 159726 78520 159732 78532
rect 158956 78492 159732 78520
rect 158956 78480 158962 78492
rect 159726 78480 159732 78492
rect 159784 78480 159790 78532
rect 164206 78520 164234 78560
rect 165430 78548 165436 78600
rect 165488 78588 165494 78600
rect 215846 78588 215852 78600
rect 165488 78560 215852 78588
rect 165488 78548 165494 78560
rect 215846 78548 215852 78560
rect 215904 78548 215910 78600
rect 191558 78520 191564 78532
rect 164206 78492 191564 78520
rect 191558 78480 191564 78492
rect 191616 78520 191622 78532
rect 191742 78520 191748 78532
rect 191616 78492 191748 78520
rect 191616 78480 191622 78492
rect 191742 78480 191748 78492
rect 191800 78480 191806 78532
rect 133138 78452 133144 78464
rect 122806 78424 133144 78452
rect 119522 78344 119528 78396
rect 119580 78384 119586 78396
rect 122806 78384 122834 78424
rect 133138 78412 133144 78424
rect 133196 78412 133202 78464
rect 163038 78412 163044 78464
rect 163096 78452 163102 78464
rect 167454 78452 167460 78464
rect 163096 78424 167460 78452
rect 163096 78412 163102 78424
rect 167454 78412 167460 78424
rect 167512 78412 167518 78464
rect 168098 78412 168104 78464
rect 168156 78452 168162 78464
rect 197906 78452 197912 78464
rect 168156 78424 197912 78452
rect 168156 78412 168162 78424
rect 197906 78412 197912 78424
rect 197964 78412 197970 78464
rect 119580 78356 122834 78384
rect 119580 78344 119586 78356
rect 129458 78344 129464 78396
rect 129516 78384 129522 78396
rect 142338 78384 142344 78396
rect 129516 78356 142344 78384
rect 129516 78344 129522 78356
rect 142338 78344 142344 78356
rect 142396 78344 142402 78396
rect 161014 78344 161020 78396
rect 161072 78384 161078 78396
rect 168006 78384 168012 78396
rect 161072 78356 168012 78384
rect 161072 78344 161078 78356
rect 168006 78344 168012 78356
rect 168064 78344 168070 78396
rect 168650 78344 168656 78396
rect 168708 78384 168714 78396
rect 168834 78384 168840 78396
rect 168708 78356 168840 78384
rect 168708 78344 168714 78356
rect 168834 78344 168840 78356
rect 168892 78344 168898 78396
rect 169662 78344 169668 78396
rect 169720 78384 169726 78396
rect 199010 78384 199016 78396
rect 169720 78356 199016 78384
rect 169720 78344 169726 78356
rect 199010 78344 199016 78356
rect 199068 78344 199074 78396
rect 108298 78276 108304 78328
rect 108356 78316 108362 78328
rect 131942 78316 131948 78328
rect 108356 78288 131948 78316
rect 108356 78276 108362 78288
rect 131942 78276 131948 78288
rect 132000 78276 132006 78328
rect 132218 78276 132224 78328
rect 132276 78316 132282 78328
rect 137554 78316 137560 78328
rect 132276 78288 137560 78316
rect 132276 78276 132282 78288
rect 137554 78276 137560 78288
rect 137612 78276 137618 78328
rect 168742 78276 168748 78328
rect 168800 78316 168806 78328
rect 169294 78316 169300 78328
rect 168800 78288 169300 78316
rect 168800 78276 168806 78288
rect 169294 78276 169300 78288
rect 169352 78276 169358 78328
rect 173894 78276 173900 78328
rect 173952 78316 173958 78328
rect 174630 78316 174636 78328
rect 173952 78288 174636 78316
rect 173952 78276 173958 78288
rect 174630 78276 174636 78288
rect 174688 78276 174694 78328
rect 175366 78276 175372 78328
rect 175424 78316 175430 78328
rect 178218 78316 178224 78328
rect 175424 78288 178224 78316
rect 175424 78276 175430 78288
rect 178218 78276 178224 78288
rect 178276 78276 178282 78328
rect 179322 78276 179328 78328
rect 179380 78316 179386 78328
rect 202322 78316 202328 78328
rect 179380 78288 202328 78316
rect 179380 78276 179386 78288
rect 202322 78276 202328 78288
rect 202380 78276 202386 78328
rect 104526 78208 104532 78260
rect 104584 78248 104590 78260
rect 127158 78248 127164 78260
rect 104584 78220 127164 78248
rect 104584 78208 104590 78220
rect 127158 78208 127164 78220
rect 127216 78208 127222 78260
rect 129642 78208 129648 78260
rect 129700 78248 129706 78260
rect 142246 78248 142252 78260
rect 129700 78220 142252 78248
rect 129700 78208 129706 78220
rect 142246 78208 142252 78220
rect 142304 78208 142310 78260
rect 158806 78208 158812 78260
rect 158864 78248 158870 78260
rect 159818 78248 159824 78260
rect 158864 78220 159824 78248
rect 158864 78208 158870 78220
rect 159818 78208 159824 78220
rect 159876 78208 159882 78260
rect 167914 78208 167920 78260
rect 167972 78248 167978 78260
rect 169662 78248 169668 78260
rect 167972 78220 169668 78248
rect 167972 78208 167978 78220
rect 169662 78208 169668 78220
rect 169720 78208 169726 78260
rect 172514 78208 172520 78260
rect 172572 78248 172578 78260
rect 183738 78248 183744 78260
rect 172572 78220 183744 78248
rect 172572 78208 172578 78220
rect 183738 78208 183744 78220
rect 183796 78248 183802 78260
rect 184198 78248 184204 78260
rect 183796 78220 184204 78248
rect 183796 78208 183802 78220
rect 184198 78208 184204 78220
rect 184256 78208 184262 78260
rect 107010 78140 107016 78192
rect 107068 78180 107074 78192
rect 129826 78180 129832 78192
rect 107068 78152 129832 78180
rect 107068 78140 107074 78152
rect 129826 78140 129832 78152
rect 129884 78180 129890 78192
rect 130746 78180 130752 78192
rect 129884 78152 130752 78180
rect 129884 78140 129890 78152
rect 130746 78140 130752 78152
rect 130804 78140 130810 78192
rect 138198 78140 138204 78192
rect 138256 78180 138262 78192
rect 139026 78180 139032 78192
rect 138256 78152 139032 78180
rect 138256 78140 138262 78152
rect 139026 78140 139032 78152
rect 139084 78140 139090 78192
rect 154942 78140 154948 78192
rect 155000 78180 155006 78192
rect 165430 78180 165436 78192
rect 155000 78152 165436 78180
rect 155000 78140 155006 78152
rect 165430 78140 165436 78152
rect 165488 78140 165494 78192
rect 166442 78140 166448 78192
rect 166500 78180 166506 78192
rect 180150 78180 180156 78192
rect 166500 78152 180156 78180
rect 166500 78140 166506 78152
rect 180150 78140 180156 78152
rect 180208 78180 180214 78192
rect 180426 78180 180432 78192
rect 180208 78152 180432 78180
rect 180208 78140 180214 78152
rect 180426 78140 180432 78152
rect 180484 78140 180490 78192
rect 180610 78140 180616 78192
rect 180668 78180 180674 78192
rect 200482 78180 200488 78192
rect 180668 78152 200488 78180
rect 180668 78140 180674 78152
rect 200482 78140 200488 78152
rect 200540 78140 200546 78192
rect 104066 78072 104072 78124
rect 104124 78112 104130 78124
rect 127710 78112 127716 78124
rect 104124 78084 127716 78112
rect 104124 78072 104130 78084
rect 127710 78072 127716 78084
rect 127768 78072 127774 78124
rect 141786 78112 141792 78124
rect 133846 78084 141792 78112
rect 101306 78004 101312 78056
rect 101364 78044 101370 78056
rect 128262 78044 128268 78056
rect 101364 78016 128268 78044
rect 101364 78004 101370 78016
rect 128262 78004 128268 78016
rect 128320 78004 128326 78056
rect 131022 78004 131028 78056
rect 131080 78044 131086 78056
rect 133846 78044 133874 78084
rect 141786 78072 141792 78084
rect 141844 78072 141850 78124
rect 157426 78072 157432 78124
rect 157484 78112 157490 78124
rect 163038 78112 163044 78124
rect 157484 78084 163044 78112
rect 157484 78072 157490 78084
rect 163038 78072 163044 78084
rect 163096 78072 163102 78124
rect 163590 78072 163596 78124
rect 163648 78112 163654 78124
rect 179230 78112 179236 78124
rect 163648 78084 179236 78112
rect 163648 78072 163654 78084
rect 179230 78072 179236 78084
rect 179288 78112 179294 78124
rect 179288 78084 180656 78112
rect 179288 78072 179294 78084
rect 131080 78016 133874 78044
rect 131080 78004 131086 78016
rect 168650 78004 168656 78056
rect 168708 78044 168714 78056
rect 169386 78044 169392 78056
rect 168708 78016 169392 78044
rect 168708 78004 168714 78016
rect 169386 78004 169392 78016
rect 169444 78004 169450 78056
rect 178862 78044 178868 78056
rect 172486 78016 178868 78044
rect 46934 77936 46940 77988
rect 46992 77976 46998 77988
rect 105630 77976 105636 77988
rect 46992 77948 105636 77976
rect 46992 77936 46998 77948
rect 105630 77936 105636 77948
rect 105688 77936 105694 77988
rect 106734 77936 106740 77988
rect 106792 77976 106798 77988
rect 131298 77976 131304 77988
rect 106792 77948 131304 77976
rect 106792 77936 106798 77948
rect 131298 77936 131304 77948
rect 131356 77976 131362 77988
rect 131666 77976 131672 77988
rect 131356 77948 131672 77976
rect 131356 77936 131362 77948
rect 131666 77936 131672 77948
rect 131724 77936 131730 77988
rect 132310 77936 132316 77988
rect 132368 77976 132374 77988
rect 141418 77976 141424 77988
rect 132368 77948 141424 77976
rect 132368 77936 132374 77948
rect 141418 77936 141424 77948
rect 141476 77936 141482 77988
rect 164326 77936 164332 77988
rect 164384 77976 164390 77988
rect 172486 77976 172514 78016
rect 178862 78004 178868 78016
rect 178920 78004 178926 78056
rect 180628 78044 180656 78084
rect 180702 78072 180708 78124
rect 180760 78112 180766 78124
rect 202046 78112 202052 78124
rect 180760 78084 202052 78112
rect 180760 78072 180766 78084
rect 202046 78072 202052 78084
rect 202104 78072 202110 78124
rect 214742 78044 214748 78056
rect 180628 78016 214748 78044
rect 214742 78004 214748 78016
rect 214800 78004 214806 78056
rect 215846 78004 215852 78056
rect 215904 78044 215910 78056
rect 216122 78044 216128 78056
rect 215904 78016 216128 78044
rect 215904 78004 215910 78016
rect 216122 78004 216128 78016
rect 216180 78044 216186 78056
rect 270494 78044 270500 78056
rect 216180 78016 270500 78044
rect 216180 78004 216186 78016
rect 270494 78004 270500 78016
rect 270552 78004 270558 78056
rect 164384 77948 172514 77976
rect 164384 77936 164390 77948
rect 173894 77936 173900 77988
rect 173952 77976 173958 77988
rect 174262 77976 174268 77988
rect 173952 77948 174268 77976
rect 173952 77936 173958 77948
rect 174262 77936 174268 77948
rect 174320 77936 174326 77988
rect 181622 77976 181628 77988
rect 176626 77948 181628 77976
rect 103146 77868 103152 77920
rect 103204 77908 103210 77920
rect 124214 77908 124220 77920
rect 103204 77880 124220 77908
rect 103204 77868 103210 77880
rect 124214 77868 124220 77880
rect 124272 77908 124278 77920
rect 125502 77908 125508 77920
rect 124272 77880 125508 77908
rect 124272 77868 124278 77880
rect 125502 77868 125508 77880
rect 125560 77868 125566 77920
rect 133966 77868 133972 77920
rect 134024 77908 134030 77920
rect 134610 77908 134616 77920
rect 134024 77880 134616 77908
rect 134024 77868 134030 77880
rect 134610 77868 134616 77880
rect 134668 77868 134674 77920
rect 141878 77908 141884 77920
rect 136928 77880 141884 77908
rect 109586 77800 109592 77852
rect 109644 77840 109650 77852
rect 127618 77840 127624 77852
rect 109644 77812 127624 77840
rect 109644 77800 109650 77812
rect 127618 77800 127624 77812
rect 127676 77800 127682 77852
rect 130838 77800 130844 77852
rect 130896 77840 130902 77852
rect 136928 77840 136956 77880
rect 141878 77868 141884 77880
rect 141936 77868 141942 77920
rect 166902 77868 166908 77920
rect 166960 77908 166966 77920
rect 176626 77908 176654 77948
rect 181622 77936 181628 77948
rect 181680 77976 181686 77988
rect 182082 77976 182088 77988
rect 181680 77948 182088 77976
rect 181680 77936 181686 77948
rect 182082 77936 182088 77948
rect 182140 77936 182146 77988
rect 191742 77936 191748 77988
rect 191800 77976 191806 77988
rect 306374 77976 306380 77988
rect 191800 77948 306380 77976
rect 191800 77936 191806 77948
rect 306374 77936 306380 77948
rect 306432 77936 306438 77988
rect 166960 77880 176654 77908
rect 166960 77868 166966 77880
rect 179322 77868 179328 77920
rect 179380 77908 179386 77920
rect 197998 77908 198004 77920
rect 179380 77880 198004 77908
rect 179380 77868 179386 77880
rect 197998 77868 198004 77880
rect 198056 77868 198062 77920
rect 130896 77812 136956 77840
rect 130896 77800 130902 77812
rect 137002 77800 137008 77852
rect 137060 77840 137066 77852
rect 144914 77840 144920 77852
rect 137060 77812 144920 77840
rect 137060 77800 137066 77812
rect 144914 77800 144920 77812
rect 144972 77800 144978 77852
rect 160462 77800 160468 77852
rect 160520 77840 160526 77852
rect 162118 77840 162124 77852
rect 160520 77812 162124 77840
rect 160520 77800 160526 77812
rect 162118 77800 162124 77812
rect 162176 77800 162182 77852
rect 172514 77800 172520 77852
rect 172572 77840 172578 77852
rect 172790 77840 172796 77852
rect 172572 77812 172796 77840
rect 172572 77800 172578 77812
rect 172790 77800 172796 77812
rect 172848 77800 172854 77852
rect 175918 77800 175924 77852
rect 175976 77840 175982 77852
rect 177206 77840 177212 77852
rect 175976 77812 177212 77840
rect 175976 77800 175982 77812
rect 177206 77800 177212 77812
rect 177264 77800 177270 77852
rect 180426 77800 180432 77852
rect 180484 77840 180490 77852
rect 195238 77840 195244 77852
rect 180484 77812 195244 77840
rect 180484 77800 180490 77812
rect 195238 77800 195244 77812
rect 195296 77800 195302 77852
rect 129550 77732 129556 77784
rect 129608 77772 129614 77784
rect 142154 77772 142160 77784
rect 129608 77744 142160 77772
rect 129608 77732 129614 77744
rect 142154 77732 142160 77744
rect 142212 77732 142218 77784
rect 166350 77732 166356 77784
rect 166408 77772 166414 77784
rect 180334 77772 180340 77784
rect 166408 77744 180340 77772
rect 166408 77732 166414 77744
rect 180334 77732 180340 77744
rect 180392 77732 180398 77784
rect 123754 77664 123760 77716
rect 123812 77704 123818 77716
rect 141694 77704 141700 77716
rect 123812 77676 141700 77704
rect 123812 77664 123818 77676
rect 141694 77664 141700 77676
rect 141752 77664 141758 77716
rect 162486 77664 162492 77716
rect 162544 77704 162550 77716
rect 178954 77704 178960 77716
rect 162544 77676 178960 77704
rect 162544 77664 162550 77676
rect 178954 77664 178960 77676
rect 179012 77664 179018 77716
rect 180058 77664 180064 77716
rect 180116 77704 180122 77716
rect 194042 77704 194048 77716
rect 180116 77676 194048 77704
rect 180116 77664 180122 77676
rect 194042 77664 194048 77676
rect 194100 77664 194106 77716
rect 105722 77596 105728 77648
rect 105780 77636 105786 77648
rect 137186 77636 137192 77648
rect 105780 77608 137192 77636
rect 105780 77596 105786 77608
rect 137186 77596 137192 77608
rect 137244 77596 137250 77648
rect 153470 77596 153476 77648
rect 153528 77636 153534 77648
rect 215846 77636 215852 77648
rect 153528 77608 215852 77636
rect 153528 77596 153534 77608
rect 215846 77596 215852 77608
rect 215904 77596 215910 77648
rect 105630 77528 105636 77580
rect 105688 77568 105694 77580
rect 135070 77568 135076 77580
rect 105688 77540 135076 77568
rect 105688 77528 105694 77540
rect 135070 77528 135076 77540
rect 135128 77528 135134 77580
rect 142246 77528 142252 77580
rect 142304 77568 142310 77580
rect 142982 77568 142988 77580
rect 142304 77540 142988 77568
rect 142304 77528 142310 77540
rect 142982 77528 142988 77540
rect 143040 77528 143046 77580
rect 152458 77528 152464 77580
rect 152516 77568 152522 77580
rect 152734 77568 152740 77580
rect 152516 77540 152740 77568
rect 152516 77528 152522 77540
rect 152734 77528 152740 77540
rect 152792 77528 152798 77580
rect 157150 77528 157156 77580
rect 157208 77568 157214 77580
rect 162578 77568 162584 77580
rect 157208 77540 162584 77568
rect 157208 77528 157214 77540
rect 162578 77528 162584 77540
rect 162636 77528 162642 77580
rect 165798 77528 165804 77580
rect 165856 77568 165862 77580
rect 165856 77540 167408 77568
rect 165856 77528 165862 77540
rect 126974 77460 126980 77512
rect 127032 77500 127038 77512
rect 129642 77500 129648 77512
rect 127032 77472 129648 77500
rect 127032 77460 127038 77472
rect 129642 77460 129648 77472
rect 129700 77460 129706 77512
rect 130930 77460 130936 77512
rect 130988 77500 130994 77512
rect 140038 77500 140044 77512
rect 130988 77472 140044 77500
rect 130988 77460 130994 77472
rect 140038 77460 140044 77472
rect 140096 77460 140102 77512
rect 142706 77460 142712 77512
rect 142764 77500 142770 77512
rect 142890 77500 142896 77512
rect 142764 77472 142896 77500
rect 142764 77460 142770 77472
rect 142890 77460 142896 77472
rect 142948 77460 142954 77512
rect 161842 77460 161848 77512
rect 161900 77500 161906 77512
rect 166902 77500 166908 77512
rect 161900 77472 166908 77500
rect 161900 77460 161906 77472
rect 166902 77460 166908 77472
rect 166960 77460 166966 77512
rect 167380 77500 167408 77540
rect 167454 77528 167460 77580
rect 167512 77568 167518 77580
rect 179322 77568 179328 77580
rect 167512 77540 179328 77568
rect 167512 77528 167518 77540
rect 179322 77528 179328 77540
rect 179380 77528 179386 77580
rect 180610 77500 180616 77512
rect 167380 77472 180616 77500
rect 180610 77460 180616 77472
rect 180668 77460 180674 77512
rect 133138 77392 133144 77444
rect 133196 77432 133202 77444
rect 143534 77432 143540 77444
rect 133196 77404 143540 77432
rect 133196 77392 133202 77404
rect 143534 77392 143540 77404
rect 143592 77392 143598 77444
rect 143994 77392 144000 77444
rect 144052 77432 144058 77444
rect 144052 77404 144132 77432
rect 144052 77392 144058 77404
rect 144104 77376 144132 77404
rect 144086 77324 144092 77376
rect 144144 77324 144150 77376
rect 161474 77324 161480 77376
rect 161532 77364 161538 77376
rect 161842 77364 161848 77376
rect 161532 77336 161848 77364
rect 161532 77324 161538 77336
rect 161842 77324 161848 77336
rect 161900 77324 161906 77376
rect 197906 77324 197912 77376
rect 197964 77364 197970 77376
rect 287698 77364 287704 77376
rect 197964 77336 287704 77364
rect 197964 77324 197970 77336
rect 287698 77324 287704 77336
rect 287756 77324 287762 77376
rect 135714 77256 135720 77308
rect 135772 77296 135778 77308
rect 136082 77296 136088 77308
rect 135772 77268 136088 77296
rect 135772 77256 135778 77268
rect 136082 77256 136088 77268
rect 136140 77256 136146 77308
rect 137002 77256 137008 77308
rect 137060 77296 137066 77308
rect 137278 77296 137284 77308
rect 137060 77268 137284 77296
rect 137060 77256 137066 77268
rect 137278 77256 137284 77268
rect 137336 77256 137342 77308
rect 142614 77256 142620 77308
rect 142672 77296 142678 77308
rect 143350 77296 143356 77308
rect 142672 77268 143356 77296
rect 142672 77256 142678 77268
rect 143350 77256 143356 77268
rect 143408 77256 143414 77308
rect 153470 77256 153476 77308
rect 153528 77296 153534 77308
rect 153838 77296 153844 77308
rect 153528 77268 153844 77296
rect 153528 77256 153534 77268
rect 153838 77256 153844 77268
rect 153896 77256 153902 77308
rect 164234 77256 164240 77308
rect 164292 77296 164298 77308
rect 165522 77296 165528 77308
rect 164292 77268 165528 77296
rect 164292 77256 164298 77268
rect 165522 77256 165528 77268
rect 165580 77256 165586 77308
rect 199010 77256 199016 77308
rect 199068 77296 199074 77308
rect 453298 77296 453304 77308
rect 199068 77268 453304 77296
rect 199068 77256 199074 77268
rect 453298 77256 453304 77268
rect 453356 77256 453362 77308
rect 101214 77188 101220 77240
rect 101272 77228 101278 77240
rect 101272 77200 147674 77228
rect 101272 77188 101278 77200
rect 99006 77120 99012 77172
rect 99064 77160 99070 77172
rect 146386 77160 146392 77172
rect 99064 77132 146392 77160
rect 99064 77120 99070 77132
rect 146386 77120 146392 77132
rect 146444 77120 146450 77172
rect 96154 77052 96160 77104
rect 96212 77092 96218 77104
rect 138566 77092 138572 77104
rect 96212 77064 138572 77092
rect 96212 77052 96218 77064
rect 138566 77052 138572 77064
rect 138624 77052 138630 77104
rect 114278 76984 114284 77036
rect 114336 77024 114342 77036
rect 146570 77024 146576 77036
rect 114336 76996 146576 77024
rect 114336 76984 114342 76996
rect 146570 76984 146576 76996
rect 146628 76984 146634 77036
rect 111610 76916 111616 76968
rect 111668 76956 111674 76968
rect 143350 76956 143356 76968
rect 111668 76928 143356 76956
rect 111668 76916 111674 76928
rect 143350 76916 143356 76928
rect 143408 76916 143414 76968
rect 105354 76848 105360 76900
rect 105412 76888 105418 76900
rect 132218 76888 132224 76900
rect 105412 76860 132224 76888
rect 105412 76848 105418 76860
rect 132218 76848 132224 76860
rect 132276 76848 132282 76900
rect 134518 76848 134524 76900
rect 134576 76888 134582 76900
rect 134794 76888 134800 76900
rect 134576 76860 134800 76888
rect 134576 76848 134582 76860
rect 134794 76848 134800 76860
rect 134852 76848 134858 76900
rect 144178 76848 144184 76900
rect 144236 76888 144242 76900
rect 144362 76888 144368 76900
rect 144236 76860 144368 76888
rect 144236 76848 144242 76860
rect 144362 76848 144368 76860
rect 144420 76848 144426 76900
rect 115658 76780 115664 76832
rect 115716 76820 115722 76832
rect 147030 76820 147036 76832
rect 115716 76792 147036 76820
rect 115716 76780 115722 76792
rect 147030 76780 147036 76792
rect 147088 76780 147094 76832
rect 114002 76712 114008 76764
rect 114060 76752 114066 76764
rect 143442 76752 143448 76764
rect 114060 76724 143448 76752
rect 114060 76712 114066 76724
rect 143442 76712 143448 76724
rect 143500 76712 143506 76764
rect 116946 76644 116952 76696
rect 117004 76684 117010 76696
rect 147306 76684 147312 76696
rect 117004 76656 147312 76684
rect 117004 76644 117010 76656
rect 147306 76644 147312 76656
rect 147364 76644 147370 76696
rect 96430 76576 96436 76628
rect 96488 76616 96494 76628
rect 125594 76616 125600 76628
rect 96488 76588 125600 76616
rect 96488 76576 96494 76588
rect 125594 76576 125600 76588
rect 125652 76576 125658 76628
rect 128262 76576 128268 76628
rect 128320 76616 128326 76628
rect 131390 76616 131396 76628
rect 128320 76588 131396 76616
rect 128320 76576 128326 76588
rect 131390 76576 131396 76588
rect 131448 76616 131454 76628
rect 135346 76616 135352 76628
rect 131448 76588 135352 76616
rect 131448 76576 131454 76588
rect 135346 76576 135352 76588
rect 135404 76576 135410 76628
rect 136634 76576 136640 76628
rect 136692 76616 136698 76628
rect 137462 76616 137468 76628
rect 136692 76588 137468 76616
rect 136692 76576 136698 76588
rect 137462 76576 137468 76588
rect 137520 76576 137526 76628
rect 144914 76576 144920 76628
rect 144972 76616 144978 76628
rect 146018 76616 146024 76628
rect 144972 76588 146024 76616
rect 144972 76576 144978 76588
rect 146018 76576 146024 76588
rect 146076 76576 146082 76628
rect 147646 76616 147674 77200
rect 155402 77188 155408 77240
rect 155460 77228 155466 77240
rect 218054 77228 218060 77240
rect 155460 77200 218060 77228
rect 155460 77188 155466 77200
rect 218054 77188 218060 77200
rect 218112 77188 218118 77240
rect 218330 77188 218336 77240
rect 218388 77228 218394 77240
rect 218388 77200 218560 77228
rect 218388 77188 218394 77200
rect 218422 77160 218428 77172
rect 162136 77132 218428 77160
rect 155126 76984 155132 77036
rect 155184 77024 155190 77036
rect 162136 77024 162164 77132
rect 218422 77120 218428 77132
rect 218480 77120 218486 77172
rect 218532 77092 218560 77200
rect 218882 77092 218888 77104
rect 155184 76996 162164 77024
rect 162228 77064 218888 77092
rect 155184 76984 155190 76996
rect 157334 76916 157340 76968
rect 157392 76956 157398 76968
rect 157702 76956 157708 76968
rect 157392 76928 157708 76956
rect 157392 76916 157398 76928
rect 157702 76916 157708 76928
rect 157760 76916 157766 76968
rect 159910 76916 159916 76968
rect 159968 76956 159974 76968
rect 162228 76956 162256 77064
rect 218882 77052 218888 77064
rect 218940 77052 218946 77104
rect 164326 76984 164332 77036
rect 164384 77024 164390 77036
rect 164786 77024 164792 77036
rect 164384 76996 164792 77024
rect 164384 76984 164390 76996
rect 164786 76984 164792 76996
rect 164844 76984 164850 77036
rect 208854 77024 208860 77036
rect 166966 76996 208860 77024
rect 159968 76928 162256 76956
rect 159968 76916 159974 76928
rect 164602 76916 164608 76968
rect 164660 76956 164666 76968
rect 165522 76956 165528 76968
rect 164660 76928 165528 76956
rect 164660 76916 164666 76928
rect 165522 76916 165528 76928
rect 165580 76916 165586 76968
rect 153194 76848 153200 76900
rect 153252 76888 153258 76900
rect 154298 76888 154304 76900
rect 153252 76860 154304 76888
rect 153252 76848 153258 76860
rect 154298 76848 154304 76860
rect 154356 76848 154362 76900
rect 154758 76848 154764 76900
rect 154816 76888 154822 76900
rect 154942 76888 154948 76900
rect 154816 76860 154948 76888
rect 154816 76848 154822 76860
rect 154942 76848 154948 76860
rect 155000 76848 155006 76900
rect 160738 76848 160744 76900
rect 160796 76888 160802 76900
rect 166966 76888 166994 76996
rect 208854 76984 208860 76996
rect 208912 76984 208918 77036
rect 167454 76916 167460 76968
rect 167512 76956 167518 76968
rect 168190 76956 168196 76968
rect 167512 76928 168196 76956
rect 167512 76916 167518 76928
rect 168190 76916 168196 76928
rect 168248 76916 168254 76968
rect 171778 76916 171784 76968
rect 171836 76956 171842 76968
rect 196158 76956 196164 76968
rect 171836 76928 196164 76956
rect 171836 76916 171842 76928
rect 196158 76916 196164 76928
rect 196216 76916 196222 76968
rect 160796 76860 166994 76888
rect 160796 76848 160802 76860
rect 168834 76848 168840 76900
rect 168892 76888 168898 76900
rect 169202 76888 169208 76900
rect 168892 76860 169208 76888
rect 168892 76848 168898 76860
rect 169202 76848 169208 76860
rect 169260 76848 169266 76900
rect 173526 76848 173532 76900
rect 173584 76888 173590 76900
rect 174262 76888 174268 76900
rect 173584 76860 174268 76888
rect 173584 76848 173590 76860
rect 174262 76848 174268 76860
rect 174320 76848 174326 76900
rect 175366 76848 175372 76900
rect 175424 76888 175430 76900
rect 176562 76888 176568 76900
rect 175424 76860 176568 76888
rect 175424 76848 175430 76860
rect 176562 76848 176568 76860
rect 176620 76848 176626 76900
rect 177942 76848 177948 76900
rect 178000 76888 178006 76900
rect 211798 76888 211804 76900
rect 178000 76860 211804 76888
rect 178000 76848 178006 76860
rect 211798 76848 211804 76860
rect 211856 76848 211862 76900
rect 157334 76780 157340 76832
rect 157392 76820 157398 76832
rect 157978 76820 157984 76832
rect 157392 76792 157984 76820
rect 157392 76780 157398 76792
rect 157978 76780 157984 76792
rect 158036 76780 158042 76832
rect 168190 76780 168196 76832
rect 168248 76820 168254 76832
rect 169662 76820 169668 76832
rect 168248 76792 169668 76820
rect 168248 76780 168254 76792
rect 169662 76780 169668 76792
rect 169720 76820 169726 76832
rect 201954 76820 201960 76832
rect 169720 76792 201960 76820
rect 169720 76780 169726 76792
rect 201954 76780 201960 76792
rect 202012 76780 202018 76832
rect 154758 76712 154764 76764
rect 154816 76752 154822 76764
rect 155034 76752 155040 76764
rect 154816 76724 155040 76752
rect 154816 76712 154822 76724
rect 155034 76712 155040 76724
rect 155092 76712 155098 76764
rect 170214 76712 170220 76764
rect 170272 76752 170278 76764
rect 171962 76752 171968 76764
rect 170272 76724 171968 76752
rect 170272 76712 170278 76724
rect 171962 76712 171968 76724
rect 172020 76712 172026 76764
rect 172606 76712 172612 76764
rect 172664 76752 172670 76764
rect 173526 76752 173532 76764
rect 172664 76724 173532 76752
rect 172664 76712 172670 76724
rect 173526 76712 173532 76724
rect 173584 76752 173590 76764
rect 206278 76752 206284 76764
rect 173584 76724 206284 76752
rect 173584 76712 173590 76724
rect 206278 76712 206284 76724
rect 206336 76712 206342 76764
rect 218422 76712 218428 76764
rect 218480 76752 218486 76764
rect 289814 76752 289820 76764
rect 218480 76724 289820 76752
rect 218480 76712 218486 76724
rect 289814 76712 289820 76724
rect 289872 76712 289878 76764
rect 148962 76644 148968 76696
rect 149020 76684 149026 76696
rect 182818 76684 182824 76696
rect 149020 76656 182824 76684
rect 149020 76644 149026 76656
rect 182818 76644 182824 76656
rect 182876 76644 182882 76696
rect 218054 76644 218060 76696
rect 218112 76684 218118 76696
rect 218606 76684 218612 76696
rect 218112 76656 218612 76684
rect 218112 76644 218118 76656
rect 218606 76644 218612 76656
rect 218664 76684 218670 76696
rect 296714 76684 296720 76696
rect 218664 76656 296720 76684
rect 218664 76644 218670 76656
rect 296714 76644 296720 76656
rect 296772 76644 296778 76696
rect 149238 76616 149244 76628
rect 147646 76588 149244 76616
rect 149238 76576 149244 76588
rect 149296 76616 149302 76628
rect 150342 76616 150348 76628
rect 149296 76588 150348 76616
rect 149296 76576 149302 76588
rect 150342 76576 150348 76588
rect 150400 76576 150406 76628
rect 151446 76576 151452 76628
rect 151504 76616 151510 76628
rect 197998 76616 198004 76628
rect 151504 76588 198004 76616
rect 151504 76576 151510 76588
rect 197998 76576 198004 76588
rect 198056 76576 198062 76628
rect 218882 76576 218888 76628
rect 218940 76616 218946 76628
rect 353294 76616 353300 76628
rect 218940 76588 353300 76616
rect 218940 76576 218946 76588
rect 353294 76576 353300 76588
rect 353352 76576 353358 76628
rect 67634 76508 67640 76560
rect 67692 76548 67698 76560
rect 105354 76548 105360 76560
rect 67692 76520 105360 76548
rect 67692 76508 67698 76520
rect 105354 76508 105360 76520
rect 105412 76508 105418 76560
rect 111242 76508 111248 76560
rect 111300 76548 111306 76560
rect 111300 76520 133184 76548
rect 111300 76508 111306 76520
rect 113266 76440 113272 76492
rect 113324 76480 113330 76492
rect 113324 76452 133092 76480
rect 113324 76440 113330 76452
rect 112622 76372 112628 76424
rect 112680 76412 112686 76424
rect 129918 76412 129924 76424
rect 112680 76384 129924 76412
rect 112680 76372 112686 76384
rect 129918 76372 129924 76384
rect 129976 76412 129982 76424
rect 130838 76412 130844 76424
rect 129976 76384 130844 76412
rect 129976 76372 129982 76384
rect 130838 76372 130844 76384
rect 130896 76372 130902 76424
rect 125594 76304 125600 76356
rect 125652 76344 125658 76356
rect 133064 76344 133092 76452
rect 133156 76412 133184 76520
rect 134426 76508 134432 76560
rect 134484 76548 134490 76560
rect 134886 76548 134892 76560
rect 134484 76520 134892 76548
rect 134484 76508 134490 76520
rect 134886 76508 134892 76520
rect 134944 76508 134950 76560
rect 143350 76508 143356 76560
rect 143408 76548 143414 76560
rect 146294 76548 146300 76560
rect 143408 76520 146300 76548
rect 143408 76508 143414 76520
rect 146294 76508 146300 76520
rect 146352 76508 146358 76560
rect 146570 76508 146576 76560
rect 146628 76548 146634 76560
rect 182174 76548 182180 76560
rect 146628 76520 182180 76548
rect 146628 76508 146634 76520
rect 182174 76508 182180 76520
rect 182232 76508 182238 76560
rect 196158 76508 196164 76560
rect 196216 76548 196222 76560
rect 196802 76548 196808 76560
rect 196216 76520 196808 76548
rect 196216 76508 196222 76520
rect 196802 76508 196808 76520
rect 196860 76548 196866 76560
rect 389174 76548 389180 76560
rect 196860 76520 389180 76548
rect 196860 76508 196866 76520
rect 389174 76508 389180 76520
rect 389232 76508 389238 76560
rect 145558 76440 145564 76492
rect 145616 76480 145622 76492
rect 146018 76480 146024 76492
rect 145616 76452 146024 76480
rect 145616 76440 145622 76452
rect 146018 76440 146024 76452
rect 146076 76440 146082 76492
rect 147214 76440 147220 76492
rect 147272 76480 147278 76492
rect 178678 76480 178684 76492
rect 147272 76452 178684 76480
rect 147272 76440 147278 76452
rect 178678 76440 178684 76452
rect 178736 76440 178742 76492
rect 140682 76412 140688 76424
rect 133156 76384 140688 76412
rect 140682 76372 140688 76384
rect 140740 76372 140746 76424
rect 163682 76372 163688 76424
rect 163740 76412 163746 76424
rect 171778 76412 171784 76424
rect 163740 76384 171784 76412
rect 163740 76372 163746 76384
rect 171778 76372 171784 76384
rect 171836 76372 171842 76424
rect 173434 76372 173440 76424
rect 173492 76412 173498 76424
rect 173710 76412 173716 76424
rect 173492 76384 173716 76412
rect 173492 76372 173498 76384
rect 173710 76372 173716 76384
rect 173768 76372 173774 76424
rect 174170 76372 174176 76424
rect 174228 76412 174234 76424
rect 177666 76412 177672 76424
rect 174228 76384 177672 76412
rect 174228 76372 174234 76384
rect 177666 76372 177672 76384
rect 177724 76372 177730 76424
rect 177850 76372 177856 76424
rect 177908 76412 177914 76424
rect 199286 76412 199292 76424
rect 177908 76384 199292 76412
rect 177908 76372 177914 76384
rect 199286 76372 199292 76384
rect 199344 76372 199350 76424
rect 139670 76344 139676 76356
rect 125652 76316 128354 76344
rect 133064 76316 139676 76344
rect 125652 76304 125658 76316
rect 128326 76208 128354 76316
rect 139670 76304 139676 76316
rect 139728 76304 139734 76356
rect 145374 76304 145380 76356
rect 145432 76344 145438 76356
rect 145558 76344 145564 76356
rect 145432 76316 145564 76344
rect 145432 76304 145438 76316
rect 145558 76304 145564 76316
rect 145616 76304 145622 76356
rect 152366 76304 152372 76356
rect 152424 76344 152430 76356
rect 152826 76344 152832 76356
rect 152424 76316 152832 76344
rect 152424 76304 152430 76316
rect 152826 76304 152832 76316
rect 152884 76304 152890 76356
rect 170582 76304 170588 76356
rect 170640 76344 170646 76356
rect 170766 76344 170772 76356
rect 170640 76316 170772 76344
rect 170640 76304 170646 76316
rect 170766 76304 170772 76316
rect 170824 76304 170830 76356
rect 176378 76304 176384 76356
rect 176436 76344 176442 76356
rect 180426 76344 180432 76356
rect 176436 76316 180432 76344
rect 176436 76304 176442 76316
rect 180426 76304 180432 76316
rect 180484 76304 180490 76356
rect 195698 76344 195704 76356
rect 183526 76316 195704 76344
rect 170122 76236 170128 76288
rect 170180 76276 170186 76288
rect 177850 76276 177856 76288
rect 170180 76248 177856 76276
rect 170180 76236 170186 76248
rect 177850 76236 177856 76248
rect 177908 76236 177914 76288
rect 131022 76208 131028 76220
rect 128326 76180 131028 76208
rect 131022 76168 131028 76180
rect 131080 76168 131086 76220
rect 150618 76168 150624 76220
rect 150676 76208 150682 76220
rect 150986 76208 150992 76220
rect 150676 76180 150992 76208
rect 150676 76168 150682 76180
rect 150986 76168 150992 76180
rect 151044 76168 151050 76220
rect 172698 76168 172704 76220
rect 172756 76208 172762 76220
rect 173618 76208 173624 76220
rect 172756 76180 173624 76208
rect 172756 76168 172762 76180
rect 173618 76168 173624 76180
rect 173676 76168 173682 76220
rect 174170 76168 174176 76220
rect 174228 76208 174234 76220
rect 175182 76208 175188 76220
rect 174228 76180 175188 76208
rect 174228 76168 174234 76180
rect 175182 76168 175188 76180
rect 175240 76168 175246 76220
rect 183526 76208 183554 76316
rect 195698 76304 195704 76316
rect 195756 76304 195762 76356
rect 175292 76180 183554 76208
rect 163222 76100 163228 76152
rect 163280 76140 163286 76152
rect 163406 76140 163412 76152
rect 163280 76112 163412 76140
rect 163280 76100 163286 76112
rect 163406 76100 163412 76112
rect 163464 76100 163470 76152
rect 170766 76100 170772 76152
rect 170824 76140 170830 76152
rect 175292 76140 175320 76180
rect 170824 76112 175320 76140
rect 170824 76100 170830 76112
rect 175826 76100 175832 76152
rect 175884 76140 175890 76152
rect 176102 76140 176108 76152
rect 175884 76112 176108 76140
rect 175884 76100 175890 76112
rect 176102 76100 176108 76112
rect 176160 76100 176166 76152
rect 101306 76032 101312 76084
rect 101364 76072 101370 76084
rect 101490 76072 101496 76084
rect 101364 76044 101496 76072
rect 101364 76032 101370 76044
rect 101490 76032 101496 76044
rect 101548 76032 101554 76084
rect 136634 76032 136640 76084
rect 136692 76072 136698 76084
rect 137370 76072 137376 76084
rect 136692 76044 137376 76072
rect 136692 76032 136698 76044
rect 137370 76032 137376 76044
rect 137428 76032 137434 76084
rect 132770 75964 132776 76016
rect 132828 76004 132834 76016
rect 133506 76004 133512 76016
rect 132828 75976 133512 76004
rect 132828 75964 132834 75976
rect 133506 75964 133512 75976
rect 133564 75964 133570 76016
rect 138014 75964 138020 76016
rect 138072 76004 138078 76016
rect 138750 76004 138756 76016
rect 138072 75976 138756 76004
rect 138072 75964 138078 75976
rect 138750 75964 138756 75976
rect 138808 75964 138814 76016
rect 165982 75964 165988 76016
rect 166040 76004 166046 76016
rect 166718 76004 166724 76016
rect 166040 75976 166724 76004
rect 166040 75964 166046 75976
rect 166718 75964 166724 75976
rect 166776 75964 166782 76016
rect 88978 75896 88984 75948
rect 89036 75936 89042 75948
rect 96154 75936 96160 75948
rect 89036 75908 96160 75936
rect 89036 75896 89042 75908
rect 96154 75896 96160 75908
rect 96212 75896 96218 75948
rect 99926 75896 99932 75948
rect 99984 75936 99990 75948
rect 100478 75936 100484 75948
rect 99984 75908 100484 75936
rect 99984 75896 99990 75908
rect 100478 75896 100484 75908
rect 100536 75896 100542 75948
rect 121454 75896 121460 75948
rect 121512 75936 121518 75948
rect 123754 75936 123760 75948
rect 121512 75908 123760 75936
rect 121512 75896 121518 75908
rect 123754 75896 123760 75908
rect 123812 75896 123818 75948
rect 135530 75896 135536 75948
rect 135588 75936 135594 75948
rect 136450 75936 136456 75948
rect 135588 75908 136456 75936
rect 135588 75896 135594 75908
rect 136450 75896 136456 75908
rect 136508 75896 136514 75948
rect 138474 75896 138480 75948
rect 138532 75936 138538 75948
rect 138842 75936 138848 75948
rect 138532 75908 138848 75936
rect 138532 75896 138538 75908
rect 138842 75896 138848 75908
rect 138900 75896 138906 75948
rect 143442 75896 143448 75948
rect 143500 75936 143506 75948
rect 145374 75936 145380 75948
rect 143500 75908 145380 75936
rect 143500 75896 143506 75908
rect 145374 75896 145380 75908
rect 145432 75936 145438 75948
rect 152458 75936 152464 75948
rect 145432 75908 152464 75936
rect 145432 75896 145438 75908
rect 152458 75896 152464 75908
rect 152516 75896 152522 75948
rect 160738 75896 160744 75948
rect 160796 75936 160802 75948
rect 161382 75936 161388 75948
rect 160796 75908 161388 75936
rect 160796 75896 160802 75908
rect 161382 75896 161388 75908
rect 161440 75896 161446 75948
rect 164786 75896 164792 75948
rect 164844 75936 164850 75948
rect 165062 75936 165068 75948
rect 164844 75908 165068 75936
rect 164844 75896 164850 75908
rect 165062 75896 165068 75908
rect 165120 75896 165126 75948
rect 168466 75896 168472 75948
rect 168524 75936 168530 75948
rect 168834 75936 168840 75948
rect 168524 75908 168840 75936
rect 168524 75896 168530 75908
rect 168834 75896 168840 75908
rect 168892 75896 168898 75948
rect 172238 75896 172244 75948
rect 172296 75936 172302 75948
rect 172422 75936 172428 75948
rect 172296 75908 172428 75936
rect 172296 75896 172302 75908
rect 172422 75896 172428 75908
rect 172480 75896 172486 75948
rect 176930 75896 176936 75948
rect 176988 75936 176994 75948
rect 177942 75936 177948 75948
rect 176988 75908 177948 75936
rect 176988 75896 176994 75908
rect 177942 75896 177948 75908
rect 178000 75896 178006 75948
rect 97350 75828 97356 75880
rect 97408 75868 97414 75880
rect 132034 75868 132040 75880
rect 97408 75840 132040 75868
rect 97408 75828 97414 75840
rect 132034 75828 132040 75840
rect 132092 75828 132098 75880
rect 137370 75828 137376 75880
rect 137428 75868 137434 75880
rect 137738 75868 137744 75880
rect 137428 75840 137744 75868
rect 137428 75828 137434 75840
rect 137738 75828 137744 75840
rect 137796 75828 137802 75880
rect 158070 75828 158076 75880
rect 158128 75868 158134 75880
rect 206462 75868 206468 75880
rect 158128 75840 206468 75868
rect 158128 75828 158134 75840
rect 206462 75828 206468 75840
rect 206520 75828 206526 75880
rect 98822 75760 98828 75812
rect 98880 75800 98886 75812
rect 145834 75800 145840 75812
rect 98880 75772 145840 75800
rect 98880 75760 98886 75772
rect 145834 75760 145840 75772
rect 145892 75760 145898 75812
rect 163130 75760 163136 75812
rect 163188 75800 163194 75812
rect 163314 75800 163320 75812
rect 163188 75772 163320 75800
rect 163188 75760 163194 75772
rect 163314 75760 163320 75772
rect 163372 75760 163378 75812
rect 170950 75760 170956 75812
rect 171008 75800 171014 75812
rect 202230 75800 202236 75812
rect 171008 75772 202236 75800
rect 171008 75760 171014 75772
rect 202230 75760 202236 75772
rect 202288 75800 202294 75812
rect 202782 75800 202788 75812
rect 202288 75772 202788 75800
rect 202288 75760 202294 75772
rect 202782 75760 202788 75772
rect 202840 75760 202846 75812
rect 96062 75692 96068 75744
rect 96120 75732 96126 75744
rect 99374 75732 99380 75744
rect 96120 75704 99380 75732
rect 96120 75692 96126 75704
rect 99374 75692 99380 75704
rect 99432 75732 99438 75744
rect 100478 75732 100484 75744
rect 99432 75704 100484 75732
rect 99432 75692 99438 75704
rect 100478 75692 100484 75704
rect 100536 75692 100542 75744
rect 104158 75692 104164 75744
rect 104216 75732 104222 75744
rect 137830 75732 137836 75744
rect 104216 75704 137836 75732
rect 104216 75692 104222 75704
rect 137830 75692 137836 75704
rect 137888 75692 137894 75744
rect 172330 75692 172336 75744
rect 172388 75732 172394 75744
rect 205542 75732 205548 75744
rect 172388 75704 205548 75732
rect 172388 75692 172394 75704
rect 205542 75692 205548 75704
rect 205600 75732 205606 75744
rect 206370 75732 206376 75744
rect 205600 75704 206376 75732
rect 205600 75692 205606 75704
rect 206370 75692 206376 75704
rect 206428 75692 206434 75744
rect 113082 75624 113088 75676
rect 113140 75664 113146 75676
rect 147490 75664 147496 75676
rect 113140 75636 147496 75664
rect 113140 75624 113146 75636
rect 147490 75624 147496 75636
rect 147548 75624 147554 75676
rect 157886 75624 157892 75676
rect 157944 75664 157950 75676
rect 157944 75636 166994 75664
rect 157944 75624 157950 75636
rect 139210 75596 139216 75608
rect 109006 75568 139216 75596
rect 89714 75420 89720 75472
rect 89772 75460 89778 75472
rect 104342 75460 104348 75472
rect 89772 75432 104348 75460
rect 89772 75420 89778 75432
rect 104342 75420 104348 75432
rect 104400 75460 104406 75472
rect 109006 75460 109034 75568
rect 139210 75556 139216 75568
rect 139268 75556 139274 75608
rect 163314 75556 163320 75608
rect 163372 75596 163378 75608
rect 163774 75596 163780 75608
rect 163372 75568 163780 75596
rect 163372 75556 163378 75568
rect 163774 75556 163780 75568
rect 163832 75556 163838 75608
rect 166966 75596 166994 75636
rect 168742 75624 168748 75676
rect 168800 75664 168806 75676
rect 169570 75664 169576 75676
rect 168800 75636 169576 75664
rect 168800 75624 168806 75636
rect 169570 75624 169576 75636
rect 169628 75624 169634 75676
rect 171870 75624 171876 75676
rect 171928 75664 171934 75676
rect 206278 75664 206284 75676
rect 171928 75636 206284 75664
rect 171928 75624 171934 75636
rect 206278 75624 206284 75636
rect 206336 75624 206342 75676
rect 192294 75596 192300 75608
rect 166966 75568 192300 75596
rect 192294 75556 192300 75568
rect 192352 75556 192358 75608
rect 119338 75488 119344 75540
rect 119396 75528 119402 75540
rect 152274 75528 152280 75540
rect 119396 75500 152280 75528
rect 119396 75488 119402 75500
rect 152274 75488 152280 75500
rect 152332 75528 152338 75540
rect 152642 75528 152648 75540
rect 152332 75500 152648 75528
rect 152332 75488 152338 75500
rect 152642 75488 152648 75500
rect 152700 75488 152706 75540
rect 161474 75488 161480 75540
rect 161532 75528 161538 75540
rect 162394 75528 162400 75540
rect 161532 75500 162400 75528
rect 161532 75488 161538 75500
rect 162394 75488 162400 75500
rect 162452 75488 162458 75540
rect 170858 75488 170864 75540
rect 170916 75528 170922 75540
rect 204530 75528 204536 75540
rect 170916 75500 204536 75528
rect 170916 75488 170922 75500
rect 204530 75488 204536 75500
rect 204588 75488 204594 75540
rect 104400 75432 109034 75460
rect 104400 75420 104406 75432
rect 112990 75420 112996 75472
rect 113048 75460 113054 75472
rect 145742 75460 145748 75472
rect 113048 75432 145748 75460
rect 113048 75420 113054 75432
rect 145742 75420 145748 75432
rect 145800 75420 145806 75472
rect 150894 75420 150900 75472
rect 150952 75460 150958 75472
rect 151262 75460 151268 75472
rect 150952 75432 151268 75460
rect 150952 75420 150958 75432
rect 151262 75420 151268 75432
rect 151320 75420 151326 75472
rect 168742 75420 168748 75472
rect 168800 75460 168806 75472
rect 169478 75460 169484 75472
rect 168800 75432 169484 75460
rect 168800 75420 168806 75432
rect 169478 75420 169484 75432
rect 169536 75420 169542 75472
rect 169846 75420 169852 75472
rect 169904 75460 169910 75472
rect 171042 75460 171048 75472
rect 169904 75432 171048 75460
rect 169904 75420 169910 75432
rect 171042 75420 171048 75432
rect 171100 75420 171106 75472
rect 171410 75420 171416 75472
rect 171468 75460 171474 75472
rect 172054 75460 172060 75472
rect 171468 75432 172060 75460
rect 171468 75420 171474 75432
rect 172054 75420 172060 75432
rect 172112 75420 172118 75472
rect 172790 75420 172796 75472
rect 172848 75460 172854 75472
rect 173802 75460 173808 75472
rect 172848 75432 173808 75460
rect 172848 75420 172854 75432
rect 173802 75420 173808 75432
rect 173860 75420 173866 75472
rect 174630 75420 174636 75472
rect 174688 75460 174694 75472
rect 207290 75460 207296 75472
rect 174688 75432 207296 75460
rect 174688 75420 174694 75432
rect 207290 75420 207296 75432
rect 207348 75420 207354 75472
rect 84166 75364 99374 75392
rect 52454 75148 52460 75200
rect 52512 75188 52518 75200
rect 84166 75188 84194 75364
rect 52512 75160 84194 75188
rect 99346 75188 99374 75364
rect 100294 75352 100300 75404
rect 100352 75392 100358 75404
rect 100352 75364 107700 75392
rect 100352 75352 100358 75364
rect 100478 75284 100484 75336
rect 100536 75324 100542 75336
rect 107672 75324 107700 75364
rect 107746 75352 107752 75404
rect 107804 75392 107810 75404
rect 136542 75392 136548 75404
rect 107804 75364 136548 75392
rect 107804 75352 107810 75364
rect 136542 75352 136548 75364
rect 136600 75352 136606 75404
rect 150342 75352 150348 75404
rect 150400 75392 150406 75404
rect 150400 75364 157334 75392
rect 150400 75352 150406 75364
rect 131114 75324 131120 75336
rect 100536 75296 107608 75324
rect 107672 75296 131120 75324
rect 100536 75284 100542 75296
rect 107010 75216 107016 75268
rect 107068 75256 107074 75268
rect 107470 75256 107476 75268
rect 107068 75228 107476 75256
rect 107068 75216 107074 75228
rect 107470 75216 107476 75228
rect 107528 75216 107534 75268
rect 107580 75256 107608 75296
rect 131114 75284 131120 75296
rect 131172 75324 131178 75336
rect 133782 75324 133788 75336
rect 131172 75296 133788 75324
rect 131172 75284 131178 75296
rect 133782 75284 133788 75296
rect 133840 75284 133846 75336
rect 139946 75324 139952 75336
rect 137986 75296 139952 75324
rect 137986 75256 138014 75296
rect 139946 75284 139952 75296
rect 140004 75284 140010 75336
rect 140774 75284 140780 75336
rect 140832 75324 140838 75336
rect 141970 75324 141976 75336
rect 140832 75296 141976 75324
rect 140832 75284 140838 75296
rect 141970 75284 141976 75296
rect 142028 75284 142034 75336
rect 150802 75284 150808 75336
rect 150860 75324 150866 75336
rect 151262 75324 151268 75336
rect 150860 75296 151268 75324
rect 150860 75284 150866 75296
rect 151262 75284 151268 75296
rect 151320 75284 151326 75336
rect 157306 75324 157334 75364
rect 158898 75352 158904 75404
rect 158956 75392 158962 75404
rect 159450 75392 159456 75404
rect 158956 75364 159456 75392
rect 158956 75352 158962 75364
rect 159450 75352 159456 75364
rect 159508 75352 159514 75404
rect 160186 75352 160192 75404
rect 160244 75392 160250 75404
rect 160922 75392 160928 75404
rect 160244 75364 160928 75392
rect 160244 75352 160250 75364
rect 160922 75352 160928 75364
rect 160980 75352 160986 75404
rect 178126 75352 178132 75404
rect 178184 75392 178190 75404
rect 205910 75392 205916 75404
rect 178184 75364 205916 75392
rect 178184 75352 178190 75364
rect 205910 75352 205916 75364
rect 205968 75352 205974 75404
rect 216766 75324 216772 75336
rect 157306 75296 216772 75324
rect 216766 75284 216772 75296
rect 216824 75284 216830 75336
rect 107580 75228 138014 75256
rect 138290 75216 138296 75268
rect 138348 75256 138354 75268
rect 138842 75256 138848 75268
rect 138348 75228 138848 75256
rect 138348 75216 138354 75228
rect 138842 75216 138848 75228
rect 138900 75216 138906 75268
rect 139762 75216 139768 75268
rect 139820 75256 139826 75268
rect 140314 75256 140320 75268
rect 139820 75228 140320 75256
rect 139820 75216 139826 75228
rect 140314 75216 140320 75228
rect 140372 75216 140378 75268
rect 142890 75216 142896 75268
rect 142948 75256 142954 75268
rect 143258 75256 143264 75268
rect 142948 75228 143264 75256
rect 142948 75216 142954 75228
rect 143258 75216 143264 75228
rect 143316 75216 143322 75268
rect 146662 75216 146668 75268
rect 146720 75256 146726 75268
rect 176286 75256 176292 75268
rect 146720 75228 176292 75256
rect 146720 75216 146726 75228
rect 176286 75216 176292 75228
rect 176344 75216 176350 75268
rect 202782 75216 202788 75268
rect 202840 75256 202846 75268
rect 454678 75256 454684 75268
rect 202840 75228 454684 75256
rect 202840 75216 202846 75228
rect 454678 75216 454684 75228
rect 454736 75216 454742 75268
rect 102870 75188 102876 75200
rect 99346 75160 102876 75188
rect 52512 75148 52518 75160
rect 102870 75148 102876 75160
rect 102928 75188 102934 75200
rect 107746 75188 107752 75200
rect 102928 75160 107752 75188
rect 102928 75148 102934 75160
rect 107746 75148 107752 75160
rect 107804 75148 107810 75200
rect 117130 75148 117136 75200
rect 117188 75188 117194 75200
rect 145926 75188 145932 75200
rect 117188 75160 145932 75188
rect 117188 75148 117194 75160
rect 145926 75148 145932 75160
rect 145984 75148 145990 75200
rect 176194 75188 176200 75200
rect 157306 75160 176200 75188
rect 123110 75080 123116 75132
rect 123168 75120 123174 75132
rect 123168 75092 147904 75120
rect 123168 75080 123174 75092
rect 108482 75012 108488 75064
rect 108540 75052 108546 75064
rect 130010 75052 130016 75064
rect 108540 75024 130016 75052
rect 108540 75012 108546 75024
rect 130010 75012 130016 75024
rect 130068 75052 130074 75064
rect 137922 75052 137928 75064
rect 130068 75024 137928 75052
rect 130068 75012 130074 75024
rect 137922 75012 137928 75024
rect 137980 75012 137986 75064
rect 135990 74944 135996 74996
rect 136048 74984 136054 74996
rect 136266 74984 136272 74996
rect 136048 74956 136272 74984
rect 136048 74944 136054 74956
rect 136266 74944 136272 74956
rect 136324 74944 136330 74996
rect 147876 74984 147904 75092
rect 148042 75080 148048 75132
rect 148100 75120 148106 75132
rect 157306 75120 157334 75160
rect 176194 75148 176200 75160
rect 176252 75148 176258 75200
rect 177298 75148 177304 75200
rect 177356 75188 177362 75200
rect 201954 75188 201960 75200
rect 177356 75160 201960 75188
rect 177356 75148 177362 75160
rect 201954 75148 201960 75160
rect 202012 75148 202018 75200
rect 205910 75148 205916 75200
rect 205968 75188 205974 75200
rect 499574 75188 499580 75200
rect 205968 75160 499580 75188
rect 205968 75148 205974 75160
rect 499574 75148 499580 75160
rect 499632 75148 499638 75200
rect 148100 75092 157334 75120
rect 148100 75080 148106 75092
rect 157426 75080 157432 75132
rect 157484 75120 157490 75132
rect 158622 75120 158628 75132
rect 157484 75092 158628 75120
rect 157484 75080 157490 75092
rect 158622 75080 158628 75092
rect 158680 75080 158686 75132
rect 159082 75080 159088 75132
rect 159140 75120 159146 75132
rect 159634 75120 159640 75132
rect 159140 75092 159640 75120
rect 159140 75080 159146 75092
rect 159634 75080 159640 75092
rect 159692 75080 159698 75132
rect 160186 75080 160192 75132
rect 160244 75120 160250 75132
rect 160554 75120 160560 75132
rect 160244 75092 160560 75120
rect 160244 75080 160250 75092
rect 160554 75080 160560 75092
rect 160612 75080 160618 75132
rect 160646 75080 160652 75132
rect 160704 75120 160710 75132
rect 161198 75120 161204 75132
rect 160704 75092 161204 75120
rect 160704 75080 160710 75092
rect 161198 75080 161204 75092
rect 161256 75080 161262 75132
rect 169018 75080 169024 75132
rect 169076 75120 169082 75132
rect 176378 75120 176384 75132
rect 169076 75092 176384 75120
rect 169076 75080 169082 75092
rect 176378 75080 176384 75092
rect 176436 75080 176442 75132
rect 180334 75080 180340 75132
rect 180392 75120 180398 75132
rect 219894 75120 219900 75132
rect 180392 75092 219900 75120
rect 180392 75080 180398 75092
rect 219894 75080 219900 75092
rect 219952 75080 219958 75132
rect 166718 75052 166724 75064
rect 157306 75024 166724 75052
rect 153746 74984 153752 74996
rect 147876 74956 153752 74984
rect 153746 74944 153752 74956
rect 153804 74944 153810 74996
rect 146386 74808 146392 74860
rect 146444 74848 146450 74860
rect 157306 74848 157334 75024
rect 166718 75012 166724 75024
rect 166776 75012 166782 75064
rect 172882 75012 172888 75064
rect 172940 75052 172946 75064
rect 173802 75052 173808 75064
rect 172940 75024 173808 75052
rect 172940 75012 172946 75024
rect 173802 75012 173808 75024
rect 173860 75012 173866 75064
rect 176286 75012 176292 75064
rect 176344 75052 176350 75064
rect 176344 75024 176700 75052
rect 176344 75012 176350 75024
rect 157886 74944 157892 74996
rect 157944 74984 157950 74996
rect 158622 74984 158628 74996
rect 157944 74956 158628 74984
rect 157944 74944 157950 74956
rect 158622 74944 158628 74956
rect 158680 74944 158686 74996
rect 168466 74944 168472 74996
rect 168524 74984 168530 74996
rect 169386 74984 169392 74996
rect 168524 74956 169392 74984
rect 168524 74944 168530 74956
rect 169386 74944 169392 74956
rect 169444 74944 169450 74996
rect 176672 74984 176700 75024
rect 183554 75012 183560 75064
rect 183612 75052 183618 75064
rect 184842 75052 184848 75064
rect 183612 75024 184848 75052
rect 183612 75012 183618 75024
rect 184842 75012 184848 75024
rect 184900 75052 184906 75064
rect 210602 75052 210608 75064
rect 184900 75024 210608 75052
rect 184900 75012 184906 75024
rect 210602 75012 210608 75024
rect 210660 75012 210666 75064
rect 185026 74984 185032 74996
rect 176672 74956 185032 74984
rect 185026 74944 185032 74956
rect 185084 74944 185090 74996
rect 161198 74876 161204 74928
rect 161256 74916 161262 74928
rect 169018 74916 169024 74928
rect 161256 74888 169024 74916
rect 161256 74876 161262 74888
rect 169018 74876 169024 74888
rect 169076 74876 169082 74928
rect 175550 74876 175556 74928
rect 175608 74916 175614 74928
rect 176286 74916 176292 74928
rect 175608 74888 176292 74916
rect 175608 74876 175614 74888
rect 176286 74876 176292 74888
rect 176344 74876 176350 74928
rect 146444 74820 157334 74848
rect 146444 74808 146450 74820
rect 162302 74808 162308 74860
rect 162360 74848 162366 74860
rect 162670 74848 162676 74860
rect 162360 74820 162676 74848
rect 162360 74808 162366 74820
rect 162670 74808 162676 74820
rect 162728 74808 162734 74860
rect 154666 74672 154672 74724
rect 154724 74712 154730 74724
rect 155310 74712 155316 74724
rect 154724 74684 155316 74712
rect 154724 74672 154730 74684
rect 155310 74672 155316 74684
rect 155368 74672 155374 74724
rect 166718 74672 166724 74724
rect 166776 74712 166782 74724
rect 180794 74712 180800 74724
rect 166776 74684 180800 74712
rect 166776 74672 166782 74684
rect 180794 74672 180800 74684
rect 180852 74672 180858 74724
rect 149698 74604 149704 74656
rect 149756 74644 149762 74656
rect 150250 74644 150256 74656
rect 149756 74616 150256 74644
rect 149756 74604 149762 74616
rect 150250 74604 150256 74616
rect 150308 74604 150314 74656
rect 206278 74604 206284 74656
rect 206336 74644 206342 74656
rect 475378 74644 475384 74656
rect 206336 74616 475384 74644
rect 206336 74604 206342 74616
rect 475378 74604 475384 74616
rect 475436 74604 475442 74656
rect 165706 74536 165712 74588
rect 165764 74576 165770 74588
rect 166166 74576 166172 74588
rect 165764 74548 166172 74576
rect 165764 74536 165770 74548
rect 166166 74536 166172 74548
rect 166224 74536 166230 74588
rect 206370 74536 206376 74588
rect 206428 74576 206434 74588
rect 511258 74576 511264 74588
rect 206428 74548 511264 74576
rect 206428 74536 206434 74548
rect 511258 74536 511264 74548
rect 511316 74536 511322 74588
rect 96338 74468 96344 74520
rect 96396 74508 96402 74520
rect 149698 74508 149704 74520
rect 96396 74480 149704 74508
rect 96396 74468 96402 74480
rect 149698 74468 149704 74480
rect 149756 74508 149762 74520
rect 150066 74508 150072 74520
rect 149756 74480 150072 74508
rect 149756 74468 149762 74480
rect 150066 74468 150072 74480
rect 150124 74468 150130 74520
rect 153378 74468 153384 74520
rect 153436 74508 153442 74520
rect 220814 74508 220820 74520
rect 153436 74480 220820 74508
rect 153436 74468 153442 74480
rect 220814 74468 220820 74480
rect 220872 74468 220878 74520
rect 114830 74400 114836 74452
rect 114888 74440 114894 74452
rect 149974 74440 149980 74452
rect 114888 74412 149980 74440
rect 114888 74400 114894 74412
rect 149974 74400 149980 74412
rect 150032 74400 150038 74452
rect 159266 74400 159272 74452
rect 159324 74440 159330 74452
rect 159910 74440 159916 74452
rect 159324 74412 159916 74440
rect 159324 74400 159330 74412
rect 159910 74400 159916 74412
rect 159968 74400 159974 74452
rect 161842 74400 161848 74452
rect 161900 74440 161906 74452
rect 218238 74440 218244 74452
rect 161900 74412 218244 74440
rect 161900 74400 161906 74412
rect 218238 74400 218244 74412
rect 218296 74400 218302 74452
rect 122374 74332 122380 74384
rect 122432 74372 122438 74384
rect 151538 74372 151544 74384
rect 122432 74344 151544 74372
rect 122432 74332 122438 74344
rect 151538 74332 151544 74344
rect 151596 74332 151602 74384
rect 155862 74332 155868 74384
rect 155920 74372 155926 74384
rect 189810 74372 189816 74384
rect 155920 74344 189816 74372
rect 155920 74332 155926 74344
rect 189810 74332 189816 74344
rect 189868 74332 189874 74384
rect 98914 74264 98920 74316
rect 98972 74304 98978 74316
rect 132954 74304 132960 74316
rect 98972 74276 132960 74304
rect 98972 74264 98978 74276
rect 132954 74264 132960 74276
rect 133012 74264 133018 74316
rect 166258 74264 166264 74316
rect 166316 74304 166322 74316
rect 166902 74304 166908 74316
rect 166316 74276 166908 74304
rect 166316 74264 166322 74276
rect 166902 74264 166908 74276
rect 166960 74304 166966 74316
rect 200758 74304 200764 74316
rect 166960 74276 200764 74304
rect 166960 74264 166966 74276
rect 200758 74264 200764 74276
rect 200816 74264 200822 74316
rect 119246 74196 119252 74248
rect 119304 74236 119310 74248
rect 151814 74236 151820 74248
rect 119304 74208 151820 74236
rect 119304 74196 119310 74208
rect 151814 74196 151820 74208
rect 151872 74196 151878 74248
rect 172422 74196 172428 74248
rect 172480 74236 172486 74248
rect 206094 74236 206100 74248
rect 172480 74208 206100 74236
rect 172480 74196 172486 74208
rect 206094 74196 206100 74208
rect 206152 74196 206158 74248
rect 117958 74128 117964 74180
rect 118016 74168 118022 74180
rect 150894 74168 150900 74180
rect 118016 74140 150900 74168
rect 118016 74128 118022 74140
rect 150894 74128 150900 74140
rect 150952 74168 150958 74180
rect 151630 74168 151636 74180
rect 150952 74140 151636 74168
rect 150952 74128 150958 74140
rect 151630 74128 151636 74140
rect 151688 74128 151694 74180
rect 155586 74128 155592 74180
rect 155644 74168 155650 74180
rect 155862 74168 155868 74180
rect 155644 74140 155868 74168
rect 155644 74128 155650 74140
rect 155862 74128 155868 74140
rect 155920 74128 155926 74180
rect 171042 74128 171048 74180
rect 171100 74168 171106 74180
rect 204438 74168 204444 74180
rect 171100 74140 204444 74168
rect 171100 74128 171106 74140
rect 204438 74128 204444 74140
rect 204496 74128 204502 74180
rect 101490 74060 101496 74112
rect 101548 74100 101554 74112
rect 134978 74100 134984 74112
rect 101548 74072 134984 74100
rect 101548 74060 101554 74072
rect 134978 74060 134984 74072
rect 135036 74060 135042 74112
rect 173802 74060 173808 74112
rect 173860 74100 173866 74112
rect 206186 74100 206192 74112
rect 173860 74072 206192 74100
rect 173860 74060 173866 74072
rect 206186 74060 206192 74072
rect 206244 74060 206250 74112
rect 116762 73992 116768 74044
rect 116820 74032 116826 74044
rect 116820 74004 147674 74032
rect 116820 73992 116826 74004
rect 139394 73964 139400 73976
rect 109006 73936 139400 73964
rect 95970 73856 95976 73908
rect 96028 73896 96034 73908
rect 107102 73896 107108 73908
rect 96028 73868 107108 73896
rect 96028 73856 96034 73868
rect 107102 73856 107108 73868
rect 107160 73896 107166 73908
rect 109006 73896 109034 73936
rect 139394 73924 139400 73936
rect 139452 73924 139458 73976
rect 107160 73868 109034 73896
rect 147646 73896 147674 74004
rect 159910 73992 159916 74044
rect 159968 74032 159974 74044
rect 180058 74032 180064 74044
rect 159968 74004 180064 74032
rect 159968 73992 159974 74004
rect 180058 73992 180064 74004
rect 180116 73992 180122 74044
rect 181990 73992 181996 74044
rect 182048 74032 182054 74044
rect 219710 74032 219716 74044
rect 182048 74004 219716 74032
rect 182048 73992 182054 74004
rect 219710 73992 219716 74004
rect 219768 73992 219774 74044
rect 220814 73992 220820 74044
rect 220872 74032 220878 74044
rect 269114 74032 269120 74044
rect 220872 74004 269120 74032
rect 220872 73992 220878 74004
rect 269114 73992 269120 74004
rect 269172 73992 269178 74044
rect 163038 73924 163044 73976
rect 163096 73964 163102 73976
rect 192202 73964 192208 73976
rect 163096 73936 192208 73964
rect 163096 73924 163102 73936
rect 192202 73924 192208 73936
rect 192260 73964 192266 73976
rect 322934 73964 322940 73976
rect 192260 73936 322940 73964
rect 192260 73924 192266 73936
rect 322934 73924 322940 73936
rect 322992 73924 322998 73976
rect 149882 73896 149888 73908
rect 147646 73868 149888 73896
rect 107160 73856 107166 73868
rect 149882 73856 149888 73868
rect 149940 73896 149946 73908
rect 207658 73896 207664 73908
rect 149940 73868 207664 73896
rect 149940 73856 149946 73868
rect 207658 73856 207664 73868
rect 207716 73856 207722 73908
rect 218238 73856 218244 73908
rect 218296 73896 218302 73908
rect 354674 73896 354680 73908
rect 218296 73868 354680 73896
rect 218296 73856 218302 73868
rect 354674 73856 354680 73868
rect 354732 73856 354738 73908
rect 35894 73788 35900 73840
rect 35952 73828 35958 73840
rect 101490 73828 101496 73840
rect 35952 73800 101496 73828
rect 35952 73788 35958 73800
rect 101490 73788 101496 73800
rect 101548 73788 101554 73840
rect 106274 73788 106280 73840
rect 106332 73828 106338 73840
rect 136358 73828 136364 73840
rect 106332 73800 136364 73828
rect 106332 73788 106338 73800
rect 136358 73788 136364 73800
rect 136416 73788 136422 73840
rect 151538 73788 151544 73840
rect 151596 73828 151602 73840
rect 248414 73828 248420 73840
rect 151596 73800 248420 73828
rect 151596 73788 151602 73800
rect 248414 73788 248420 73800
rect 248472 73788 248478 73840
rect 268378 73788 268384 73840
rect 268436 73828 268442 73840
rect 580994 73828 581000 73840
rect 268436 73800 581000 73828
rect 268436 73788 268442 73800
rect 580994 73788 581000 73800
rect 581052 73788 581058 73840
rect 118050 73720 118056 73772
rect 118108 73760 118114 73772
rect 141510 73760 141516 73772
rect 118108 73732 141516 73760
rect 118108 73720 118114 73732
rect 141510 73720 141516 73732
rect 141568 73720 141574 73772
rect 151814 73720 151820 73772
rect 151872 73760 151878 73772
rect 152918 73760 152924 73772
rect 151872 73732 152924 73760
rect 151872 73720 151878 73732
rect 152918 73720 152924 73732
rect 152976 73720 152982 73772
rect 163038 73720 163044 73772
rect 163096 73760 163102 73772
rect 164142 73760 164148 73772
rect 163096 73732 164148 73760
rect 163096 73720 163102 73732
rect 164142 73720 164148 73732
rect 164200 73720 164206 73772
rect 175182 73720 175188 73772
rect 175240 73760 175246 73772
rect 207566 73760 207572 73772
rect 175240 73732 207572 73760
rect 175240 73720 175246 73732
rect 207566 73720 207572 73732
rect 207624 73720 207630 73772
rect 158070 73652 158076 73704
rect 158128 73692 158134 73704
rect 158438 73692 158444 73704
rect 158128 73664 158444 73692
rect 158128 73652 158134 73664
rect 158438 73652 158444 73664
rect 158496 73652 158502 73704
rect 169202 73652 169208 73704
rect 169260 73692 169266 73704
rect 179046 73692 179052 73704
rect 169260 73664 179052 73692
rect 169260 73652 169266 73664
rect 179046 73652 179052 73664
rect 179104 73692 179110 73704
rect 203150 73692 203156 73704
rect 179104 73664 203156 73692
rect 179104 73652 179110 73664
rect 203150 73652 203156 73664
rect 203208 73652 203214 73704
rect 97626 73584 97632 73636
rect 97684 73624 97690 73636
rect 131482 73624 131488 73636
rect 97684 73596 131488 73624
rect 97684 73584 97690 73596
rect 131482 73584 131488 73596
rect 131540 73624 131546 73636
rect 132310 73624 132316 73636
rect 131540 73596 132316 73624
rect 131540 73584 131546 73596
rect 132310 73584 132316 73596
rect 132368 73584 132374 73636
rect 164050 73584 164056 73636
rect 164108 73624 164114 73636
rect 166258 73624 166264 73636
rect 164108 73596 166264 73624
rect 164108 73584 164114 73596
rect 166258 73584 166264 73596
rect 166316 73584 166322 73636
rect 168282 73584 168288 73636
rect 168340 73624 168346 73636
rect 181990 73624 181996 73636
rect 168340 73596 181996 73624
rect 168340 73584 168346 73596
rect 181990 73584 181996 73596
rect 182048 73584 182054 73636
rect 118510 73516 118516 73568
rect 118568 73556 118574 73568
rect 149790 73556 149796 73568
rect 118568 73528 149796 73556
rect 118568 73516 118574 73528
rect 149790 73516 149796 73528
rect 149848 73516 149854 73568
rect 135806 73380 135812 73432
rect 135864 73420 135870 73432
rect 136174 73420 136180 73432
rect 135864 73392 136180 73420
rect 135864 73380 135870 73392
rect 136174 73380 136180 73392
rect 136232 73380 136238 73432
rect 122098 73176 122104 73228
rect 122156 73216 122162 73228
rect 122834 73216 122840 73228
rect 122156 73188 122840 73216
rect 122156 73176 122162 73188
rect 122834 73176 122840 73188
rect 122892 73176 122898 73228
rect 127710 73108 127716 73160
rect 127768 73148 127774 73160
rect 136634 73148 136640 73160
rect 127768 73120 136640 73148
rect 127768 73108 127774 73120
rect 136634 73108 136640 73120
rect 136692 73108 136698 73160
rect 167638 73108 167644 73160
rect 167696 73148 167702 73160
rect 168282 73148 168288 73160
rect 167696 73120 168288 73148
rect 167696 73108 167702 73120
rect 168282 73108 168288 73120
rect 168340 73148 168346 73160
rect 180702 73148 180708 73160
rect 168340 73120 180708 73148
rect 168340 73108 168346 73120
rect 180702 73108 180708 73120
rect 180760 73108 180766 73160
rect 327718 73108 327724 73160
rect 327776 73148 327782 73160
rect 580166 73148 580172 73160
rect 327776 73120 580172 73148
rect 327776 73108 327782 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 115750 73040 115756 73092
rect 115808 73080 115814 73092
rect 149146 73080 149152 73092
rect 115808 73052 149152 73080
rect 115808 73040 115814 73052
rect 149146 73040 149152 73052
rect 149204 73080 149210 73092
rect 149606 73080 149612 73092
rect 149204 73052 149612 73080
rect 149204 73040 149210 73052
rect 149606 73040 149612 73052
rect 149664 73040 149670 73092
rect 157794 73040 157800 73092
rect 157852 73080 157858 73092
rect 221090 73080 221096 73092
rect 157852 73052 221096 73080
rect 157852 73040 157858 73052
rect 221090 73040 221096 73052
rect 221148 73080 221154 73092
rect 222102 73080 222108 73092
rect 221148 73052 222108 73080
rect 221148 73040 221154 73052
rect 222102 73040 222108 73052
rect 222160 73040 222166 73092
rect 128998 72972 129004 73024
rect 129056 73012 129062 73024
rect 152826 73012 152832 73024
rect 129056 72984 152832 73012
rect 129056 72972 129062 72984
rect 152826 72972 152832 72984
rect 152884 72972 152890 73024
rect 161290 72972 161296 73024
rect 161348 73012 161354 73024
rect 209222 73012 209228 73024
rect 161348 72984 209228 73012
rect 161348 72972 161354 72984
rect 209222 72972 209228 72984
rect 209280 72972 209286 73024
rect 114370 72904 114376 72956
rect 114428 72944 114434 72956
rect 147858 72944 147864 72956
rect 114428 72916 147864 72944
rect 114428 72904 114434 72916
rect 147858 72904 147864 72916
rect 147916 72944 147922 72956
rect 148778 72944 148784 72956
rect 147916 72916 148784 72944
rect 147916 72904 147922 72916
rect 148778 72904 148784 72916
rect 148836 72904 148842 72956
rect 155770 72904 155776 72956
rect 155828 72944 155834 72956
rect 190822 72944 190828 72956
rect 155828 72916 190828 72944
rect 155828 72904 155834 72916
rect 190822 72904 190828 72916
rect 190880 72904 190886 72956
rect 117222 72836 117228 72888
rect 117280 72876 117286 72888
rect 149330 72876 149336 72888
rect 117280 72848 149336 72876
rect 117280 72836 117286 72848
rect 149330 72836 149336 72848
rect 149388 72876 149394 72888
rect 150158 72876 150164 72888
rect 149388 72848 150164 72876
rect 149388 72836 149394 72848
rect 150158 72836 150164 72848
rect 150216 72836 150222 72888
rect 166534 72836 166540 72888
rect 166592 72876 166598 72888
rect 200942 72876 200948 72888
rect 166592 72848 200948 72876
rect 166592 72836 166598 72848
rect 200942 72836 200948 72848
rect 201000 72836 201006 72888
rect 115842 72768 115848 72820
rect 115900 72808 115906 72820
rect 148134 72808 148140 72820
rect 115900 72780 148140 72808
rect 115900 72768 115906 72780
rect 148134 72768 148140 72780
rect 148192 72808 148198 72820
rect 148410 72808 148416 72820
rect 148192 72780 148416 72808
rect 148192 72768 148198 72780
rect 148410 72768 148416 72780
rect 148468 72768 148474 72820
rect 155218 72768 155224 72820
rect 155276 72808 155282 72820
rect 189718 72808 189724 72820
rect 155276 72780 189724 72808
rect 155276 72768 155282 72780
rect 155788 72752 155816 72780
rect 189718 72768 189724 72780
rect 189776 72768 189782 72820
rect 221366 72768 221372 72820
rect 221424 72808 221430 72820
rect 311158 72808 311164 72820
rect 221424 72780 311164 72808
rect 221424 72768 221430 72780
rect 311158 72768 311164 72780
rect 311216 72768 311222 72820
rect 109862 72700 109868 72752
rect 109920 72740 109926 72752
rect 142246 72740 142252 72752
rect 109920 72712 142252 72740
rect 109920 72700 109926 72712
rect 142246 72700 142252 72712
rect 142304 72700 142310 72752
rect 155770 72700 155776 72752
rect 155828 72700 155834 72752
rect 189074 72700 189080 72752
rect 189132 72740 189138 72752
rect 189626 72740 189632 72752
rect 189132 72712 189632 72740
rect 189132 72700 189138 72712
rect 189626 72700 189632 72712
rect 189684 72740 189690 72752
rect 283558 72740 283564 72752
rect 189684 72712 283564 72740
rect 189684 72700 189690 72712
rect 283558 72700 283564 72712
rect 283616 72700 283622 72752
rect 139118 72672 139124 72684
rect 109006 72644 139124 72672
rect 96614 72428 96620 72480
rect 96672 72468 96678 72480
rect 107286 72468 107292 72480
rect 96672 72440 107292 72468
rect 96672 72428 96678 72440
rect 107286 72428 107292 72440
rect 107344 72468 107350 72480
rect 109006 72468 109034 72644
rect 139118 72632 139124 72644
rect 139176 72632 139182 72684
rect 145650 72632 145656 72684
rect 145708 72672 145714 72684
rect 156874 72672 156880 72684
rect 145708 72644 156880 72672
rect 145708 72632 145714 72644
rect 156874 72632 156880 72644
rect 156932 72632 156938 72684
rect 162670 72632 162676 72684
rect 162728 72672 162734 72684
rect 196526 72672 196532 72684
rect 162728 72644 196532 72672
rect 162728 72632 162734 72644
rect 196526 72632 196532 72644
rect 196584 72632 196590 72684
rect 222102 72632 222108 72684
rect 222160 72672 222166 72684
rect 324958 72672 324964 72684
rect 222160 72644 324964 72672
rect 222160 72632 222166 72644
rect 324958 72632 324964 72644
rect 325016 72632 325022 72684
rect 117038 72564 117044 72616
rect 117096 72604 117102 72616
rect 147950 72604 147956 72616
rect 117096 72576 147956 72604
rect 117096 72564 117102 72576
rect 147950 72564 147956 72576
rect 148008 72604 148014 72616
rect 148502 72604 148508 72616
rect 148008 72576 148508 72604
rect 148008 72564 148014 72576
rect 148502 72564 148508 72576
rect 148560 72564 148566 72616
rect 155678 72564 155684 72616
rect 155736 72604 155742 72616
rect 155736 72576 176654 72604
rect 155736 72564 155742 72576
rect 118602 72496 118608 72548
rect 118660 72536 118666 72548
rect 148042 72536 148048 72548
rect 118660 72508 148048 72536
rect 118660 72496 118666 72508
rect 148042 72496 148048 72508
rect 148100 72536 148106 72548
rect 148962 72536 148968 72548
rect 148100 72508 148968 72536
rect 148100 72496 148106 72508
rect 148962 72496 148968 72508
rect 149020 72496 149026 72548
rect 176626 72536 176654 72576
rect 176930 72564 176936 72616
rect 176988 72604 176994 72616
rect 177390 72604 177396 72616
rect 176988 72576 177396 72604
rect 176988 72564 176994 72576
rect 177390 72564 177396 72576
rect 177448 72564 177454 72616
rect 191466 72604 191472 72616
rect 189184 72576 191472 72604
rect 189074 72536 189080 72548
rect 176626 72508 189080 72536
rect 189074 72496 189080 72508
rect 189132 72496 189138 72548
rect 107344 72440 109034 72468
rect 107344 72428 107350 72440
rect 111794 72428 111800 72480
rect 111852 72468 111858 72480
rect 112438 72468 112444 72480
rect 111852 72440 112444 72468
rect 111852 72428 111858 72440
rect 112438 72428 112444 72440
rect 112496 72468 112502 72480
rect 140958 72468 140964 72480
rect 112496 72440 140964 72468
rect 112496 72428 112502 72440
rect 140958 72428 140964 72440
rect 141016 72428 141022 72480
rect 157058 72428 157064 72480
rect 157116 72468 157122 72480
rect 189184 72468 189212 72576
rect 191466 72564 191472 72576
rect 191524 72604 191530 72616
rect 304994 72604 305000 72616
rect 191524 72576 305000 72604
rect 191524 72564 191530 72576
rect 304994 72564 305000 72576
rect 305052 72564 305058 72616
rect 193950 72536 193956 72548
rect 157116 72440 189212 72468
rect 190426 72508 193956 72536
rect 157116 72428 157122 72440
rect 110874 72360 110880 72412
rect 110932 72400 110938 72412
rect 138198 72400 138204 72412
rect 110932 72372 138204 72400
rect 110932 72360 110938 72372
rect 138198 72360 138204 72372
rect 138256 72360 138262 72412
rect 160094 72360 160100 72412
rect 160152 72400 160158 72412
rect 190426 72400 190454 72508
rect 193950 72496 193956 72508
rect 194008 72536 194014 72548
rect 340874 72536 340880 72548
rect 194008 72508 340880 72536
rect 194008 72496 194014 72508
rect 340874 72496 340880 72508
rect 340932 72496 340938 72548
rect 382274 72468 382280 72480
rect 160152 72372 190454 72400
rect 200086 72440 382280 72468
rect 160152 72360 160158 72372
rect 109954 72292 109960 72344
rect 110012 72332 110018 72344
rect 128354 72332 128360 72344
rect 110012 72304 128360 72332
rect 110012 72292 110018 72304
rect 128354 72292 128360 72304
rect 128412 72332 128418 72344
rect 129458 72332 129464 72344
rect 128412 72304 129464 72332
rect 128412 72292 128418 72304
rect 129458 72292 129464 72304
rect 129516 72292 129522 72344
rect 162210 72292 162216 72344
rect 162268 72332 162274 72344
rect 196618 72332 196624 72344
rect 162268 72304 196624 72332
rect 162268 72292 162274 72304
rect 196618 72292 196624 72304
rect 196676 72332 196682 72344
rect 200086 72332 200114 72440
rect 382274 72428 382280 72440
rect 382332 72428 382338 72480
rect 196676 72304 200114 72332
rect 196676 72292 196682 72304
rect 105538 72224 105544 72276
rect 105596 72264 105602 72276
rect 140130 72264 140136 72276
rect 105596 72236 140136 72264
rect 105596 72224 105602 72236
rect 140130 72224 140136 72236
rect 140188 72224 140194 72276
rect 156598 72224 156604 72276
rect 156656 72264 156662 72276
rect 221366 72264 221372 72276
rect 156656 72236 221372 72264
rect 156656 72224 156662 72236
rect 221366 72224 221372 72236
rect 221424 72224 221430 72276
rect 114186 72156 114192 72208
rect 114244 72196 114250 72208
rect 148318 72196 148324 72208
rect 114244 72168 148324 72196
rect 114244 72156 114250 72168
rect 148318 72156 148324 72168
rect 148376 72196 148382 72208
rect 148502 72196 148508 72208
rect 148376 72168 148508 72196
rect 148376 72156 148382 72168
rect 148502 72156 148508 72168
rect 148560 72156 148566 72208
rect 156690 72156 156696 72208
rect 156748 72196 156754 72208
rect 157242 72196 157248 72208
rect 156748 72168 157248 72196
rect 156748 72156 156754 72168
rect 157242 72156 157248 72168
rect 157300 72196 157306 72208
rect 190914 72196 190920 72208
rect 157300 72168 190920 72196
rect 157300 72156 157306 72168
rect 190914 72156 190920 72168
rect 190972 72156 190978 72208
rect 160094 72088 160100 72140
rect 160152 72128 160158 72140
rect 161106 72128 161112 72140
rect 160152 72100 161112 72128
rect 160152 72088 160158 72100
rect 161106 72088 161112 72100
rect 161164 72088 161170 72140
rect 194226 72128 194232 72140
rect 166966 72100 194232 72128
rect 159726 72020 159732 72072
rect 159784 72060 159790 72072
rect 166966 72060 166994 72100
rect 194226 72088 194232 72100
rect 194284 72088 194290 72140
rect 159784 72032 166994 72060
rect 159784 72020 159790 72032
rect 176286 72020 176292 72072
rect 176344 72060 176350 72072
rect 176470 72060 176476 72072
rect 176344 72032 176476 72060
rect 176344 72020 176350 72032
rect 176470 72020 176476 72032
rect 176528 72020 176534 72072
rect 108666 71680 108672 71732
rect 108724 71720 108730 71732
rect 114554 71720 114560 71732
rect 108724 71692 114560 71720
rect 108724 71680 108730 71692
rect 114554 71680 114560 71692
rect 114612 71680 114618 71732
rect 127618 71680 127624 71732
rect 127676 71720 127682 71732
rect 138014 71720 138020 71732
rect 127676 71692 138020 71720
rect 127676 71680 127682 71692
rect 138014 71680 138020 71692
rect 138072 71720 138078 71732
rect 138290 71720 138296 71732
rect 138072 71692 138296 71720
rect 138072 71680 138078 71692
rect 138290 71680 138296 71692
rect 138348 71680 138354 71732
rect 157702 71680 157708 71732
rect 157760 71720 157766 71732
rect 158346 71720 158352 71732
rect 157760 71692 158352 71720
rect 157760 71680 157766 71692
rect 158346 71680 158352 71692
rect 158404 71680 158410 71732
rect 159542 71680 159548 71732
rect 159600 71720 159606 71732
rect 160002 71720 160008 71732
rect 159600 71692 160008 71720
rect 159600 71680 159606 71692
rect 160002 71680 160008 71692
rect 160060 71680 160066 71732
rect 169938 71680 169944 71732
rect 169996 71720 170002 71732
rect 211522 71720 211528 71732
rect 169996 71692 211528 71720
rect 169996 71680 170002 71692
rect 211522 71680 211528 71692
rect 211580 71720 211586 71732
rect 212442 71720 212448 71732
rect 211580 71692 212448 71720
rect 211580 71680 211586 71692
rect 212442 71680 212448 71692
rect 212500 71680 212506 71732
rect 3510 71612 3516 71664
rect 3568 71652 3574 71664
rect 8938 71652 8944 71664
rect 3568 71624 8944 71652
rect 3568 71612 3574 71624
rect 8938 71612 8944 71624
rect 8996 71612 9002 71664
rect 102594 71612 102600 71664
rect 102652 71652 102658 71664
rect 151354 71652 151360 71664
rect 102652 71624 151360 71652
rect 102652 71612 102658 71624
rect 151354 71612 151360 71624
rect 151412 71612 151418 71664
rect 158364 71652 158392 71680
rect 192846 71652 192852 71664
rect 158364 71624 192852 71652
rect 192846 71612 192852 71624
rect 192904 71612 192910 71664
rect 99098 71544 99104 71596
rect 99156 71584 99162 71596
rect 99156 71556 138014 71584
rect 99156 71544 99162 71556
rect 101490 71476 101496 71528
rect 101548 71516 101554 71528
rect 135438 71516 135444 71528
rect 101548 71488 135444 71516
rect 101548 71476 101554 71488
rect 135438 71476 135444 71488
rect 135496 71476 135502 71528
rect 137986 71516 138014 71556
rect 156782 71544 156788 71596
rect 156840 71584 156846 71596
rect 157150 71584 157156 71596
rect 156840 71556 157156 71584
rect 156840 71544 156846 71556
rect 157150 71544 157156 71556
rect 157208 71584 157214 71596
rect 191190 71584 191196 71596
rect 157208 71556 191196 71584
rect 157208 71544 157214 71556
rect 191190 71544 191196 71556
rect 191248 71544 191254 71596
rect 192478 71544 192484 71596
rect 192536 71584 192542 71596
rect 193122 71584 193128 71596
rect 192536 71556 193128 71584
rect 192536 71544 192542 71556
rect 193122 71544 193128 71556
rect 193180 71584 193186 71596
rect 202138 71584 202144 71596
rect 193180 71556 202144 71584
rect 193180 71544 193186 71556
rect 202138 71544 202144 71556
rect 202196 71544 202202 71596
rect 146938 71516 146944 71528
rect 137986 71488 146944 71516
rect 146938 71476 146944 71488
rect 146996 71476 147002 71528
rect 156506 71476 156512 71528
rect 156564 71516 156570 71528
rect 157058 71516 157064 71528
rect 156564 71488 157064 71516
rect 156564 71476 156570 71488
rect 157058 71476 157064 71488
rect 157116 71516 157122 71528
rect 191650 71516 191656 71528
rect 157116 71488 191656 71516
rect 157116 71476 157122 71488
rect 191650 71476 191656 71488
rect 191708 71476 191714 71528
rect 115290 71408 115296 71460
rect 115348 71448 115354 71460
rect 148226 71448 148232 71460
rect 115348 71420 148232 71448
rect 115348 71408 115354 71420
rect 148226 71408 148232 71420
rect 148284 71448 148290 71460
rect 148686 71448 148692 71460
rect 148284 71420 148692 71448
rect 148284 71408 148290 71420
rect 148686 71408 148692 71420
rect 148744 71408 148750 71460
rect 160002 71408 160008 71460
rect 160060 71448 160066 71460
rect 193858 71448 193864 71460
rect 160060 71420 193864 71448
rect 160060 71408 160066 71420
rect 193858 71408 193864 71420
rect 193916 71408 193922 71460
rect 122190 71340 122196 71392
rect 122248 71380 122254 71392
rect 122248 71352 147674 71380
rect 122248 71340 122254 71352
rect 107654 71272 107660 71324
rect 107712 71312 107718 71324
rect 108022 71312 108028 71324
rect 107712 71284 108028 71312
rect 107712 71272 107718 71284
rect 108022 71272 108028 71284
rect 108080 71312 108086 71324
rect 140498 71312 140504 71324
rect 108080 71284 140504 71312
rect 108080 71272 108086 71284
rect 140498 71272 140504 71284
rect 140556 71272 140562 71324
rect 147646 71312 147674 71352
rect 170030 71340 170036 71392
rect 170088 71380 170094 71392
rect 170858 71380 170864 71392
rect 170088 71352 170864 71380
rect 170088 71340 170094 71352
rect 170858 71340 170864 71352
rect 170916 71340 170922 71392
rect 171778 71340 171784 71392
rect 171836 71380 171842 71392
rect 199562 71380 199568 71392
rect 171836 71352 199568 71380
rect 171836 71340 171842 71352
rect 199562 71340 199568 71352
rect 199620 71340 199626 71392
rect 153654 71312 153660 71324
rect 147646 71284 153660 71312
rect 153654 71272 153660 71284
rect 153712 71312 153718 71324
rect 154298 71312 154304 71324
rect 153712 71284 154304 71312
rect 153712 71272 153718 71284
rect 154298 71272 154304 71284
rect 154356 71272 154362 71324
rect 169570 71272 169576 71324
rect 169628 71312 169634 71324
rect 203518 71312 203524 71324
rect 169628 71284 203524 71312
rect 169628 71272 169634 71284
rect 203518 71272 203524 71284
rect 203576 71272 203582 71324
rect 111058 71204 111064 71256
rect 111116 71244 111122 71256
rect 142338 71244 142344 71256
rect 111116 71216 142344 71244
rect 111116 71204 111122 71216
rect 142338 71204 142344 71216
rect 142396 71204 142402 71256
rect 161014 71204 161020 71256
rect 161072 71244 161078 71256
rect 195606 71244 195612 71256
rect 161072 71216 195612 71244
rect 161072 71204 161078 71216
rect 195606 71204 195612 71216
rect 195664 71204 195670 71256
rect 118878 71136 118884 71188
rect 118936 71176 118942 71188
rect 150250 71176 150256 71188
rect 118936 71148 150256 71176
rect 118936 71136 118942 71148
rect 150250 71136 150256 71148
rect 150308 71136 150314 71188
rect 160922 71136 160928 71188
rect 160980 71176 160986 71188
rect 195514 71176 195520 71188
rect 160980 71148 195520 71176
rect 160980 71136 160986 71148
rect 195514 71136 195520 71148
rect 195572 71136 195578 71188
rect 71038 71068 71044 71120
rect 71096 71108 71102 71120
rect 107378 71108 107384 71120
rect 71096 71080 107384 71108
rect 71096 71068 71102 71080
rect 107378 71068 107384 71080
rect 107436 71108 107442 71120
rect 137646 71108 137652 71120
rect 107436 71080 137652 71108
rect 107436 71068 107442 71080
rect 137646 71068 137652 71080
rect 137704 71068 137710 71120
rect 147030 71068 147036 71120
rect 147088 71108 147094 71120
rect 184290 71108 184296 71120
rect 147088 71080 184296 71108
rect 147088 71068 147094 71080
rect 184290 71068 184296 71080
rect 184348 71068 184354 71120
rect 42794 71000 42800 71052
rect 42852 71040 42858 71052
rect 101490 71040 101496 71052
rect 42852 71012 101496 71040
rect 42852 71000 42858 71012
rect 101490 71000 101496 71012
rect 101548 71000 101554 71052
rect 104894 71000 104900 71052
rect 104952 71040 104958 71052
rect 132402 71040 132408 71052
rect 104952 71012 132408 71040
rect 104952 71000 104958 71012
rect 132402 71000 132408 71012
rect 132460 71000 132466 71052
rect 148962 71000 148968 71052
rect 149020 71040 149026 71052
rect 200114 71040 200120 71052
rect 149020 71012 200120 71040
rect 149020 71000 149026 71012
rect 200114 71000 200120 71012
rect 200172 71000 200178 71052
rect 212442 71000 212448 71052
rect 212500 71040 212506 71052
rect 480898 71040 480904 71052
rect 212500 71012 480904 71040
rect 212500 71000 212506 71012
rect 480898 71000 480904 71012
rect 480956 71000 480962 71052
rect 120350 70932 120356 70984
rect 120408 70972 120414 70984
rect 149238 70972 149244 70984
rect 120408 70944 149244 70972
rect 120408 70932 120414 70944
rect 149238 70932 149244 70944
rect 149296 70932 149302 70984
rect 170858 70932 170864 70984
rect 170916 70972 170922 70984
rect 204346 70972 204352 70984
rect 170916 70944 204352 70972
rect 170916 70932 170922 70944
rect 204346 70932 204352 70944
rect 204404 70932 204410 70984
rect 97442 70864 97448 70916
rect 97500 70904 97506 70916
rect 151170 70904 151176 70916
rect 97500 70876 151176 70904
rect 97500 70864 97506 70876
rect 151170 70864 151176 70876
rect 151228 70864 151234 70916
rect 158530 70864 158536 70916
rect 158588 70904 158594 70916
rect 191374 70904 191380 70916
rect 158588 70876 191380 70904
rect 158588 70864 158594 70876
rect 191374 70864 191380 70876
rect 191432 70864 191438 70916
rect 113542 70796 113548 70848
rect 113600 70836 113606 70848
rect 128446 70836 128452 70848
rect 113600 70808 128452 70836
rect 113600 70796 113606 70808
rect 128446 70796 128452 70808
rect 128504 70836 128510 70848
rect 129550 70836 129556 70848
rect 128504 70808 129556 70836
rect 128504 70796 128510 70808
rect 129550 70796 129556 70808
rect 129608 70796 129614 70848
rect 165522 70796 165528 70848
rect 165580 70836 165586 70848
rect 171778 70836 171784 70848
rect 165580 70808 171784 70836
rect 165580 70796 165586 70808
rect 171778 70796 171784 70808
rect 171836 70796 171842 70848
rect 178862 70796 178868 70848
rect 178920 70836 178926 70848
rect 219802 70836 219808 70848
rect 178920 70808 219808 70836
rect 178920 70796 178926 70808
rect 219802 70796 219808 70808
rect 219860 70796 219866 70848
rect 149238 70728 149244 70780
rect 149296 70768 149302 70780
rect 150066 70768 150072 70780
rect 149296 70740 150072 70768
rect 149296 70728 149302 70740
rect 150066 70728 150072 70740
rect 150124 70728 150130 70780
rect 97074 70320 97080 70372
rect 97132 70360 97138 70372
rect 151906 70360 151912 70372
rect 97132 70332 151912 70360
rect 97132 70320 97138 70332
rect 151906 70320 151912 70332
rect 151964 70320 151970 70372
rect 168098 70320 168104 70372
rect 168156 70360 168162 70372
rect 195054 70360 195060 70372
rect 168156 70332 195060 70360
rect 168156 70320 168162 70332
rect 195054 70320 195060 70332
rect 195112 70320 195118 70372
rect 151078 70292 151084 70304
rect 106246 70264 109034 70292
rect 97534 70184 97540 70236
rect 97592 70224 97598 70236
rect 106246 70224 106274 70264
rect 97592 70196 106274 70224
rect 109006 70224 109034 70264
rect 113146 70264 151084 70292
rect 113146 70224 113174 70264
rect 151078 70252 151084 70264
rect 151136 70252 151142 70304
rect 165246 70252 165252 70304
rect 165304 70292 165310 70304
rect 212994 70292 213000 70304
rect 165304 70264 213000 70292
rect 165304 70252 165310 70264
rect 212994 70252 213000 70264
rect 213052 70252 213058 70304
rect 109006 70196 113174 70224
rect 97592 70184 97598 70196
rect 115014 70184 115020 70236
rect 115072 70224 115078 70236
rect 150710 70224 150716 70236
rect 115072 70196 150716 70224
rect 115072 70184 115078 70196
rect 150710 70184 150716 70196
rect 150768 70184 150774 70236
rect 162394 70184 162400 70236
rect 162452 70224 162458 70236
rect 196434 70224 196440 70236
rect 162452 70196 196440 70224
rect 162452 70184 162458 70196
rect 196434 70184 196440 70196
rect 196492 70184 196498 70236
rect 98546 70116 98552 70168
rect 98604 70156 98610 70168
rect 132770 70156 132776 70168
rect 98604 70128 132776 70156
rect 98604 70116 98610 70128
rect 132770 70116 132776 70128
rect 132828 70116 132834 70168
rect 162302 70116 162308 70168
rect 162360 70156 162366 70168
rect 197078 70156 197084 70168
rect 162360 70128 197084 70156
rect 162360 70116 162366 70128
rect 197078 70116 197084 70128
rect 197136 70116 197142 70168
rect 108574 70048 108580 70100
rect 108632 70088 108638 70100
rect 142430 70088 142436 70100
rect 108632 70060 142436 70088
rect 108632 70048 108638 70060
rect 142430 70048 142436 70060
rect 142488 70048 142494 70100
rect 164602 70048 164608 70100
rect 164660 70088 164666 70100
rect 199746 70088 199752 70100
rect 164660 70060 199752 70088
rect 164660 70048 164666 70060
rect 199746 70048 199752 70060
rect 199804 70048 199810 70100
rect 108942 69980 108948 70032
rect 109000 70020 109006 70032
rect 142522 70020 142528 70032
rect 109000 69992 142528 70020
rect 109000 69980 109006 69992
rect 142522 69980 142528 69992
rect 142580 69980 142586 70032
rect 164786 69980 164792 70032
rect 164844 70020 164850 70032
rect 165246 70020 165252 70032
rect 164844 69992 165252 70020
rect 164844 69980 164850 69992
rect 165246 69980 165252 69992
rect 165304 69980 165310 70032
rect 199378 70020 199384 70032
rect 165448 69992 199384 70020
rect 165448 69964 165476 69992
rect 199378 69980 199384 69992
rect 199436 69980 199442 70032
rect 110966 69912 110972 69964
rect 111024 69952 111030 69964
rect 143994 69952 144000 69964
rect 111024 69924 144000 69952
rect 111024 69912 111030 69924
rect 143994 69912 144000 69924
rect 144052 69952 144058 69964
rect 146938 69952 146944 69964
rect 144052 69924 146944 69952
rect 144052 69912 144058 69924
rect 146938 69912 146944 69924
rect 146996 69912 147002 69964
rect 161566 69912 161572 69964
rect 161624 69952 161630 69964
rect 162302 69952 162308 69964
rect 161624 69924 162308 69952
rect 161624 69912 161630 69924
rect 162302 69912 162308 69924
rect 162360 69912 162366 69964
rect 164878 69912 164884 69964
rect 164936 69952 164942 69964
rect 165430 69952 165436 69964
rect 164936 69924 165436 69952
rect 164936 69912 164942 69924
rect 165430 69912 165436 69924
rect 165488 69912 165494 69964
rect 166166 69912 166172 69964
rect 166224 69952 166230 69964
rect 196986 69952 196992 69964
rect 166224 69924 196992 69952
rect 166224 69912 166230 69924
rect 196986 69912 196992 69924
rect 197044 69912 197050 69964
rect 101674 69844 101680 69896
rect 101732 69884 101738 69896
rect 101732 69856 109034 69884
rect 101732 69844 101738 69856
rect 85574 69776 85580 69828
rect 85632 69816 85638 69828
rect 105814 69816 105820 69828
rect 85632 69788 105820 69816
rect 85632 69776 85638 69788
rect 105814 69776 105820 69788
rect 105872 69776 105878 69828
rect 35986 69640 35992 69692
rect 36044 69680 36050 69692
rect 101674 69680 101680 69692
rect 36044 69652 101680 69680
rect 36044 69640 36050 69652
rect 101674 69640 101680 69652
rect 101732 69640 101738 69692
rect 105832 69680 105860 69776
rect 109006 69748 109034 69856
rect 110230 69844 110236 69896
rect 110288 69884 110294 69896
rect 142798 69884 142804 69896
rect 110288 69856 142804 69884
rect 110288 69844 110294 69856
rect 142798 69844 142804 69856
rect 142856 69844 142862 69896
rect 148410 69844 148416 69896
rect 148468 69884 148474 69896
rect 196618 69884 196624 69896
rect 148468 69856 196624 69884
rect 148468 69844 148474 69856
rect 196618 69844 196624 69856
rect 196676 69844 196682 69896
rect 118786 69776 118792 69828
rect 118844 69816 118850 69828
rect 152734 69816 152740 69828
rect 118844 69788 152740 69816
rect 118844 69776 118850 69788
rect 152734 69776 152740 69788
rect 152792 69776 152798 69828
rect 161658 69776 161664 69828
rect 161716 69816 161722 69828
rect 162394 69816 162400 69828
rect 161716 69788 162400 69816
rect 161716 69776 161722 69788
rect 162394 69776 162400 69788
rect 162452 69776 162458 69828
rect 162578 69776 162584 69828
rect 162636 69816 162642 69828
rect 189442 69816 189448 69828
rect 162636 69788 189448 69816
rect 162636 69776 162642 69788
rect 189442 69776 189448 69788
rect 189500 69816 189506 69828
rect 317414 69816 317420 69828
rect 189500 69788 317420 69816
rect 189500 69776 189506 69788
rect 317414 69776 317420 69788
rect 317472 69776 317478 69828
rect 134978 69748 134984 69760
rect 109006 69720 134984 69748
rect 134978 69708 134984 69720
rect 135036 69708 135042 69760
rect 159174 69708 159180 69760
rect 159232 69748 159238 69760
rect 193490 69748 193496 69760
rect 159232 69720 193496 69748
rect 159232 69708 159238 69720
rect 193490 69708 193496 69720
rect 193548 69748 193554 69760
rect 345014 69748 345020 69760
rect 193548 69720 345020 69748
rect 193548 69708 193554 69720
rect 345014 69708 345020 69720
rect 345072 69708 345078 69760
rect 138750 69680 138756 69692
rect 105832 69652 138756 69680
rect 138750 69640 138756 69652
rect 138808 69640 138814 69692
rect 147490 69640 147496 69692
rect 147548 69680 147554 69692
rect 182910 69680 182916 69692
rect 147548 69652 182916 69680
rect 147548 69640 147554 69652
rect 182910 69640 182916 69652
rect 182968 69640 182974 69692
rect 195054 69640 195060 69692
rect 195112 69680 195118 69692
rect 368474 69680 368480 69692
rect 195112 69652 368480 69680
rect 195112 69640 195118 69652
rect 368474 69640 368480 69652
rect 368532 69640 368538 69692
rect 111702 69572 111708 69624
rect 111760 69612 111766 69624
rect 142154 69612 142160 69624
rect 111760 69584 142160 69612
rect 111760 69572 111766 69584
rect 142154 69572 142160 69584
rect 142212 69612 142218 69624
rect 143074 69612 143080 69624
rect 142212 69584 143080 69612
rect 142212 69572 142218 69584
rect 143074 69572 143080 69584
rect 143132 69572 143138 69624
rect 161842 69572 161848 69624
rect 161900 69612 161906 69624
rect 162578 69612 162584 69624
rect 161900 69584 162584 69612
rect 161900 69572 161906 69584
rect 162578 69572 162584 69584
rect 162636 69572 162642 69624
rect 163498 69572 163504 69624
rect 163556 69612 163562 69624
rect 163958 69612 163964 69624
rect 163556 69584 163964 69612
rect 163556 69572 163562 69584
rect 163958 69572 163964 69584
rect 164016 69612 164022 69624
rect 164016 69584 171134 69612
rect 164016 69572 164022 69584
rect 102778 69504 102784 69556
rect 102836 69544 102842 69556
rect 132494 69544 132500 69556
rect 102836 69516 132500 69544
rect 102836 69504 102842 69516
rect 132494 69504 132500 69516
rect 132552 69504 132558 69556
rect 162596 69544 162624 69572
rect 166166 69544 166172 69556
rect 162596 69516 166172 69544
rect 166166 69504 166172 69516
rect 166224 69504 166230 69556
rect 171106 69544 171134 69584
rect 174262 69572 174268 69624
rect 174320 69612 174326 69624
rect 175090 69612 175096 69624
rect 174320 69584 175096 69612
rect 174320 69572 174326 69584
rect 175090 69572 175096 69584
rect 175148 69612 175154 69624
rect 208670 69612 208676 69624
rect 175148 69584 208676 69612
rect 175148 69572 175154 69584
rect 208670 69572 208676 69584
rect 208728 69572 208734 69624
rect 198366 69544 198372 69556
rect 171106 69516 198372 69544
rect 198366 69504 198372 69516
rect 198424 69504 198430 69556
rect 107194 69436 107200 69488
rect 107252 69476 107258 69488
rect 120074 69476 120080 69488
rect 107252 69448 120080 69476
rect 107252 69436 107258 69448
rect 120074 69436 120080 69448
rect 120132 69436 120138 69488
rect 161750 69436 161756 69488
rect 161808 69476 161814 69488
rect 162762 69476 162768 69488
rect 161808 69448 162768 69476
rect 161808 69436 161814 69448
rect 162762 69436 162768 69448
rect 162820 69476 162826 69488
rect 210418 69476 210424 69488
rect 162820 69448 210424 69476
rect 162820 69436 162826 69448
rect 210418 69436 210424 69448
rect 210476 69436 210482 69488
rect 120166 69368 120172 69420
rect 120224 69408 120230 69420
rect 120718 69408 120724 69420
rect 120224 69380 120724 69408
rect 120224 69368 120230 69380
rect 120718 69368 120724 69380
rect 120776 69408 120782 69420
rect 120776 69380 122834 69408
rect 120776 69368 120782 69380
rect 122806 69340 122834 69380
rect 141234 69340 141240 69352
rect 122806 69312 141240 69340
rect 141234 69300 141240 69312
rect 141292 69300 141298 69352
rect 102778 69028 102784 69080
rect 102836 69068 102842 69080
rect 105538 69068 105544 69080
rect 102836 69040 105544 69068
rect 102836 69028 102842 69040
rect 105538 69028 105544 69040
rect 105596 69028 105602 69080
rect 150710 69028 150716 69080
rect 150768 69068 150774 69080
rect 151538 69068 151544 69080
rect 150768 69040 151544 69068
rect 150768 69028 150774 69040
rect 151538 69028 151544 69040
rect 151596 69028 151602 69080
rect 99282 68960 99288 69012
rect 99340 69000 99346 69012
rect 153470 69000 153476 69012
rect 99340 68972 153476 69000
rect 99340 68960 99346 68972
rect 153470 68960 153476 68972
rect 153528 68960 153534 69012
rect 160370 68960 160376 69012
rect 160428 69000 160434 69012
rect 214558 69000 214564 69012
rect 160428 68972 214564 69000
rect 160428 68960 160434 68972
rect 214558 68960 214564 68972
rect 214616 68960 214622 69012
rect 114094 68892 114100 68944
rect 114152 68932 114158 68944
rect 114152 68904 145052 68932
rect 114152 68892 114158 68904
rect 115474 68824 115480 68876
rect 115532 68864 115538 68876
rect 145024 68864 145052 68904
rect 145098 68892 145104 68944
rect 145156 68932 145162 68944
rect 147030 68932 147036 68944
rect 145156 68904 147036 68932
rect 145156 68892 145162 68904
rect 147030 68892 147036 68904
rect 147088 68892 147094 68944
rect 166074 68892 166080 68944
rect 166132 68932 166138 68944
rect 166810 68932 166816 68944
rect 166132 68904 166816 68932
rect 166132 68892 166138 68904
rect 166810 68892 166816 68904
rect 166868 68892 166874 68944
rect 211890 68932 211896 68944
rect 171106 68904 211896 68932
rect 148594 68864 148600 68876
rect 115532 68836 142154 68864
rect 145024 68836 148600 68864
rect 115532 68824 115538 68836
rect 102962 68796 102968 68808
rect 99346 68768 102968 68796
rect 60734 68620 60740 68672
rect 60792 68660 60798 68672
rect 99346 68660 99374 68768
rect 102962 68756 102968 68768
rect 103020 68796 103026 68808
rect 137094 68796 137100 68808
rect 103020 68768 137100 68796
rect 103020 68756 103026 68768
rect 137094 68756 137100 68768
rect 137152 68756 137158 68808
rect 142126 68796 142154 68836
rect 148594 68824 148600 68836
rect 148652 68864 148658 68876
rect 148870 68864 148876 68876
rect 148652 68836 148876 68864
rect 148652 68824 148658 68836
rect 148870 68824 148876 68836
rect 148928 68824 148934 68876
rect 165982 68824 165988 68876
rect 166040 68864 166046 68876
rect 171106 68864 171134 68904
rect 211890 68892 211896 68904
rect 211948 68892 211954 68944
rect 166040 68836 171134 68864
rect 166040 68824 166046 68836
rect 171502 68824 171508 68876
rect 171560 68864 171566 68876
rect 172146 68864 172152 68876
rect 171560 68836 172152 68864
rect 171560 68824 171566 68836
rect 172146 68824 172152 68836
rect 172204 68824 172210 68876
rect 172882 68824 172888 68876
rect 172940 68864 172946 68876
rect 173710 68864 173716 68876
rect 172940 68836 173716 68864
rect 172940 68824 172946 68836
rect 173710 68824 173716 68836
rect 173768 68824 173774 68876
rect 177666 68824 177672 68876
rect 177724 68864 177730 68876
rect 209958 68864 209964 68876
rect 177724 68836 209964 68864
rect 177724 68824 177730 68836
rect 209958 68824 209964 68836
rect 210016 68864 210022 68876
rect 211062 68864 211068 68876
rect 210016 68836 211068 68864
rect 210016 68824 210022 68836
rect 211062 68824 211068 68836
rect 211120 68824 211126 68876
rect 149514 68796 149520 68808
rect 142126 68768 149520 68796
rect 149514 68756 149520 68768
rect 149572 68756 149578 68808
rect 165798 68756 165804 68808
rect 165856 68796 165862 68808
rect 166442 68796 166448 68808
rect 165856 68768 166448 68796
rect 165856 68756 165862 68768
rect 166442 68756 166448 68768
rect 166500 68756 166506 68808
rect 171410 68756 171416 68808
rect 171468 68796 171474 68808
rect 172330 68796 172336 68808
rect 171468 68768 172336 68796
rect 171468 68756 171474 68768
rect 172330 68756 172336 68768
rect 172388 68756 172394 68808
rect 175918 68756 175924 68808
rect 175976 68796 175982 68808
rect 200666 68796 200672 68808
rect 175976 68768 200672 68796
rect 175976 68756 175982 68768
rect 200666 68756 200672 68768
rect 200724 68756 200730 68808
rect 108758 68688 108764 68740
rect 108816 68728 108822 68740
rect 142706 68728 142712 68740
rect 108816 68700 142712 68728
rect 108816 68688 108822 68700
rect 142706 68688 142712 68700
rect 142764 68728 142770 68740
rect 142890 68728 142896 68740
rect 142764 68700 142896 68728
rect 142764 68688 142770 68700
rect 142890 68688 142896 68700
rect 142948 68688 142954 68740
rect 165706 68688 165712 68740
rect 165764 68728 165770 68740
rect 166350 68728 166356 68740
rect 165764 68700 166356 68728
rect 165764 68688 165770 68700
rect 166350 68688 166356 68700
rect 166408 68688 166414 68740
rect 168834 68688 168840 68740
rect 168892 68728 168898 68740
rect 169386 68728 169392 68740
rect 168892 68700 169392 68728
rect 168892 68688 168898 68700
rect 169386 68688 169392 68700
rect 169444 68728 169450 68740
rect 203426 68728 203432 68740
rect 169444 68700 203432 68728
rect 169444 68688 169450 68700
rect 203426 68688 203432 68700
rect 203484 68688 203490 68740
rect 60792 68632 99374 68660
rect 60792 68620 60798 68632
rect 103330 68620 103336 68672
rect 103388 68660 103394 68672
rect 135622 68660 135628 68672
rect 103388 68632 135628 68660
rect 103388 68620 103394 68632
rect 135622 68620 135628 68632
rect 135680 68620 135686 68672
rect 166810 68620 166816 68672
rect 166868 68660 166874 68672
rect 201218 68660 201224 68672
rect 166868 68632 201224 68660
rect 166868 68620 166874 68632
rect 201218 68620 201224 68632
rect 201276 68620 201282 68672
rect 34514 68552 34520 68604
rect 34572 68592 34578 68604
rect 99834 68592 99840 68604
rect 34572 68564 99840 68592
rect 34572 68552 34578 68564
rect 99834 68552 99840 68564
rect 99892 68552 99898 68604
rect 112898 68552 112904 68604
rect 112956 68592 112962 68604
rect 112956 68564 137324 68592
rect 112956 68552 112962 68564
rect 99190 68484 99196 68536
rect 99248 68524 99254 68536
rect 131574 68524 131580 68536
rect 99248 68496 131580 68524
rect 99248 68484 99254 68496
rect 131574 68484 131580 68496
rect 131632 68524 131638 68536
rect 132678 68524 132684 68536
rect 131632 68496 132684 68524
rect 131632 68484 131638 68496
rect 132678 68484 132684 68496
rect 132736 68484 132742 68536
rect 137296 68524 137324 68564
rect 140038 68552 140044 68604
rect 140096 68592 140102 68604
rect 142246 68592 142252 68604
rect 140096 68564 142252 68592
rect 140096 68552 140102 68564
rect 142246 68552 142252 68564
rect 142304 68552 142310 68604
rect 149146 68552 149152 68604
rect 149204 68592 149210 68604
rect 220814 68592 220820 68604
rect 149204 68564 220820 68592
rect 149204 68552 149210 68564
rect 220814 68552 220820 68564
rect 220872 68552 220878 68604
rect 144362 68524 144368 68536
rect 137296 68496 144368 68524
rect 144362 68484 144368 68496
rect 144420 68484 144426 68536
rect 172330 68484 172336 68536
rect 172388 68524 172394 68536
rect 205818 68524 205824 68536
rect 172388 68496 205824 68524
rect 172388 68484 172394 68496
rect 205818 68484 205824 68496
rect 205876 68484 205882 68536
rect 214558 68484 214564 68536
rect 214616 68524 214622 68536
rect 358814 68524 358820 68536
rect 214616 68496 358820 68524
rect 214616 68484 214622 68496
rect 358814 68484 358820 68496
rect 358872 68484 358878 68536
rect 103146 68416 103152 68468
rect 103204 68456 103210 68468
rect 134242 68456 134248 68468
rect 103204 68428 134248 68456
rect 103204 68416 103210 68428
rect 134242 68416 134248 68428
rect 134300 68416 134306 68468
rect 165338 68416 165344 68468
rect 165396 68456 165402 68468
rect 197814 68456 197820 68468
rect 165396 68428 197820 68456
rect 165396 68416 165402 68428
rect 197814 68416 197820 68428
rect 197872 68456 197878 68468
rect 396074 68456 396080 68468
rect 197872 68428 396080 68456
rect 197872 68416 197878 68428
rect 396074 68416 396080 68428
rect 396132 68416 396138 68468
rect 40034 68348 40040 68400
rect 40092 68388 40098 68400
rect 103330 68388 103336 68400
rect 40092 68360 103336 68388
rect 40092 68348 40098 68360
rect 103330 68348 103336 68360
rect 103388 68348 103394 68400
rect 110782 68348 110788 68400
rect 110840 68388 110846 68400
rect 142706 68388 142712 68400
rect 110840 68360 142712 68388
rect 110840 68348 110846 68360
rect 142706 68348 142712 68360
rect 142764 68388 142770 68400
rect 142982 68388 142988 68400
rect 142764 68360 142988 68388
rect 142764 68348 142770 68360
rect 142982 68348 142988 68360
rect 143040 68348 143046 68400
rect 165890 68348 165896 68400
rect 165948 68388 165954 68400
rect 193766 68388 193772 68400
rect 165948 68360 193772 68388
rect 165948 68348 165954 68360
rect 193766 68348 193772 68360
rect 193824 68388 193830 68400
rect 440234 68388 440240 68400
rect 193824 68360 440240 68388
rect 193824 68348 193830 68360
rect 440234 68348 440240 68360
rect 440292 68348 440298 68400
rect 97166 68280 97172 68332
rect 97224 68320 97230 68332
rect 106274 68320 106280 68332
rect 97224 68292 106280 68320
rect 97224 68280 97230 68292
rect 106274 68280 106280 68292
rect 106332 68320 106338 68332
rect 139670 68320 139676 68332
rect 106332 68292 139676 68320
rect 106332 68280 106338 68292
rect 139670 68280 139676 68292
rect 139728 68280 139734 68332
rect 147306 68280 147312 68332
rect 147364 68320 147370 68332
rect 189718 68320 189724 68332
rect 147364 68292 189724 68320
rect 147364 68280 147370 68292
rect 189718 68280 189724 68292
rect 189776 68280 189782 68332
rect 211062 68280 211068 68332
rect 211120 68320 211126 68332
rect 536834 68320 536840 68332
rect 211120 68292 536840 68320
rect 211120 68280 211126 68292
rect 536834 68280 536840 68292
rect 536892 68280 536898 68332
rect 118970 68212 118976 68264
rect 119028 68252 119034 68264
rect 141970 68252 141976 68264
rect 119028 68224 141976 68252
rect 119028 68212 119034 68224
rect 141970 68212 141976 68224
rect 142028 68212 142034 68264
rect 173710 68212 173716 68264
rect 173768 68252 173774 68264
rect 207198 68252 207204 68264
rect 173768 68224 207204 68252
rect 173768 68212 173774 68224
rect 207198 68212 207204 68224
rect 207256 68212 207262 68264
rect 172146 68144 172152 68196
rect 172204 68184 172210 68196
rect 205634 68184 205640 68196
rect 172204 68156 205640 68184
rect 172204 68144 172210 68156
rect 205634 68144 205640 68156
rect 205692 68144 205698 68196
rect 166442 68076 166448 68128
rect 166500 68116 166506 68128
rect 175918 68116 175924 68128
rect 166500 68088 175924 68116
rect 166500 68076 166506 68088
rect 175918 68076 175924 68088
rect 175976 68076 175982 68128
rect 200850 68116 200856 68128
rect 180766 68088 200856 68116
rect 166350 68008 166356 68060
rect 166408 68048 166414 68060
rect 180766 68048 180794 68088
rect 200850 68076 200856 68088
rect 200908 68076 200914 68128
rect 166408 68020 180794 68048
rect 166408 68008 166414 68020
rect 149514 67600 149520 67652
rect 149572 67640 149578 67652
rect 149882 67640 149888 67652
rect 149572 67612 149888 67640
rect 149572 67600 149578 67612
rect 149882 67600 149888 67612
rect 149940 67600 149946 67652
rect 153470 67600 153476 67652
rect 153528 67640 153534 67652
rect 154206 67640 154212 67652
rect 153528 67612 154212 67640
rect 153528 67600 153534 67612
rect 154206 67600 154212 67612
rect 154264 67600 154270 67652
rect 166092 67612 166304 67640
rect 124858 67532 124864 67584
rect 124916 67572 124922 67584
rect 135346 67572 135352 67584
rect 124916 67544 135352 67572
rect 124916 67532 124922 67544
rect 135346 67532 135352 67544
rect 135404 67572 135410 67584
rect 135898 67572 135904 67584
rect 135404 67544 135904 67572
rect 135404 67532 135410 67544
rect 135898 67532 135904 67544
rect 135956 67532 135962 67584
rect 145650 67572 145656 67584
rect 142126 67544 145656 67572
rect 96982 67464 96988 67516
rect 97040 67504 97046 67516
rect 142126 67504 142154 67544
rect 145650 67532 145656 67544
rect 145708 67572 145714 67584
rect 146018 67572 146024 67584
rect 145708 67544 146024 67572
rect 145708 67532 145714 67544
rect 146018 67532 146024 67544
rect 146076 67532 146082 67584
rect 163406 67532 163412 67584
rect 163464 67572 163470 67584
rect 164142 67572 164148 67584
rect 163464 67544 164148 67572
rect 163464 67532 163470 67544
rect 164142 67532 164148 67544
rect 164200 67532 164206 67584
rect 164510 67532 164516 67584
rect 164568 67572 164574 67584
rect 165154 67572 165160 67584
rect 164568 67544 165160 67572
rect 164568 67532 164574 67544
rect 165154 67532 165160 67544
rect 165212 67532 165218 67584
rect 97040 67476 142154 67504
rect 164160 67504 164188 67532
rect 166092 67504 166120 67612
rect 166276 67572 166304 67612
rect 211614 67572 211620 67584
rect 166276 67544 211620 67572
rect 211614 67532 211620 67544
rect 211672 67532 211678 67584
rect 164160 67476 166120 67504
rect 97040 67464 97046 67476
rect 166166 67464 166172 67516
rect 166224 67504 166230 67516
rect 212718 67504 212724 67516
rect 166224 67476 212724 67504
rect 166224 67464 166230 67476
rect 212718 67464 212724 67476
rect 212776 67464 212782 67516
rect 119798 67396 119804 67448
rect 119856 67436 119862 67448
rect 153286 67436 153292 67448
rect 119856 67408 153292 67436
rect 119856 67396 119862 67408
rect 153286 67396 153292 67408
rect 153344 67396 153350 67448
rect 157702 67396 157708 67448
rect 157760 67436 157766 67448
rect 192570 67436 192576 67448
rect 157760 67408 192576 67436
rect 157760 67396 157766 67408
rect 192570 67396 192576 67408
rect 192628 67436 192634 67448
rect 193030 67436 193036 67448
rect 192628 67408 193036 67436
rect 192628 67396 192634 67408
rect 193030 67396 193036 67408
rect 193088 67396 193094 67448
rect 100018 67328 100024 67380
rect 100076 67368 100082 67380
rect 133966 67368 133972 67380
rect 100076 67340 133972 67368
rect 100076 67328 100082 67340
rect 133966 67328 133972 67340
rect 134024 67368 134030 67380
rect 134518 67368 134524 67380
rect 134024 67340 134524 67368
rect 134024 67328 134030 67340
rect 134518 67328 134524 67340
rect 134576 67328 134582 67380
rect 165154 67328 165160 67380
rect 165212 67368 165218 67380
rect 199654 67368 199660 67380
rect 165212 67340 199660 67368
rect 165212 67328 165218 67340
rect 199654 67328 199660 67340
rect 199712 67328 199718 67380
rect 100110 67260 100116 67312
rect 100168 67300 100174 67312
rect 134058 67300 134064 67312
rect 100168 67272 134064 67300
rect 100168 67260 100174 67272
rect 134058 67260 134064 67272
rect 134116 67300 134122 67312
rect 134610 67300 134616 67312
rect 134116 67272 134616 67300
rect 134116 67260 134122 67272
rect 134610 67260 134616 67272
rect 134668 67260 134674 67312
rect 165614 67260 165620 67312
rect 165672 67300 165678 67312
rect 166166 67300 166172 67312
rect 165672 67272 166172 67300
rect 165672 67260 165678 67272
rect 166166 67260 166172 67272
rect 166224 67260 166230 67312
rect 177022 67260 177028 67312
rect 177080 67300 177086 67312
rect 177850 67300 177856 67312
rect 177080 67272 177856 67300
rect 177080 67260 177086 67272
rect 177850 67260 177856 67272
rect 177908 67300 177914 67312
rect 211338 67300 211344 67312
rect 177908 67272 211344 67300
rect 177908 67260 177914 67272
rect 211338 67260 211344 67272
rect 211396 67260 211402 67312
rect 100386 67192 100392 67244
rect 100444 67232 100450 67244
rect 134150 67232 134156 67244
rect 100444 67204 134156 67232
rect 100444 67192 100450 67204
rect 134150 67192 134156 67204
rect 134208 67192 134214 67244
rect 166718 67192 166724 67244
rect 166776 67232 166782 67244
rect 196158 67232 196164 67244
rect 166776 67204 196164 67232
rect 166776 67192 166782 67204
rect 196158 67192 196164 67204
rect 196216 67192 196222 67244
rect 104434 67124 104440 67176
rect 104492 67164 104498 67176
rect 138842 67164 138848 67176
rect 104492 67136 138848 67164
rect 104492 67124 104498 67136
rect 138842 67124 138848 67136
rect 138900 67124 138906 67176
rect 175458 67124 175464 67176
rect 175516 67164 175522 67176
rect 204898 67164 204904 67176
rect 175516 67136 204904 67164
rect 175516 67124 175522 67136
rect 204898 67124 204904 67136
rect 204956 67124 204962 67176
rect 136174 67096 136180 67108
rect 104544 67068 136180 67096
rect 77294 66920 77300 66972
rect 77352 66960 77358 66972
rect 104434 66960 104440 66972
rect 77352 66932 104440 66960
rect 77352 66920 77358 66932
rect 104434 66920 104440 66932
rect 104492 66920 104498 66972
rect 44174 66852 44180 66904
rect 44232 66892 44238 66904
rect 101766 66892 101772 66904
rect 44232 66864 101772 66892
rect 44232 66852 44238 66864
rect 101766 66852 101772 66864
rect 101824 66892 101830 66904
rect 104544 66892 104572 67068
rect 136174 67056 136180 67068
rect 136232 67056 136238 67108
rect 147950 67056 147956 67108
rect 148008 67096 148014 67108
rect 203518 67096 203524 67108
rect 148008 67068 203524 67096
rect 148008 67056 148014 67068
rect 203518 67056 203524 67068
rect 203576 67056 203582 67108
rect 106918 66988 106924 67040
rect 106976 67028 106982 67040
rect 109402 67028 109408 67040
rect 106976 67000 109408 67028
rect 106976 66988 106982 67000
rect 109402 66988 109408 67000
rect 109460 67028 109466 67040
rect 140130 67028 140136 67040
rect 109460 67000 140136 67028
rect 109460 66988 109466 67000
rect 140130 66988 140136 67000
rect 140188 66988 140194 67040
rect 154298 66988 154304 67040
rect 154356 67028 154362 67040
rect 274634 67028 274640 67040
rect 154356 67000 274640 67028
rect 154356 66988 154362 67000
rect 274634 66988 274640 67000
rect 274692 66988 274698 67040
rect 107562 66920 107568 66972
rect 107620 66960 107626 66972
rect 135530 66960 135536 66972
rect 107620 66932 135536 66960
rect 107620 66920 107626 66932
rect 135530 66920 135536 66932
rect 135588 66920 135594 66972
rect 159082 66920 159088 66972
rect 159140 66960 159146 66972
rect 159726 66960 159732 66972
rect 159140 66932 159732 66960
rect 159140 66920 159146 66932
rect 159726 66920 159732 66932
rect 159784 66960 159790 66972
rect 188338 66960 188344 66972
rect 159784 66932 188344 66960
rect 159784 66920 159790 66932
rect 188338 66920 188344 66932
rect 188396 66920 188402 66972
rect 193030 66920 193036 66972
rect 193088 66960 193094 66972
rect 332686 66960 332692 66972
rect 193088 66932 332692 66960
rect 193088 66920 193094 66932
rect 332686 66920 332692 66932
rect 332744 66920 332750 66972
rect 101824 66864 104572 66892
rect 101824 66852 101830 66864
rect 120074 66852 120080 66904
rect 120132 66892 120138 66904
rect 120718 66892 120724 66904
rect 120132 66864 120724 66892
rect 120132 66852 120138 66864
rect 120718 66852 120724 66864
rect 120776 66892 120782 66904
rect 141142 66892 141148 66904
rect 120776 66864 141148 66892
rect 120776 66852 120782 66864
rect 141142 66852 141148 66864
rect 141200 66852 141206 66904
rect 165982 66852 165988 66904
rect 166040 66892 166046 66904
rect 166810 66892 166816 66904
rect 166040 66864 166816 66892
rect 166040 66852 166046 66864
rect 166810 66852 166816 66864
rect 166868 66852 166874 66904
rect 188430 66892 188436 66904
rect 171106 66864 188436 66892
rect 120258 66784 120264 66836
rect 120316 66824 120322 66836
rect 120810 66824 120816 66836
rect 120316 66796 120816 66824
rect 120316 66784 120322 66796
rect 120810 66784 120816 66796
rect 120868 66824 120874 66836
rect 141050 66824 141056 66836
rect 120868 66796 141056 66824
rect 120868 66784 120874 66796
rect 141050 66784 141056 66796
rect 141108 66784 141114 66836
rect 162118 66784 162124 66836
rect 162176 66824 162182 66836
rect 171106 66824 171134 66864
rect 188430 66852 188436 66864
rect 188488 66852 188494 66904
rect 196158 66852 196164 66904
rect 196216 66892 196222 66904
rect 196894 66892 196900 66904
rect 196216 66864 196900 66892
rect 196216 66852 196222 66864
rect 196894 66852 196900 66864
rect 196952 66892 196958 66904
rect 375374 66892 375380 66904
rect 196952 66864 375380 66892
rect 196952 66852 196958 66864
rect 375374 66852 375380 66864
rect 375432 66852 375438 66904
rect 162176 66796 171134 66824
rect 162176 66784 162182 66796
rect 97718 66716 97724 66768
rect 97776 66756 97782 66768
rect 151262 66756 151268 66768
rect 97776 66728 151268 66756
rect 97776 66716 97782 66728
rect 151262 66716 151268 66728
rect 151320 66716 151326 66768
rect 153286 66240 153292 66292
rect 153344 66280 153350 66292
rect 154022 66280 154028 66292
rect 153344 66252 154028 66280
rect 153344 66240 153350 66252
rect 154022 66240 154028 66252
rect 154080 66240 154086 66292
rect 176856 66252 177804 66280
rect 110046 66172 110052 66224
rect 110104 66212 110110 66224
rect 143902 66212 143908 66224
rect 110104 66184 143908 66212
rect 110104 66172 110110 66184
rect 143902 66172 143908 66184
rect 143960 66212 143966 66224
rect 147122 66212 147128 66224
rect 143960 66184 147128 66212
rect 143960 66172 143966 66184
rect 147122 66172 147128 66184
rect 147180 66172 147186 66224
rect 163314 66172 163320 66224
rect 163372 66212 163378 66224
rect 164050 66212 164056 66224
rect 163372 66184 164056 66212
rect 163372 66172 163378 66184
rect 164050 66172 164056 66184
rect 164108 66172 164114 66224
rect 172790 66172 172796 66224
rect 172848 66212 172854 66224
rect 173618 66212 173624 66224
rect 172848 66184 173624 66212
rect 172848 66172 172854 66184
rect 173618 66172 173624 66184
rect 173676 66172 173682 66224
rect 175366 66172 175372 66224
rect 175424 66212 175430 66224
rect 176286 66212 176292 66224
rect 175424 66184 176292 66212
rect 175424 66172 175430 66184
rect 176286 66172 176292 66184
rect 176344 66212 176350 66224
rect 176856 66212 176884 66252
rect 176344 66184 176884 66212
rect 176344 66172 176350 66184
rect 176930 66172 176936 66224
rect 176988 66212 176994 66224
rect 177666 66212 177672 66224
rect 176988 66184 177672 66212
rect 176988 66172 176994 66184
rect 177666 66172 177672 66184
rect 177724 66172 177730 66224
rect 177776 66212 177804 66252
rect 204898 66240 204904 66292
rect 204956 66280 204962 66292
rect 554038 66280 554044 66292
rect 204956 66252 554044 66280
rect 204956 66240 204962 66252
rect 554038 66240 554044 66252
rect 554096 66240 554102 66292
rect 210234 66212 210240 66224
rect 177776 66184 210240 66212
rect 210234 66172 210240 66184
rect 210292 66172 210298 66224
rect 104434 66104 104440 66156
rect 104492 66144 104498 66156
rect 136910 66144 136916 66156
rect 104492 66116 136916 66144
rect 104492 66104 104498 66116
rect 136910 66104 136916 66116
rect 136968 66104 136974 66156
rect 177684 66144 177712 66172
rect 211706 66144 211712 66156
rect 177684 66116 211712 66144
rect 211706 66104 211712 66116
rect 211764 66104 211770 66156
rect 103238 66036 103244 66088
rect 103296 66076 103302 66088
rect 103422 66076 103428 66088
rect 103296 66048 103428 66076
rect 103296 66036 103302 66048
rect 103422 66036 103428 66048
rect 103480 66076 103486 66088
rect 135806 66076 135812 66088
rect 103480 66048 135812 66076
rect 103480 66036 103486 66048
rect 135806 66036 135812 66048
rect 135864 66036 135870 66088
rect 164418 66036 164424 66088
rect 164476 66076 164482 66088
rect 198918 66076 198924 66088
rect 164476 66048 198924 66076
rect 164476 66036 164482 66048
rect 198918 66036 198924 66048
rect 198976 66036 198982 66088
rect 139854 66008 139860 66020
rect 109006 65980 139860 66008
rect 93118 65900 93124 65952
rect 93176 65940 93182 65952
rect 107010 65940 107016 65952
rect 93176 65912 107016 65940
rect 93176 65900 93182 65912
rect 107010 65900 107016 65912
rect 107068 65940 107074 65952
rect 109006 65940 109034 65980
rect 139854 65968 139860 65980
rect 139912 65968 139918 66020
rect 173618 65968 173624 66020
rect 173676 66008 173682 66020
rect 205726 66008 205732 66020
rect 173676 65980 205732 66008
rect 173676 65968 173682 65980
rect 205726 65968 205732 65980
rect 205784 65968 205790 66020
rect 107068 65912 109034 65940
rect 107068 65900 107074 65912
rect 110322 65900 110328 65952
rect 110380 65940 110386 65952
rect 142154 65940 142160 65952
rect 110380 65912 142160 65940
rect 110380 65900 110386 65912
rect 142154 65900 142160 65912
rect 142212 65940 142218 65952
rect 142614 65940 142620 65952
rect 142212 65912 142620 65940
rect 142212 65900 142218 65912
rect 142614 65900 142620 65912
rect 142672 65900 142678 65952
rect 154942 65900 154948 65952
rect 155000 65940 155006 65952
rect 155678 65940 155684 65952
rect 155000 65912 155684 65940
rect 155000 65900 155006 65912
rect 155678 65900 155684 65912
rect 155736 65940 155742 65952
rect 186958 65940 186964 65952
rect 155736 65912 186964 65940
rect 155736 65900 155742 65912
rect 186958 65900 186964 65912
rect 187016 65900 187022 65952
rect 134426 65872 134432 65884
rect 109006 65844 134432 65872
rect 78674 65764 78680 65816
rect 78732 65804 78738 65816
rect 104710 65804 104716 65816
rect 78732 65776 104716 65804
rect 78732 65764 78738 65776
rect 104710 65764 104716 65776
rect 104768 65764 104774 65816
rect 75914 65696 75920 65748
rect 75972 65736 75978 65748
rect 104158 65736 104164 65748
rect 75972 65708 104164 65736
rect 75972 65696 75978 65708
rect 104158 65696 104164 65708
rect 104216 65696 104222 65748
rect 60826 65628 60832 65680
rect 60884 65668 60890 65680
rect 105722 65668 105728 65680
rect 60884 65640 105728 65668
rect 60884 65628 60890 65640
rect 105722 65628 105728 65640
rect 105780 65628 105786 65680
rect 52546 65560 52552 65612
rect 52604 65600 52610 65612
rect 103422 65600 103428 65612
rect 52604 65572 103428 65600
rect 52604 65560 52610 65572
rect 103422 65560 103428 65572
rect 103480 65560 103486 65612
rect 35158 65492 35164 65544
rect 35216 65532 35222 65544
rect 103330 65532 103336 65544
rect 35216 65504 103336 65532
rect 35216 65492 35222 65504
rect 103330 65492 103336 65504
rect 103388 65532 103394 65544
rect 109006 65532 109034 65844
rect 134426 65832 134432 65844
rect 134484 65832 134490 65884
rect 164050 65832 164056 65884
rect 164108 65872 164114 65884
rect 191282 65872 191288 65884
rect 164108 65844 191288 65872
rect 164108 65832 164114 65844
rect 191282 65832 191288 65844
rect 191340 65832 191346 65884
rect 113174 65764 113180 65816
rect 113232 65804 113238 65816
rect 120258 65804 120264 65816
rect 113232 65776 120264 65804
rect 113232 65764 113238 65776
rect 120258 65764 120264 65776
rect 120316 65764 120322 65816
rect 160278 65764 160284 65816
rect 160336 65804 160342 65816
rect 161014 65804 161020 65816
rect 160336 65776 161020 65804
rect 160336 65764 160342 65776
rect 161014 65764 161020 65776
rect 161072 65804 161078 65816
rect 187050 65804 187056 65816
rect 161072 65776 187056 65804
rect 161072 65764 161078 65776
rect 187050 65764 187056 65776
rect 187108 65764 187114 65816
rect 147858 65560 147864 65612
rect 147916 65600 147922 65612
rect 209958 65600 209964 65612
rect 147916 65572 209964 65600
rect 147916 65560 147922 65572
rect 209958 65560 209964 65572
rect 210016 65560 210022 65612
rect 103388 65504 109034 65532
rect 103388 65492 103394 65504
rect 198918 65492 198924 65544
rect 198976 65532 198982 65544
rect 418798 65532 418804 65544
rect 198976 65504 418804 65532
rect 198976 65492 198982 65504
rect 418798 65492 418804 65504
rect 418856 65492 418862 65544
rect 141510 64880 141516 64932
rect 141568 64920 141574 64932
rect 142246 64920 142252 64932
rect 141568 64892 142252 64920
rect 141568 64880 141574 64892
rect 142246 64880 142252 64892
rect 142304 64880 142310 64932
rect 97810 64812 97816 64864
rect 97868 64852 97874 64864
rect 144086 64852 144092 64864
rect 97868 64824 144092 64852
rect 97868 64812 97874 64824
rect 144086 64812 144092 64824
rect 144144 64812 144150 64864
rect 174170 64812 174176 64864
rect 174228 64852 174234 64864
rect 214374 64852 214380 64864
rect 174228 64824 214380 64852
rect 174228 64812 174234 64824
rect 214374 64812 214380 64824
rect 214432 64812 214438 64864
rect 104158 64744 104164 64796
rect 104216 64784 104222 64796
rect 138474 64784 138480 64796
rect 104216 64756 138480 64784
rect 104216 64744 104222 64756
rect 138474 64744 138480 64756
rect 138532 64744 138538 64796
rect 158990 64744 158996 64796
rect 159048 64784 159054 64796
rect 193398 64784 193404 64796
rect 159048 64756 193404 64784
rect 159048 64744 159054 64756
rect 193398 64744 193404 64756
rect 193456 64744 193462 64796
rect 103790 64676 103796 64728
rect 103848 64716 103854 64728
rect 137462 64716 137468 64728
rect 103848 64688 137468 64716
rect 103848 64676 103854 64688
rect 137462 64676 137468 64688
rect 137520 64676 137526 64728
rect 168650 64676 168656 64728
rect 168708 64716 168714 64728
rect 203058 64716 203064 64728
rect 168708 64688 203064 64716
rect 168708 64676 168714 64688
rect 203058 64676 203064 64688
rect 203116 64676 203122 64728
rect 103974 64608 103980 64660
rect 104032 64648 104038 64660
rect 132586 64648 132592 64660
rect 104032 64620 132592 64648
rect 104032 64608 104038 64620
rect 132586 64608 132592 64620
rect 132644 64608 132650 64660
rect 149790 64404 149796 64456
rect 149848 64444 149854 64456
rect 224954 64444 224960 64456
rect 149848 64416 224960 64444
rect 149848 64404 149854 64416
rect 224954 64404 224960 64416
rect 225012 64404 225018 64456
rect 152642 64336 152648 64388
rect 152700 64376 152706 64388
rect 256694 64376 256700 64388
rect 152700 64348 256700 64376
rect 152700 64336 152706 64348
rect 256694 64336 256700 64348
rect 256752 64336 256758 64388
rect 193398 64268 193404 64320
rect 193456 64308 193462 64320
rect 340966 64308 340972 64320
rect 193456 64280 340972 64308
rect 193456 64268 193462 64280
rect 340966 64268 340972 64280
rect 341024 64268 341030 64320
rect 203058 64200 203064 64252
rect 203116 64240 203122 64252
rect 472618 64240 472624 64252
rect 203116 64212 472624 64240
rect 203116 64200 203122 64212
rect 472618 64200 472624 64212
rect 472676 64200 472682 64252
rect 88334 64132 88340 64184
rect 88392 64172 88398 64184
rect 104158 64172 104164 64184
rect 88392 64144 104164 64172
rect 88392 64132 88398 64144
rect 104158 64132 104164 64144
rect 104216 64132 104222 64184
rect 147398 64132 147404 64184
rect 147456 64172 147462 64184
rect 183554 64172 183560 64184
rect 147456 64144 183560 64172
rect 147456 64132 147462 64144
rect 183554 64132 183560 64144
rect 183612 64132 183618 64184
rect 214374 64132 214380 64184
rect 214432 64172 214438 64184
rect 543734 64172 543740 64184
rect 214432 64144 543740 64172
rect 214432 64132 214438 64144
rect 543734 64132 543740 64144
rect 543792 64132 543798 64184
rect 144362 63996 144368 64048
rect 144420 64036 144426 64048
rect 147214 64036 147220 64048
rect 144420 64008 147220 64036
rect 144420 63996 144426 64008
rect 147214 63996 147220 64008
rect 147272 63996 147278 64048
rect 144086 63520 144092 63572
rect 144144 63560 144150 63572
rect 144270 63560 144276 63572
rect 144144 63532 144276 63560
rect 144144 63520 144150 63532
rect 144270 63520 144276 63532
rect 144328 63520 144334 63572
rect 100570 63452 100576 63504
rect 100628 63492 100634 63504
rect 134334 63492 134340 63504
rect 100628 63464 134340 63492
rect 100628 63452 100634 63464
rect 134334 63452 134340 63464
rect 134392 63452 134398 63504
rect 154758 63452 154764 63504
rect 154816 63492 154822 63504
rect 215478 63492 215484 63504
rect 154816 63464 215484 63492
rect 154816 63452 154822 63464
rect 215478 63452 215484 63464
rect 215536 63452 215542 63504
rect 104342 63384 104348 63436
rect 104400 63424 104406 63436
rect 104802 63424 104808 63436
rect 104400 63396 104808 63424
rect 104400 63384 104406 63396
rect 104802 63384 104808 63396
rect 104860 63424 104866 63436
rect 137186 63424 137192 63436
rect 104860 63396 137192 63424
rect 104860 63384 104866 63396
rect 137186 63384 137192 63396
rect 137244 63384 137250 63436
rect 168558 63384 168564 63436
rect 168616 63424 168622 63436
rect 169294 63424 169300 63436
rect 168616 63396 169300 63424
rect 168616 63384 168622 63396
rect 169294 63384 169300 63396
rect 169352 63424 169358 63436
rect 203610 63424 203616 63436
rect 169352 63396 203616 63424
rect 169352 63384 169358 63396
rect 203610 63384 203616 63396
rect 203668 63384 203674 63436
rect 157610 63316 157616 63368
rect 157668 63356 157674 63368
rect 192018 63356 192024 63368
rect 157668 63328 192024 63356
rect 157668 63316 157674 63328
rect 192018 63316 192024 63328
rect 192076 63356 192082 63368
rect 193030 63356 193036 63368
rect 192076 63328 193036 63356
rect 192076 63316 192082 63328
rect 193030 63316 193036 63328
rect 193088 63316 193094 63368
rect 168098 63248 168104 63300
rect 168156 63288 168162 63300
rect 201494 63288 201500 63300
rect 168156 63260 201500 63288
rect 168156 63248 168162 63260
rect 201494 63248 201500 63260
rect 201552 63248 201558 63300
rect 167454 62908 167460 62960
rect 167512 62948 167518 62960
rect 168098 62948 168104 62960
rect 167512 62920 168104 62948
rect 167512 62908 167518 62920
rect 168098 62908 168104 62920
rect 168156 62908 168162 62960
rect 72418 62840 72424 62892
rect 72476 62880 72482 62892
rect 104342 62880 104348 62892
rect 72476 62852 104348 62880
rect 72476 62840 72482 62852
rect 104342 62840 104348 62852
rect 104400 62840 104406 62892
rect 197630 62840 197636 62892
rect 197688 62880 197694 62892
rect 197814 62880 197820 62892
rect 197688 62852 197820 62880
rect 197688 62840 197694 62852
rect 197814 62840 197820 62852
rect 197872 62840 197878 62892
rect 215478 62840 215484 62892
rect 215536 62880 215542 62892
rect 292574 62880 292580 62892
rect 215536 62852 292580 62880
rect 215536 62840 215542 62852
rect 292574 62840 292580 62852
rect 292632 62840 292638 62892
rect 27614 62772 27620 62824
rect 27672 62812 27678 62824
rect 100570 62812 100576 62824
rect 27672 62784 100576 62812
rect 27672 62772 27678 62784
rect 100570 62772 100576 62784
rect 100628 62772 100634 62824
rect 108850 62772 108856 62824
rect 108908 62812 108914 62824
rect 115934 62812 115940 62824
rect 108908 62784 115940 62812
rect 108908 62772 108914 62784
rect 115934 62772 115940 62784
rect 115992 62812 115998 62824
rect 116946 62812 116952 62824
rect 115992 62784 116952 62812
rect 115992 62772 115998 62784
rect 116946 62772 116952 62784
rect 117004 62772 117010 62824
rect 138658 62772 138664 62824
rect 138716 62812 138722 62824
rect 142338 62812 142344 62824
rect 138716 62784 142344 62812
rect 138716 62772 138722 62784
rect 142338 62772 142344 62784
rect 142396 62772 142402 62824
rect 193030 62772 193036 62824
rect 193088 62812 193094 62824
rect 331214 62812 331220 62824
rect 193088 62784 331220 62812
rect 193088 62772 193094 62784
rect 331214 62772 331220 62784
rect 331272 62772 331278 62824
rect 103514 62704 103520 62756
rect 103572 62744 103578 62756
rect 108298 62744 108304 62756
rect 103572 62716 108304 62744
rect 103572 62704 103578 62716
rect 108298 62704 108304 62716
rect 108356 62704 108362 62756
rect 145926 62228 145932 62280
rect 145984 62268 145990 62280
rect 148318 62268 148324 62280
rect 145984 62240 148324 62268
rect 145984 62228 145990 62240
rect 148318 62228 148324 62240
rect 148376 62228 148382 62280
rect 106826 62024 106832 62076
rect 106884 62064 106890 62076
rect 117222 62064 117228 62076
rect 106884 62036 117228 62064
rect 106884 62024 106890 62036
rect 117222 62024 117228 62036
rect 117280 62024 117286 62076
rect 172698 62024 172704 62076
rect 172756 62064 172762 62076
rect 212534 62064 212540 62076
rect 172756 62036 212540 62064
rect 172756 62024 172762 62036
rect 212534 62024 212540 62036
rect 212592 62064 212598 62076
rect 213822 62064 213828 62076
rect 212592 62036 213828 62064
rect 212592 62024 212598 62036
rect 213822 62024 213828 62036
rect 213880 62024 213886 62076
rect 163222 61956 163228 62008
rect 163280 61996 163286 62008
rect 197630 61996 197636 62008
rect 163280 61968 197636 61996
rect 163280 61956 163286 61968
rect 197630 61956 197636 61968
rect 197688 61956 197694 62008
rect 151906 61548 151912 61600
rect 151964 61588 151970 61600
rect 251174 61588 251180 61600
rect 151964 61560 251180 61588
rect 151964 61548 151970 61560
rect 251174 61548 251180 61560
rect 251232 61548 251238 61600
rect 154482 61480 154488 61532
rect 154540 61520 154546 61532
rect 277394 61520 277400 61532
rect 154540 61492 277400 61520
rect 154540 61480 154546 61492
rect 277394 61480 277400 61492
rect 277452 61480 277458 61532
rect 197630 61412 197636 61464
rect 197688 61452 197694 61464
rect 394694 61452 394700 61464
rect 197688 61424 394700 61452
rect 197688 61412 197694 61424
rect 394694 61412 394700 61424
rect 394752 61412 394758 61464
rect 146386 61344 146392 61396
rect 146444 61384 146450 61396
rect 185578 61384 185584 61396
rect 146444 61356 185584 61384
rect 146444 61344 146450 61356
rect 185578 61344 185584 61356
rect 185636 61344 185642 61396
rect 213822 61344 213828 61396
rect 213880 61384 213886 61396
rect 529934 61384 529940 61396
rect 213880 61356 529940 61384
rect 213880 61344 213886 61356
rect 529934 61344 529940 61356
rect 529992 61344 529998 61396
rect 98638 60664 98644 60716
rect 98696 60704 98702 60716
rect 132954 60704 132960 60716
rect 98696 60676 132960 60704
rect 98696 60664 98702 60676
rect 132954 60664 132960 60676
rect 133012 60664 133018 60716
rect 145834 60664 145840 60716
rect 145892 60704 145898 60716
rect 152642 60704 152648 60716
rect 145892 60676 152648 60704
rect 145892 60664 145898 60676
rect 152642 60664 152648 60676
rect 152700 60664 152706 60716
rect 154666 60664 154672 60716
rect 154724 60704 154730 60716
rect 189074 60704 189080 60716
rect 154724 60676 189080 60704
rect 154724 60664 154730 60676
rect 189074 60664 189080 60676
rect 189132 60704 189138 60716
rect 189350 60704 189356 60716
rect 189132 60676 189356 60704
rect 189132 60664 189138 60676
rect 189350 60664 189356 60676
rect 189408 60664 189414 60716
rect 97994 60596 98000 60648
rect 98052 60636 98058 60648
rect 105906 60636 105912 60648
rect 98052 60608 105912 60636
rect 98052 60596 98058 60608
rect 105906 60596 105912 60608
rect 105964 60636 105970 60648
rect 139762 60636 139768 60648
rect 105964 60608 139768 60636
rect 105964 60596 105970 60608
rect 139762 60596 139768 60608
rect 139820 60596 139826 60648
rect 158898 60596 158904 60648
rect 158956 60636 158962 60648
rect 193306 60636 193312 60648
rect 158956 60608 193312 60636
rect 158956 60596 158962 60608
rect 193306 60596 193312 60608
rect 193364 60636 193370 60648
rect 194502 60636 194508 60648
rect 193364 60608 194508 60636
rect 193364 60596 193370 60608
rect 194502 60596 194508 60608
rect 194560 60596 194566 60648
rect 105814 60528 105820 60580
rect 105872 60568 105878 60580
rect 106090 60568 106096 60580
rect 105872 60540 106096 60568
rect 105872 60528 105878 60540
rect 106090 60528 106096 60540
rect 106148 60568 106154 60580
rect 137002 60568 137008 60580
rect 106148 60540 137008 60568
rect 106148 60528 106154 60540
rect 137002 60528 137008 60540
rect 137060 60528 137066 60580
rect 167362 60528 167368 60580
rect 167420 60568 167426 60580
rect 193674 60568 193680 60580
rect 167420 60540 193680 60568
rect 167420 60528 167426 60540
rect 193674 60528 193680 60540
rect 193732 60568 193738 60580
rect 194410 60568 194416 60580
rect 193732 60540 194416 60568
rect 193732 60528 193738 60540
rect 194410 60528 194416 60540
rect 194468 60528 194474 60580
rect 153102 60120 153108 60172
rect 153160 60160 153166 60172
rect 259454 60160 259460 60172
rect 153160 60132 259460 60160
rect 153160 60120 153166 60132
rect 259454 60120 259460 60132
rect 259512 60120 259518 60172
rect 62114 60052 62120 60104
rect 62172 60092 62178 60104
rect 105814 60092 105820 60104
rect 62172 60064 105820 60092
rect 62172 60052 62178 60064
rect 105814 60052 105820 60064
rect 105872 60052 105878 60104
rect 189074 60052 189080 60104
rect 189132 60092 189138 60104
rect 299474 60092 299480 60104
rect 189132 60064 299480 60092
rect 189132 60052 189138 60064
rect 299474 60052 299480 60064
rect 299532 60052 299538 60104
rect 21358 59984 21364 60036
rect 21416 60024 21422 60036
rect 98638 60024 98644 60036
rect 21416 59996 98644 60024
rect 21416 59984 21422 59996
rect 98638 59984 98644 59996
rect 98696 59984 98702 60036
rect 147306 59984 147312 60036
rect 147364 60024 147370 60036
rect 187694 60024 187700 60036
rect 147364 59996 187700 60024
rect 147364 59984 147370 59996
rect 187694 59984 187700 59996
rect 187752 59984 187758 60036
rect 194502 59984 194508 60036
rect 194560 60024 194566 60036
rect 349154 60024 349160 60036
rect 194560 59996 349160 60024
rect 194560 59984 194566 59996
rect 349154 59984 349160 59996
rect 349212 59984 349218 60036
rect 140130 59780 140136 59832
rect 140188 59820 140194 59832
rect 142522 59820 142528 59832
rect 140188 59792 142528 59820
rect 140188 59780 140194 59792
rect 142522 59780 142528 59792
rect 142580 59780 142586 59832
rect 194410 59372 194416 59424
rect 194468 59412 194474 59424
rect 459554 59412 459560 59424
rect 194468 59384 459560 59412
rect 194468 59372 194474 59384
rect 459554 59372 459560 59384
rect 459612 59372 459618 59424
rect 100754 59304 100760 59356
rect 100812 59344 100818 59356
rect 101858 59344 101864 59356
rect 100812 59316 101864 59344
rect 100812 59304 100818 59316
rect 101858 59304 101864 59316
rect 101916 59344 101922 59356
rect 135714 59344 135720 59356
rect 101916 59316 135720 59344
rect 101916 59304 101922 59316
rect 135714 59304 135720 59316
rect 135772 59304 135778 59356
rect 167178 59304 167184 59356
rect 167236 59344 167242 59356
rect 201770 59344 201776 59356
rect 167236 59316 201776 59344
rect 167236 59304 167242 59316
rect 201770 59304 201776 59316
rect 201828 59344 201834 59356
rect 202782 59344 202788 59356
rect 201828 59316 202788 59344
rect 201828 59304 201834 59316
rect 202782 59304 202788 59316
rect 202840 59304 202846 59356
rect 157518 59236 157524 59288
rect 157576 59276 157582 59288
rect 192754 59276 192760 59288
rect 157576 59248 192760 59276
rect 157576 59236 157582 59248
rect 192754 59236 192760 59248
rect 192812 59276 192818 59288
rect 193030 59276 193036 59288
rect 192812 59248 193036 59276
rect 192812 59236 192818 59248
rect 193030 59236 193036 59248
rect 193088 59236 193094 59288
rect 193030 58692 193036 58744
rect 193088 58732 193094 58744
rect 327074 58732 327080 58744
rect 193088 58704 327080 58732
rect 193088 58692 193094 58704
rect 327074 58692 327080 58704
rect 327132 58692 327138 58744
rect 48314 58624 48320 58676
rect 48372 58664 48378 58676
rect 100754 58664 100760 58676
rect 48372 58636 100760 58664
rect 48372 58624 48378 58636
rect 100754 58624 100760 58636
rect 100812 58624 100818 58676
rect 202782 58624 202788 58676
rect 202840 58664 202846 58676
rect 448514 58664 448520 58676
rect 202840 58636 448520 58664
rect 202840 58624 202846 58636
rect 448514 58624 448520 58636
rect 448572 58624 448578 58676
rect 168466 57876 168472 57928
rect 168524 57916 168530 57928
rect 203242 57916 203248 57928
rect 168524 57888 203248 57916
rect 168524 57876 168530 57888
rect 203242 57876 203248 57888
rect 203300 57916 203306 57928
rect 204162 57916 204168 57928
rect 203300 57888 204168 57916
rect 203300 57876 203306 57888
rect 204162 57876 204168 57888
rect 204220 57876 204226 57928
rect 160186 57808 160192 57860
rect 160244 57848 160250 57860
rect 194686 57848 194692 57860
rect 160244 57820 194692 57848
rect 160244 57808 160250 57820
rect 194686 57808 194692 57820
rect 194744 57848 194750 57860
rect 195054 57848 195060 57860
rect 194744 57820 195060 57848
rect 194744 57808 194750 57820
rect 195054 57808 195060 57820
rect 195112 57808 195118 57860
rect 156138 57740 156144 57792
rect 156196 57780 156202 57792
rect 190454 57780 190460 57792
rect 156196 57752 190460 57780
rect 156196 57740 156202 57752
rect 190454 57740 190460 57752
rect 190512 57780 190518 57792
rect 191742 57780 191748 57792
rect 190512 57752 191748 57780
rect 190512 57740 190518 57752
rect 191742 57740 191748 57752
rect 191800 57740 191806 57792
rect 153010 57400 153016 57452
rect 153068 57440 153074 57452
rect 263594 57440 263600 57452
rect 153068 57412 263600 57440
rect 153068 57400 153074 57412
rect 263594 57400 263600 57412
rect 263652 57400 263658 57452
rect 191742 57332 191748 57384
rect 191800 57372 191806 57384
rect 309134 57372 309140 57384
rect 191800 57344 309140 57372
rect 191800 57332 191806 57344
rect 309134 57332 309140 57344
rect 309192 57332 309198 57384
rect 195054 57264 195060 57316
rect 195112 57304 195118 57316
rect 362954 57304 362960 57316
rect 195112 57276 362960 57304
rect 195112 57264 195118 57276
rect 362954 57264 362960 57276
rect 363012 57264 363018 57316
rect 204162 57196 204168 57248
rect 204220 57236 204226 57248
rect 473446 57236 473452 57248
rect 204220 57208 473452 57236
rect 204220 57196 204226 57208
rect 473446 57196 473452 57208
rect 473504 57196 473510 57248
rect 178770 56516 178776 56568
rect 178828 56556 178834 56568
rect 217042 56556 217048 56568
rect 178828 56528 217048 56556
rect 178828 56516 178834 56528
rect 217042 56516 217048 56528
rect 217100 56516 217106 56568
rect 166994 56448 167000 56500
rect 167052 56488 167058 56500
rect 201862 56488 201868 56500
rect 167052 56460 201868 56488
rect 167052 56448 167058 56460
rect 201862 56448 201868 56460
rect 201920 56488 201926 56500
rect 202782 56488 202788 56500
rect 201920 56460 202788 56488
rect 201920 56448 201926 56460
rect 202782 56448 202788 56460
rect 202840 56448 202846 56500
rect 163130 56380 163136 56432
rect 163188 56420 163194 56432
rect 197630 56420 197636 56432
rect 163188 56392 197636 56420
rect 163188 56380 163194 56392
rect 197630 56380 197636 56392
rect 197688 56380 197694 56432
rect 158806 56312 158812 56364
rect 158864 56352 158870 56364
rect 193214 56352 193220 56364
rect 158864 56324 193220 56352
rect 158864 56312 158870 56324
rect 193214 56312 193220 56324
rect 193272 56352 193278 56364
rect 194502 56352 194508 56364
rect 193272 56324 194508 56352
rect 193272 56312 193278 56324
rect 194502 56312 194508 56324
rect 194560 56312 194566 56364
rect 156046 56244 156052 56296
rect 156104 56284 156110 56296
rect 189074 56284 189080 56296
rect 156104 56256 189080 56284
rect 156104 56244 156110 56256
rect 189074 56244 189080 56256
rect 189132 56244 189138 56296
rect 150250 56176 150256 56228
rect 150308 56216 150314 56228
rect 220078 56216 220084 56228
rect 150308 56188 220084 56216
rect 150308 56176 150314 56188
rect 220078 56176 220084 56188
rect 220136 56176 220142 56228
rect 189074 56108 189080 56160
rect 189132 56148 189138 56160
rect 313274 56148 313280 56160
rect 189132 56120 313280 56148
rect 189132 56108 189138 56120
rect 313274 56108 313280 56120
rect 313332 56108 313338 56160
rect 194502 56040 194508 56092
rect 194560 56080 194566 56092
rect 351914 56080 351920 56092
rect 194560 56052 351920 56080
rect 194560 56040 194566 56052
rect 351914 56040 351920 56052
rect 351972 56040 351978 56092
rect 197630 55972 197636 56024
rect 197688 56012 197694 56024
rect 398834 56012 398840 56024
rect 197688 55984 398840 56012
rect 197688 55972 197694 55984
rect 398834 55972 398840 55984
rect 398892 55972 398898 56024
rect 202782 55904 202788 55956
rect 202840 55944 202846 55956
rect 448606 55944 448612 55956
rect 202840 55916 448612 55944
rect 202840 55904 202846 55916
rect 448606 55904 448612 55916
rect 448664 55904 448670 55956
rect 217042 55836 217048 55888
rect 217100 55876 217106 55888
rect 564526 55876 564532 55888
rect 217100 55848 564532 55876
rect 217100 55836 217106 55848
rect 564526 55836 564532 55848
rect 564584 55836 564590 55888
rect 109586 55156 109592 55208
rect 109644 55196 109650 55208
rect 138382 55196 138388 55208
rect 109644 55168 138388 55196
rect 109644 55156 109650 55168
rect 138382 55156 138388 55168
rect 138440 55156 138446 55208
rect 164326 55156 164332 55208
rect 164384 55196 164390 55208
rect 198826 55196 198832 55208
rect 164384 55168 198832 55196
rect 164384 55156 164390 55168
rect 198826 55156 198832 55168
rect 198884 55156 198890 55208
rect 168374 55088 168380 55140
rect 168432 55128 168438 55140
rect 202874 55128 202880 55140
rect 168432 55100 202880 55128
rect 168432 55088 168438 55100
rect 202874 55088 202880 55100
rect 202932 55088 202938 55140
rect 198826 54544 198832 54596
rect 198884 54584 198890 54596
rect 414658 54584 414664 54596
rect 198884 54556 414664 54584
rect 198884 54544 198890 54556
rect 414658 54544 414664 54556
rect 414716 54544 414722 54596
rect 202874 54476 202880 54528
rect 202932 54516 202938 54528
rect 464338 54516 464344 54528
rect 202932 54488 464344 54516
rect 202932 54476 202938 54488
rect 464338 54476 464344 54488
rect 464396 54476 464402 54528
rect 172054 53728 172060 53780
rect 172112 53768 172118 53780
rect 204254 53768 204260 53780
rect 172112 53740 204260 53768
rect 172112 53728 172118 53740
rect 204254 53728 204260 53740
rect 204312 53728 204318 53780
rect 166258 53660 166264 53712
rect 166316 53700 166322 53712
rect 198090 53700 198096 53712
rect 166316 53672 198096 53700
rect 166316 53660 166322 53672
rect 198090 53660 198096 53672
rect 198148 53660 198154 53712
rect 151630 53184 151636 53236
rect 151688 53224 151694 53236
rect 242894 53224 242900 53236
rect 151688 53196 242900 53224
rect 151688 53184 151694 53196
rect 242894 53184 242900 53196
rect 242952 53184 242958 53236
rect 198090 53116 198096 53168
rect 198148 53156 198154 53168
rect 402974 53156 402980 53168
rect 198148 53128 402980 53156
rect 198148 53116 198154 53128
rect 402974 53116 402980 53128
rect 403032 53116 403038 53168
rect 204254 53048 204260 53100
rect 204312 53088 204318 53100
rect 490006 53088 490012 53100
rect 204312 53060 490012 53088
rect 204312 53048 204318 53060
rect 490006 53048 490012 53060
rect 490064 53048 490070 53100
rect 197446 52504 197452 52556
rect 197504 52544 197510 52556
rect 197630 52544 197636 52556
rect 197504 52516 197636 52544
rect 197504 52504 197510 52516
rect 197630 52504 197636 52516
rect 197688 52504 197694 52556
rect 155954 52368 155960 52420
rect 156012 52408 156018 52420
rect 189626 52408 189632 52420
rect 156012 52380 189632 52408
rect 156012 52368 156018 52380
rect 189626 52368 189632 52380
rect 189684 52368 189690 52420
rect 150158 51688 150164 51740
rect 150216 51728 150222 51740
rect 217318 51728 217324 51740
rect 150216 51700 217324 51728
rect 150216 51688 150222 51700
rect 217318 51688 217324 51700
rect 217376 51688 217382 51740
rect 189626 51076 189632 51128
rect 189684 51116 189690 51128
rect 320174 51116 320180 51128
rect 189684 51088 320180 51116
rect 189684 51076 189690 51088
rect 320174 51076 320180 51088
rect 320232 51076 320238 51128
rect 157426 51008 157432 51060
rect 157484 51048 157490 51060
rect 192662 51048 192668 51060
rect 157484 51020 192668 51048
rect 157484 51008 157490 51020
rect 192662 51008 192668 51020
rect 192720 51048 192726 51060
rect 193030 51048 193036 51060
rect 192720 51020 193036 51048
rect 192720 51008 192726 51020
rect 193030 51008 193036 51020
rect 193088 51008 193094 51060
rect 176838 50940 176844 50992
rect 176896 50980 176902 50992
rect 208486 50980 208492 50992
rect 176896 50952 208492 50980
rect 176896 50940 176902 50952
rect 208486 50940 208492 50952
rect 208544 50940 208550 50992
rect 193030 50396 193036 50448
rect 193088 50436 193094 50448
rect 338114 50436 338120 50448
rect 193088 50408 338120 50436
rect 193088 50396 193094 50408
rect 338114 50396 338120 50408
rect 338172 50396 338178 50448
rect 110414 50328 110420 50380
rect 110472 50368 110478 50380
rect 119338 50368 119344 50380
rect 110472 50340 119344 50368
rect 110472 50328 110478 50340
rect 119338 50328 119344 50340
rect 119396 50328 119402 50380
rect 145742 50328 145748 50380
rect 145800 50368 145806 50380
rect 167638 50368 167644 50380
rect 145800 50340 167644 50368
rect 145800 50328 145806 50340
rect 167638 50328 167644 50340
rect 167696 50328 167702 50380
rect 208486 50328 208492 50380
rect 208544 50368 208550 50380
rect 209130 50368 209136 50380
rect 208544 50340 209136 50368
rect 208544 50328 208550 50340
rect 209130 50328 209136 50340
rect 209188 50368 209194 50380
rect 569954 50368 569960 50380
rect 209188 50340 569960 50368
rect 209188 50328 209194 50340
rect 569954 50328 569960 50340
rect 570012 50328 570018 50380
rect 143810 49648 143816 49700
rect 143868 49688 143874 49700
rect 148410 49688 148416 49700
rect 143868 49660 148416 49688
rect 143868 49648 143874 49660
rect 148410 49648 148416 49660
rect 148468 49648 148474 49700
rect 154574 49648 154580 49700
rect 154632 49688 154638 49700
rect 189442 49688 189448 49700
rect 154632 49660 189448 49688
rect 154632 49648 154638 49660
rect 189442 49648 189448 49660
rect 189500 49648 189506 49700
rect 147674 49104 147680 49156
rect 147732 49144 147738 49156
rect 201586 49144 201592 49156
rect 147732 49116 201592 49144
rect 147732 49104 147738 49116
rect 201586 49104 201592 49116
rect 201644 49104 201650 49156
rect 189442 48968 189448 49020
rect 189500 49008 189506 49020
rect 190178 49008 190184 49020
rect 189500 48980 190184 49008
rect 189500 48968 189506 48980
rect 190178 48968 190184 48980
rect 190236 49008 190242 49020
rect 285674 49008 285680 49020
rect 190236 48980 285680 49008
rect 190236 48968 190242 48980
rect 285674 48968 285680 48980
rect 285732 48968 285738 49020
rect 148686 47608 148692 47660
rect 148744 47648 148750 47660
rect 204254 47648 204260 47660
rect 148744 47620 204260 47648
rect 148744 47608 148750 47620
rect 204254 47608 204260 47620
rect 204312 47608 204318 47660
rect 150066 47540 150072 47592
rect 150124 47580 150130 47592
rect 215294 47580 215300 47592
rect 150124 47552 215300 47580
rect 150124 47540 150130 47552
rect 215294 47540 215300 47552
rect 215352 47540 215358 47592
rect 135254 46928 135260 46980
rect 135312 46968 135318 46980
rect 142430 46968 142436 46980
rect 135312 46940 142436 46968
rect 135312 46928 135318 46940
rect 142430 46928 142436 46940
rect 142488 46928 142494 46980
rect 176746 46860 176752 46912
rect 176804 46900 176810 46912
rect 208486 46900 208492 46912
rect 176804 46872 208492 46900
rect 176804 46860 176810 46872
rect 208486 46860 208492 46872
rect 208544 46900 208550 46912
rect 209038 46900 209044 46912
rect 208544 46872 209044 46900
rect 208544 46860 208550 46872
rect 209038 46860 209044 46872
rect 209096 46860 209102 46912
rect 151538 46248 151544 46300
rect 151596 46288 151602 46300
rect 233234 46288 233240 46300
rect 151596 46260 233240 46288
rect 151596 46248 151602 46260
rect 233234 46248 233240 46260
rect 233292 46248 233298 46300
rect 208486 46180 208492 46232
rect 208544 46220 208550 46232
rect 571978 46220 571984 46232
rect 208544 46192 571984 46220
rect 208544 46180 208550 46192
rect 571978 46180 571984 46192
rect 572036 46180 572042 46232
rect 172606 45500 172612 45552
rect 172664 45540 172670 45552
rect 205910 45540 205916 45552
rect 172664 45512 205916 45540
rect 172664 45500 172670 45512
rect 205910 45500 205916 45512
rect 205968 45500 205974 45552
rect 148594 44820 148600 44872
rect 148652 44860 148658 44872
rect 198734 44860 198740 44872
rect 148652 44832 198740 44860
rect 148652 44820 148658 44832
rect 198734 44820 198740 44832
rect 198792 44820 198798 44872
rect 205910 44140 205916 44192
rect 205968 44180 205974 44192
rect 520918 44180 520924 44192
rect 205968 44152 520924 44180
rect 205968 44140 205974 44152
rect 520918 44140 520924 44152
rect 520976 44140 520982 44192
rect 176654 44072 176660 44124
rect 176712 44112 176718 44124
rect 210142 44112 210148 44124
rect 176712 44084 210148 44112
rect 176712 44072 176718 44084
rect 210142 44072 210148 44084
rect 210200 44112 210206 44124
rect 211062 44112 211068 44124
rect 210200 44084 211068 44112
rect 210200 44072 210206 44084
rect 211062 44072 211068 44084
rect 211120 44072 211126 44124
rect 152918 43528 152924 43580
rect 152976 43568 152982 43580
rect 267734 43568 267740 43580
rect 152976 43540 267740 43568
rect 152976 43528 152982 43540
rect 267734 43528 267740 43540
rect 267792 43528 267798 43580
rect 163038 43460 163044 43512
rect 163096 43500 163102 43512
rect 408494 43500 408500 43512
rect 163096 43472 408500 43500
rect 163096 43460 163102 43472
rect 408494 43460 408500 43472
rect 408552 43460 408558 43512
rect 167270 43392 167276 43444
rect 167328 43432 167334 43444
rect 458174 43432 458180 43444
rect 167328 43404 458180 43432
rect 167328 43392 167334 43404
rect 458174 43392 458180 43404
rect 458232 43392 458238 43444
rect 211062 42780 211068 42832
rect 211120 42820 211126 42832
rect 576854 42820 576860 42832
rect 211120 42792 576860 42820
rect 211120 42780 211126 42792
rect 576854 42780 576860 42792
rect 576912 42780 576918 42832
rect 151446 42304 151452 42356
rect 151504 42344 151510 42356
rect 239398 42344 239404 42356
rect 151504 42316 239404 42344
rect 151504 42304 151510 42316
rect 239398 42304 239404 42316
rect 239456 42304 239462 42356
rect 159726 42236 159732 42288
rect 159784 42276 159790 42288
rect 350534 42276 350540 42288
rect 159784 42248 350540 42276
rect 159784 42236 159790 42248
rect 350534 42236 350540 42248
rect 350592 42236 350598 42288
rect 164234 42168 164240 42220
rect 164292 42208 164298 42220
rect 426434 42208 426440 42220
rect 164292 42180 426440 42208
rect 164292 42168 164298 42180
rect 426434 42168 426440 42180
rect 426492 42168 426498 42220
rect 166350 42100 166356 42152
rect 166408 42140 166414 42152
rect 438854 42140 438860 42152
rect 166408 42112 438860 42140
rect 166408 42100 166414 42112
rect 438854 42100 438860 42112
rect 438912 42100 438918 42152
rect 70394 42032 70400 42084
rect 70452 42072 70458 42084
rect 136634 42072 136640 42084
rect 70452 42044 136640 42072
rect 70452 42032 70458 42044
rect 136634 42032 136640 42044
rect 136692 42032 136698 42084
rect 145558 42032 145564 42084
rect 145616 42072 145622 42084
rect 166994 42072 167000 42084
rect 145616 42044 167000 42072
rect 145616 42032 145622 42044
rect 166994 42032 167000 42044
rect 167052 42032 167058 42084
rect 169754 42032 169760 42084
rect 169812 42072 169818 42084
rect 495434 42072 495440 42084
rect 169812 42044 495440 42072
rect 169812 42032 169818 42044
rect 495434 42032 495440 42044
rect 495492 42032 495498 42084
rect 156598 40876 156604 40928
rect 156656 40916 156662 40928
rect 307018 40916 307024 40928
rect 156656 40888 307024 40916
rect 156656 40876 156662 40888
rect 307018 40876 307024 40888
rect 307076 40876 307082 40928
rect 167086 40808 167092 40860
rect 167144 40848 167150 40860
rect 462314 40848 462320 40860
rect 167144 40820 462320 40848
rect 167144 40808 167150 40820
rect 462314 40808 462320 40820
rect 462372 40808 462378 40860
rect 172238 40740 172244 40792
rect 172296 40780 172302 40792
rect 498286 40780 498292 40792
rect 172296 40752 498292 40780
rect 172296 40740 172302 40752
rect 498286 40740 498292 40752
rect 498344 40740 498350 40792
rect 174906 40672 174912 40724
rect 174964 40712 174970 40724
rect 535454 40712 535460 40724
rect 174964 40684 535460 40712
rect 174964 40672 174970 40684
rect 535454 40672 535460 40684
rect 535512 40672 535518 40724
rect 177482 39992 177488 40044
rect 177540 40032 177546 40044
rect 213914 40032 213920 40044
rect 177540 40004 213920 40032
rect 177540 39992 177546 40004
rect 213914 39992 213920 40004
rect 213972 40032 213978 40044
rect 214374 40032 214380 40044
rect 213972 40004 214380 40032
rect 213972 39992 213978 40004
rect 214374 39992 214380 40004
rect 214432 39992 214438 40044
rect 151354 39584 151360 39636
rect 151412 39624 151418 39636
rect 235994 39624 236000 39636
rect 151412 39596 236000 39624
rect 151412 39584 151418 39596
rect 235994 39584 236000 39596
rect 236052 39584 236058 39636
rect 165062 39516 165068 39568
rect 165120 39556 165126 39568
rect 409874 39556 409880 39568
rect 165120 39528 409880 39556
rect 165120 39516 165126 39528
rect 409874 39516 409880 39528
rect 409932 39516 409938 39568
rect 214374 39448 214380 39500
rect 214432 39488 214438 39500
rect 518894 39488 518900 39500
rect 214432 39460 518900 39488
rect 214432 39448 214438 39460
rect 518894 39448 518900 39460
rect 518952 39448 518958 39500
rect 173526 39380 173532 39432
rect 173584 39420 173590 39432
rect 516134 39420 516140 39432
rect 173584 39392 516140 39420
rect 173584 39380 173590 39392
rect 516134 39380 516140 39392
rect 516192 39380 516198 39432
rect 77386 39312 77392 39364
rect 77444 39352 77450 39364
rect 138290 39352 138296 39364
rect 77444 39324 138296 39352
rect 77444 39312 77450 39324
rect 138290 39312 138296 39324
rect 138348 39312 138354 39364
rect 176102 39312 176108 39364
rect 176160 39352 176166 39364
rect 558914 39352 558920 39364
rect 176160 39324 558920 39352
rect 176160 39312 176166 39324
rect 558914 39312 558920 39324
rect 558972 39312 558978 39364
rect 138014 38972 138020 39024
rect 138072 39012 138078 39024
rect 142890 39012 142896 39024
rect 138072 38984 142896 39012
rect 138072 38972 138078 38984
rect 142890 38972 142896 38984
rect 142948 38972 142954 39024
rect 152826 38088 152832 38140
rect 152884 38128 152890 38140
rect 257338 38128 257344 38140
rect 152884 38100 257344 38128
rect 152884 38088 152890 38100
rect 257338 38088 257344 38100
rect 257396 38088 257402 38140
rect 169386 38020 169392 38072
rect 169444 38060 169450 38072
rect 463694 38060 463700 38072
rect 169444 38032 463700 38060
rect 169444 38020 169450 38032
rect 463694 38020 463700 38032
rect 463752 38020 463758 38072
rect 169478 37952 169484 38004
rect 169536 37992 169542 38004
rect 476114 37992 476120 38004
rect 169536 37964 476120 37992
rect 169536 37952 169542 37964
rect 476114 37952 476120 37964
rect 476172 37952 476178 38004
rect 13814 37884 13820 37936
rect 13872 37924 13878 37936
rect 132770 37924 132776 37936
rect 13872 37896 132776 37924
rect 13872 37884 13878 37896
rect 132770 37884 132776 37896
rect 132828 37884 132834 37936
rect 145650 37884 145656 37936
rect 145708 37924 145714 37936
rect 168466 37924 168472 37936
rect 145708 37896 168472 37924
rect 145708 37884 145714 37896
rect 168466 37884 168472 37896
rect 168524 37884 168530 37936
rect 172514 37884 172520 37936
rect 172572 37924 172578 37936
rect 525058 37924 525064 37936
rect 172572 37896 525064 37924
rect 172572 37884 172578 37896
rect 525058 37884 525064 37896
rect 525116 37884 525122 37936
rect 148502 36864 148508 36916
rect 148560 36904 148566 36916
rect 205634 36904 205640 36916
rect 148560 36876 205640 36904
rect 148560 36864 148566 36876
rect 205634 36864 205640 36876
rect 205692 36864 205698 36916
rect 154390 36796 154396 36848
rect 154448 36836 154454 36848
rect 267826 36836 267832 36848
rect 154448 36808 267832 36836
rect 154448 36796 154454 36808
rect 267826 36796 267832 36808
rect 267884 36796 267890 36848
rect 162210 36728 162216 36780
rect 162268 36768 162274 36780
rect 361574 36768 361580 36780
rect 162268 36740 361580 36768
rect 162268 36728 162274 36740
rect 361574 36728 361580 36740
rect 361632 36728 361638 36780
rect 170490 36660 170496 36712
rect 170548 36700 170554 36712
rect 481634 36700 481640 36712
rect 170548 36672 481640 36700
rect 170548 36660 170554 36672
rect 481634 36660 481640 36672
rect 481692 36660 481698 36712
rect 172146 36592 172152 36644
rect 172204 36632 172210 36644
rect 503714 36632 503720 36644
rect 172204 36604 503720 36632
rect 172204 36592 172210 36604
rect 503714 36592 503720 36604
rect 503772 36592 503778 36644
rect 174998 36524 175004 36576
rect 175056 36564 175062 36576
rect 534074 36564 534080 36576
rect 175056 36536 534080 36564
rect 175056 36524 175062 36536
rect 534074 36524 534080 36536
rect 534132 36524 534138 36576
rect 169294 35232 169300 35284
rect 169352 35272 169358 35284
rect 467834 35272 467840 35284
rect 169352 35244 467840 35272
rect 169352 35232 169358 35244
rect 467834 35232 467840 35244
rect 467892 35232 467898 35284
rect 31754 35164 31760 35216
rect 31812 35204 31818 35216
rect 133966 35204 133972 35216
rect 31812 35176 133972 35204
rect 31812 35164 31818 35176
rect 133966 35164 133972 35176
rect 134024 35164 134030 35216
rect 175274 35164 175280 35216
rect 175332 35204 175338 35216
rect 552014 35204 552020 35216
rect 175332 35176 552020 35204
rect 175332 35164 175338 35176
rect 552014 35164 552020 35176
rect 552072 35164 552078 35216
rect 159910 34008 159916 34060
rect 159968 34048 159974 34060
rect 346394 34048 346400 34060
rect 159968 34020 346400 34048
rect 159968 34008 159974 34020
rect 346394 34008 346400 34020
rect 346452 34008 346458 34060
rect 168098 33940 168104 33992
rect 168156 33980 168162 33992
rect 446398 33980 446404 33992
rect 168156 33952 446404 33980
rect 168156 33940 168162 33952
rect 446398 33940 446404 33952
rect 446456 33940 446462 33992
rect 170674 33872 170680 33924
rect 170732 33912 170738 33924
rect 488534 33912 488540 33924
rect 170732 33884 488540 33912
rect 170732 33872 170738 33884
rect 488534 33872 488540 33884
rect 488592 33872 488598 33924
rect 144270 33804 144276 33856
rect 144328 33844 144334 33856
rect 145006 33844 145012 33856
rect 144328 33816 145012 33844
rect 144328 33804 144334 33816
rect 145006 33804 145012 33816
rect 145064 33804 145070 33856
rect 176194 33804 176200 33856
rect 176252 33844 176258 33856
rect 565814 33844 565820 33856
rect 176252 33816 565820 33844
rect 176252 33804 176258 33816
rect 565814 33804 565820 33816
rect 565872 33804 565878 33856
rect 45554 33736 45560 33788
rect 45612 33776 45618 33788
rect 135346 33776 135352 33788
rect 45612 33748 135352 33776
rect 45612 33736 45618 33748
rect 135346 33736 135352 33748
rect 135404 33736 135410 33788
rect 145466 33736 145472 33788
rect 145524 33776 145530 33788
rect 171778 33776 171784 33788
rect 145524 33748 171784 33776
rect 145524 33736 145530 33748
rect 171778 33736 171784 33748
rect 171836 33736 171842 33788
rect 177666 33736 177672 33788
rect 177724 33776 177730 33788
rect 578234 33776 578240 33788
rect 177724 33748 578240 33776
rect 177724 33736 177730 33748
rect 578234 33736 578240 33748
rect 578292 33736 578298 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 95878 33096 95884 33108
rect 3568 33068 95884 33096
rect 3568 33056 3574 33068
rect 95878 33056 95884 33068
rect 95936 33056 95942 33108
rect 149974 32512 149980 32564
rect 150032 32552 150038 32564
rect 225598 32552 225604 32564
rect 150032 32524 225604 32552
rect 150032 32512 150038 32524
rect 225598 32512 225604 32524
rect 225656 32512 225662 32564
rect 151722 32444 151728 32496
rect 151780 32484 151786 32496
rect 242986 32484 242992 32496
rect 151780 32456 242992 32484
rect 151780 32444 151786 32456
rect 242986 32444 242992 32456
rect 243044 32444 243050 32496
rect 159818 32376 159824 32428
rect 159876 32416 159882 32428
rect 339494 32416 339500 32428
rect 159876 32388 339500 32416
rect 159876 32376 159882 32388
rect 339494 32376 339500 32388
rect 339552 32376 339558 32428
rect 152734 31152 152740 31204
rect 152792 31192 152798 31204
rect 264974 31192 264980 31204
rect 152792 31164 264980 31192
rect 152792 31152 152798 31164
rect 264974 31152 264980 31164
rect 265032 31152 265038 31204
rect 160922 31084 160928 31136
rect 160980 31124 160986 31136
rect 357434 31124 357440 31136
rect 160980 31096 357440 31124
rect 160980 31084 160986 31096
rect 357434 31084 357440 31096
rect 357492 31084 357498 31136
rect 17310 31016 17316 31068
rect 17368 31056 17374 31068
rect 132862 31056 132868 31068
rect 17368 31028 132868 31056
rect 17368 31016 17374 31028
rect 132862 31016 132868 31028
rect 132920 31016 132926 31068
rect 169570 31016 169576 31068
rect 169628 31056 169634 31068
rect 470594 31056 470600 31068
rect 169628 31028 470600 31056
rect 169628 31016 169634 31028
rect 470594 31016 470600 31028
rect 470652 31016 470658 31068
rect 155586 29792 155592 29844
rect 155644 29832 155650 29844
rect 299566 29832 299572 29844
rect 155644 29804 299572 29832
rect 155644 29792 155650 29804
rect 299566 29792 299572 29804
rect 299624 29792 299630 29844
rect 162946 29724 162952 29776
rect 163004 29764 163010 29776
rect 407206 29764 407212 29776
rect 163004 29736 407212 29764
rect 163004 29724 163010 29736
rect 407206 29724 407212 29736
rect 407264 29724 407270 29776
rect 170766 29656 170772 29708
rect 170824 29696 170830 29708
rect 491294 29696 491300 29708
rect 170824 29668 491300 29696
rect 170824 29656 170830 29668
rect 491294 29656 491300 29668
rect 491352 29656 491358 29708
rect 24854 29588 24860 29640
rect 24912 29628 24918 29640
rect 134150 29628 134156 29640
rect 24912 29600 134156 29628
rect 24912 29588 24918 29600
rect 134150 29588 134156 29600
rect 134208 29588 134214 29640
rect 177758 29588 177764 29640
rect 177816 29628 177822 29640
rect 574094 29628 574100 29640
rect 177816 29600 574100 29628
rect 177816 29588 177822 29600
rect 574094 29588 574100 29600
rect 574152 29588 574158 29640
rect 158346 28432 158352 28484
rect 158404 28472 158410 28484
rect 321554 28472 321560 28484
rect 158404 28444 321560 28472
rect 158404 28432 158410 28444
rect 321554 28432 321560 28444
rect 321612 28432 321618 28484
rect 166442 28364 166448 28416
rect 166500 28404 166506 28416
rect 427814 28404 427820 28416
rect 166500 28376 427820 28404
rect 166500 28364 166506 28376
rect 427814 28364 427820 28376
rect 427872 28364 427878 28416
rect 171318 28296 171324 28348
rect 171376 28336 171382 28348
rect 502334 28336 502340 28348
rect 171376 28308 502340 28336
rect 171376 28296 171382 28308
rect 502334 28296 502340 28308
rect 502392 28296 502398 28348
rect 184842 28228 184848 28280
rect 184900 28268 184906 28280
rect 582374 28268 582380 28280
rect 184900 28240 582380 28268
rect 184900 28228 184906 28240
rect 582374 28228 582380 28240
rect 582432 28228 582438 28280
rect 154206 27140 154212 27192
rect 154264 27180 154270 27192
rect 275278 27180 275284 27192
rect 154264 27152 275284 27180
rect 154264 27140 154270 27152
rect 275278 27140 275284 27152
rect 275336 27140 275342 27192
rect 162302 27072 162308 27124
rect 162360 27112 162366 27124
rect 374086 27112 374092 27124
rect 162360 27084 374092 27112
rect 162360 27072 162366 27084
rect 374086 27072 374092 27084
rect 374144 27072 374150 27124
rect 165154 27004 165160 27056
rect 165212 27044 165218 27056
rect 410518 27044 410524 27056
rect 165212 27016 410524 27044
rect 165212 27004 165218 27016
rect 410518 27004 410524 27016
rect 410576 27004 410582 27056
rect 171226 26936 171232 26988
rect 171284 26976 171290 26988
rect 506566 26976 506572 26988
rect 171284 26948 506572 26976
rect 171284 26936 171290 26948
rect 506566 26936 506572 26948
rect 506624 26936 506630 26988
rect 144914 26868 144920 26920
rect 144972 26908 144978 26920
rect 171870 26908 171876 26920
rect 144972 26880 171876 26908
rect 144972 26868 144978 26880
rect 171870 26868 171876 26880
rect 171928 26868 171934 26920
rect 172330 26868 172336 26920
rect 172388 26908 172394 26920
rect 510614 26908 510620 26920
rect 172388 26880 510620 26908
rect 172388 26868 172394 26880
rect 510614 26868 510620 26880
rect 510672 26868 510678 26920
rect 154114 25780 154120 25832
rect 154172 25820 154178 25832
rect 278774 25820 278780 25832
rect 154172 25792 278780 25820
rect 154172 25780 154178 25792
rect 278774 25780 278780 25792
rect 278832 25780 278838 25832
rect 162394 25712 162400 25764
rect 162452 25752 162458 25764
rect 378134 25752 378140 25764
rect 162452 25724 378140 25752
rect 162452 25712 162458 25724
rect 378134 25712 378140 25724
rect 378192 25712 378198 25764
rect 165246 25644 165252 25696
rect 165304 25684 165310 25696
rect 418154 25684 418160 25696
rect 165304 25656 418160 25684
rect 165304 25644 165310 25656
rect 418154 25644 418160 25656
rect 418212 25644 418218 25696
rect 171134 25576 171140 25628
rect 171192 25616 171198 25628
rect 509234 25616 509240 25628
rect 171192 25588 509240 25616
rect 171192 25576 171198 25588
rect 509234 25576 509240 25588
rect 509292 25576 509298 25628
rect 173710 25508 173716 25560
rect 173768 25548 173774 25560
rect 524414 25548 524420 25560
rect 173768 25520 524420 25548
rect 173768 25508 173774 25520
rect 524414 25508 524420 25520
rect 524472 25508 524478 25560
rect 154298 24284 154304 24336
rect 154356 24324 154362 24336
rect 282914 24324 282920 24336
rect 154356 24296 282920 24324
rect 154356 24284 154362 24296
rect 282914 24284 282920 24296
rect 282972 24284 282978 24336
rect 163958 24216 163964 24268
rect 164016 24256 164022 24268
rect 391934 24256 391940 24268
rect 164016 24228 391940 24256
rect 164016 24216 164022 24228
rect 391934 24216 391940 24228
rect 391992 24216 391998 24268
rect 172422 24148 172428 24200
rect 172480 24188 172486 24200
rect 513374 24188 513380 24200
rect 172480 24160 513380 24188
rect 172480 24148 172486 24160
rect 513374 24148 513380 24160
rect 513432 24148 513438 24200
rect 173618 24080 173624 24132
rect 173676 24120 173682 24132
rect 531406 24120 531412 24132
rect 173676 24092 531412 24120
rect 173676 24080 173682 24092
rect 531406 24080 531412 24092
rect 531464 24080 531470 24132
rect 157058 22992 157064 23044
rect 157116 23032 157122 23044
rect 310514 23032 310520 23044
rect 157116 23004 310520 23032
rect 157116 22992 157122 23004
rect 310514 22992 310520 23004
rect 310572 22992 310578 23044
rect 162854 22924 162860 22976
rect 162912 22964 162918 22976
rect 398926 22964 398932 22976
rect 162912 22936 398932 22964
rect 162912 22924 162918 22936
rect 398926 22924 398932 22936
rect 398984 22924 398990 22976
rect 166626 22856 166632 22908
rect 166684 22896 166690 22908
rect 440326 22896 440332 22908
rect 166684 22868 440332 22896
rect 166684 22856 166690 22868
rect 440326 22856 440332 22868
rect 440384 22856 440390 22908
rect 173802 22788 173808 22840
rect 173860 22828 173866 22840
rect 520274 22828 520280 22840
rect 173860 22800 520280 22828
rect 173860 22788 173866 22800
rect 520274 22788 520280 22800
rect 520332 22788 520338 22840
rect 175090 22720 175096 22772
rect 175148 22760 175154 22772
rect 538950 22760 538956 22772
rect 175148 22732 538956 22760
rect 175148 22720 175154 22732
rect 538950 22720 538956 22732
rect 539008 22720 539014 22772
rect 143718 21360 143724 21412
rect 143776 21400 143782 21412
rect 157978 21400 157984 21412
rect 143776 21372 157984 21400
rect 143776 21360 143782 21372
rect 157978 21360 157984 21372
rect 158036 21360 158042 21412
rect 158438 21360 158444 21412
rect 158496 21400 158502 21412
rect 329098 21400 329104 21412
rect 158496 21372 329104 21400
rect 158496 21360 158502 21372
rect 329098 21360 329104 21372
rect 329156 21360 329162 21412
rect 342898 21360 342904 21412
rect 342956 21400 342962 21412
rect 471974 21400 471980 21412
rect 342956 21372 471980 21400
rect 342956 21360 342962 21372
rect 471974 21360 471980 21372
rect 472032 21360 472038 21412
rect 153838 20136 153844 20188
rect 153896 20176 153902 20188
rect 280154 20176 280160 20188
rect 153896 20148 280160 20176
rect 153896 20136 153902 20148
rect 280154 20136 280160 20148
rect 280212 20136 280218 20188
rect 155218 20068 155224 20120
rect 155276 20108 155282 20120
rect 291194 20108 291200 20120
rect 155276 20080 291200 20108
rect 155276 20068 155282 20080
rect 291194 20068 291200 20080
rect 291252 20068 291258 20120
rect 155678 20000 155684 20052
rect 155736 20040 155742 20052
rect 287054 20040 287060 20052
rect 155736 20012 287060 20040
rect 155736 20000 155742 20012
rect 287054 20000 287060 20012
rect 287112 20000 287118 20052
rect 287698 20000 287704 20052
rect 287756 20040 287762 20052
rect 456886 20040 456892 20052
rect 287756 20012 456892 20040
rect 287756 20000 287762 20012
rect 456886 20000 456892 20012
rect 456944 20000 456950 20052
rect 161014 19932 161020 19984
rect 161072 19972 161078 19984
rect 357526 19972 357532 19984
rect 161072 19944 357532 19972
rect 161072 19932 161078 19944
rect 357526 19932 357532 19944
rect 357584 19932 357590 19984
rect 154022 18776 154028 18828
rect 154080 18816 154086 18828
rect 273254 18816 273260 18828
rect 154080 18788 273260 18816
rect 154080 18776 154086 18788
rect 273254 18776 273260 18788
rect 273312 18776 273318 18828
rect 166166 18708 166172 18760
rect 166224 18748 166230 18760
rect 431954 18748 431960 18760
rect 166224 18720 431960 18748
rect 166224 18708 166230 18720
rect 431954 18708 431960 18720
rect 432012 18708 432018 18760
rect 176286 18640 176292 18692
rect 176344 18680 176350 18692
rect 567194 18680 567200 18692
rect 176344 18652 567200 18680
rect 176344 18640 176350 18652
rect 567194 18640 567200 18652
rect 567252 18640 567258 18692
rect 177942 18572 177948 18624
rect 178000 18612 178006 18624
rect 571334 18612 571340 18624
rect 178000 18584 571340 18612
rect 178000 18572 178006 18584
rect 571334 18572 571340 18584
rect 571392 18572 571398 18624
rect 149882 17416 149888 17468
rect 149940 17456 149946 17468
rect 219434 17456 219440 17468
rect 149940 17428 219440 17456
rect 149940 17416 149946 17428
rect 219434 17416 219440 17428
rect 219492 17416 219498 17468
rect 168190 17348 168196 17400
rect 168248 17388 168254 17400
rect 445754 17388 445760 17400
rect 168248 17360 445760 17388
rect 168248 17348 168254 17360
rect 445754 17348 445760 17360
rect 445812 17348 445818 17400
rect 169662 17280 169668 17332
rect 169720 17320 169726 17332
rect 477494 17320 477500 17332
rect 169720 17292 477500 17320
rect 169720 17280 169726 17292
rect 477494 17280 477500 17292
rect 477552 17280 477558 17332
rect 177850 17212 177856 17264
rect 177908 17252 177914 17264
rect 570598 17252 570604 17264
rect 177908 17224 570604 17252
rect 177908 17212 177914 17224
rect 570598 17212 570604 17224
rect 570656 17212 570662 17264
rect 149698 16124 149704 16176
rect 149756 16164 149762 16176
rect 227530 16164 227536 16176
rect 149756 16136 227536 16164
rect 149756 16124 149762 16136
rect 227530 16124 227536 16136
rect 227588 16124 227594 16176
rect 161106 16056 161112 16108
rect 161164 16096 161170 16108
rect 361114 16096 361120 16108
rect 161164 16068 361120 16096
rect 161164 16056 161170 16068
rect 361114 16056 361120 16068
rect 361172 16056 361178 16108
rect 161198 15988 161204 16040
rect 161256 16028 161262 16040
rect 364610 16028 364616 16040
rect 161256 16000 364616 16028
rect 161256 15988 161262 16000
rect 364610 15988 364616 16000
rect 364668 15988 364674 16040
rect 165338 15920 165344 15972
rect 165396 15960 165402 15972
rect 420914 15960 420920 15972
rect 165396 15932 420920 15960
rect 165396 15920 165402 15932
rect 420914 15920 420920 15932
rect 420972 15920 420978 15972
rect 176378 15852 176384 15904
rect 176436 15892 176442 15904
rect 560386 15892 560392 15904
rect 176436 15864 560392 15892
rect 176436 15852 176442 15864
rect 560386 15852 560392 15864
rect 560444 15852 560450 15904
rect 155770 14696 155776 14748
rect 155828 14736 155834 14748
rect 293218 14736 293224 14748
rect 155828 14708 293224 14736
rect 155828 14696 155834 14708
rect 293218 14696 293224 14708
rect 293276 14696 293282 14748
rect 157150 14628 157156 14680
rect 157208 14668 157214 14680
rect 314654 14668 314660 14680
rect 157208 14640 314660 14668
rect 157208 14628 157214 14640
rect 314654 14628 314660 14640
rect 314712 14628 314718 14680
rect 162670 14560 162676 14612
rect 162728 14600 162734 14612
rect 385954 14600 385960 14612
rect 162728 14572 385960 14600
rect 162728 14560 162734 14572
rect 385954 14560 385960 14572
rect 386012 14560 386018 14612
rect 164050 14492 164056 14544
rect 164108 14532 164114 14544
rect 404354 14532 404360 14544
rect 164108 14504 404360 14532
rect 164108 14492 164114 14504
rect 404354 14492 404360 14504
rect 404412 14492 404418 14544
rect 30098 14424 30104 14476
rect 30156 14464 30162 14476
rect 133874 14464 133880 14476
rect 30156 14436 133880 14464
rect 30156 14424 30162 14436
rect 133874 14424 133880 14436
rect 133932 14424 133938 14476
rect 170950 14424 170956 14476
rect 171008 14464 171014 14476
rect 493042 14464 493048 14476
rect 171008 14436 493048 14464
rect 171008 14424 171014 14436
rect 493042 14424 493048 14436
rect 493100 14424 493106 14476
rect 153930 13336 153936 13388
rect 153988 13376 153994 13388
rect 272426 13376 272432 13388
rect 153988 13348 272432 13376
rect 153988 13336 153994 13348
rect 272426 13336 272432 13348
rect 272484 13336 272490 13388
rect 157242 13268 157248 13320
rect 157300 13308 157306 13320
rect 307938 13308 307944 13320
rect 157300 13280 307944 13308
rect 157300 13268 157306 13280
rect 307938 13268 307944 13280
rect 307996 13268 308002 13320
rect 162578 13200 162584 13252
rect 162636 13240 162642 13252
rect 382366 13240 382372 13252
rect 162636 13212 382372 13240
rect 162636 13200 162642 13212
rect 382366 13200 382372 13212
rect 382424 13200 382430 13252
rect 162486 13132 162492 13184
rect 162544 13172 162550 13184
rect 386690 13172 386696 13184
rect 162544 13144 386696 13172
rect 162544 13132 162550 13144
rect 386690 13132 386696 13144
rect 386748 13132 386754 13184
rect 144178 13064 144184 13116
rect 144236 13104 144242 13116
rect 155402 13104 155408 13116
rect 144236 13076 155408 13104
rect 144236 13064 144242 13076
rect 155402 13064 155408 13076
rect 155460 13064 155466 13116
rect 170858 13064 170864 13116
rect 170916 13104 170922 13116
rect 486326 13104 486332 13116
rect 170916 13076 486332 13104
rect 170916 13064 170922 13076
rect 486326 13064 486332 13076
rect 486384 13064 486390 13116
rect 486418 13064 486424 13116
rect 486476 13104 486482 13116
rect 581730 13104 581736 13116
rect 486476 13076 581736 13104
rect 486476 13064 486482 13076
rect 581730 13064 581736 13076
rect 581788 13064 581794 13116
rect 151170 11976 151176 12028
rect 151228 12016 151234 12028
rect 241698 12016 241704 12028
rect 151228 11988 241704 12016
rect 151228 11976 151234 11988
rect 241698 11976 241704 11988
rect 241756 11976 241762 12028
rect 157334 11908 157340 11960
rect 157392 11948 157398 11960
rect 328730 11948 328736 11960
rect 157392 11920 328736 11948
rect 157392 11908 157398 11920
rect 328730 11908 328736 11920
rect 328788 11908 328794 11960
rect 162762 11840 162768 11892
rect 162820 11880 162826 11892
rect 379514 11880 379520 11892
rect 162820 11852 379520 11880
rect 162820 11840 162826 11852
rect 379514 11840 379520 11852
rect 379572 11840 379578 11892
rect 165430 11772 165436 11824
rect 165488 11812 165494 11824
rect 417418 11812 417424 11824
rect 165488 11784 417424 11812
rect 165488 11772 165494 11784
rect 417418 11772 417424 11784
rect 417476 11772 417482 11824
rect 174078 11704 174084 11756
rect 174136 11744 174142 11756
rect 541986 11744 541992 11756
rect 174136 11716 541992 11744
rect 174136 11704 174142 11716
rect 541986 11704 541992 11716
rect 542044 11704 542050 11756
rect 209958 11636 209964 11688
rect 210016 11676 210022 11688
rect 210970 11676 210976 11688
rect 210016 11648 210976 11676
rect 210016 11636 210022 11648
rect 210970 11636 210976 11648
rect 211028 11636 211034 11688
rect 234614 11636 234620 11688
rect 234672 11676 234678 11688
rect 235810 11676 235816 11688
rect 234672 11648 235816 11676
rect 234672 11636 234678 11648
rect 235810 11636 235816 11648
rect 235868 11636 235874 11688
rect 259454 11636 259460 11688
rect 259512 11676 259518 11688
rect 260650 11676 260656 11688
rect 259512 11648 260656 11676
rect 259512 11636 259518 11648
rect 260650 11636 260656 11648
rect 260708 11636 260714 11688
rect 151262 10548 151268 10600
rect 151320 10588 151326 10600
rect 234614 10588 234620 10600
rect 151320 10560 234620 10588
rect 151320 10548 151326 10560
rect 234614 10548 234620 10560
rect 234672 10548 234678 10600
rect 158530 10480 158536 10532
rect 158588 10520 158594 10532
rect 336274 10520 336280 10532
rect 158588 10492 336280 10520
rect 158588 10480 158594 10492
rect 336274 10480 336280 10492
rect 336332 10480 336338 10532
rect 160094 10412 160100 10464
rect 160152 10452 160158 10464
rect 372890 10452 372896 10464
rect 160152 10424 372896 10452
rect 160152 10412 160158 10424
rect 372890 10412 372896 10424
rect 372948 10412 372954 10464
rect 166718 10344 166724 10396
rect 166776 10384 166782 10396
rect 432046 10384 432052 10396
rect 166776 10356 432052 10384
rect 166776 10344 166782 10356
rect 432046 10344 432052 10356
rect 432104 10344 432110 10396
rect 87506 10276 87512 10328
rect 87564 10316 87570 10328
rect 138106 10316 138112 10328
rect 87564 10288 138112 10316
rect 87564 10276 87570 10288
rect 138106 10276 138112 10288
rect 138164 10276 138170 10328
rect 173986 10276 173992 10328
rect 174044 10316 174050 10328
rect 548610 10316 548616 10328
rect 174044 10288 548616 10316
rect 174044 10276 174050 10288
rect 548610 10276 548616 10288
rect 548668 10276 548674 10328
rect 155862 9120 155868 9172
rect 155920 9160 155926 9172
rect 301958 9160 301964 9172
rect 155920 9132 301964 9160
rect 155920 9120 155926 9132
rect 301958 9120 301964 9132
rect 302016 9120 302022 9172
rect 158622 9052 158628 9104
rect 158680 9092 158686 9104
rect 325602 9092 325608 9104
rect 158680 9064 325608 9092
rect 158680 9052 158686 9064
rect 325602 9052 325608 9064
rect 325660 9052 325666 9104
rect 165522 8984 165528 9036
rect 165580 9024 165586 9036
rect 414290 9024 414296 9036
rect 165580 8996 414296 9024
rect 165580 8984 165586 8996
rect 414290 8984 414296 8996
rect 414348 8984 414354 9036
rect 143626 8916 143632 8968
rect 143684 8956 143690 8968
rect 157794 8956 157800 8968
rect 143684 8928 157800 8956
rect 143684 8916 143690 8928
rect 157794 8916 157800 8928
rect 157852 8916 157858 8968
rect 176470 8916 176476 8968
rect 176528 8956 176534 8968
rect 556154 8956 556160 8968
rect 176528 8928 556160 8956
rect 176528 8916 176534 8928
rect 556154 8916 556160 8928
rect 556212 8916 556218 8968
rect 160002 7828 160008 7880
rect 160060 7868 160066 7880
rect 343358 7868 343364 7880
rect 160060 7840 343364 7868
rect 160060 7828 160066 7840
rect 343358 7828 343364 7840
rect 343416 7828 343422 7880
rect 161382 7760 161388 7812
rect 161440 7800 161446 7812
rect 365806 7800 365812 7812
rect 161440 7772 365812 7800
rect 161440 7760 161446 7772
rect 365806 7760 365812 7772
rect 365864 7760 365870 7812
rect 166902 7692 166908 7744
rect 166960 7732 166966 7744
rect 435542 7732 435548 7744
rect 166960 7704 435548 7732
rect 166960 7692 166966 7704
rect 435542 7692 435548 7704
rect 435600 7692 435606 7744
rect 166810 7624 166816 7676
rect 166868 7664 166874 7676
rect 442626 7664 442632 7676
rect 166868 7636 442632 7664
rect 166868 7624 166874 7636
rect 442626 7624 442632 7636
rect 442684 7624 442690 7676
rect 54938 7556 54944 7608
rect 54996 7596 55002 7608
rect 135530 7596 135536 7608
rect 54996 7568 135536 7596
rect 54996 7556 55002 7568
rect 135530 7556 135536 7568
rect 135588 7556 135594 7608
rect 173894 7556 173900 7608
rect 173952 7596 173958 7608
rect 538398 7596 538404 7608
rect 173952 7568 538404 7596
rect 173952 7556 173958 7568
rect 538398 7556 538404 7568
rect 538456 7556 538462 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 17218 6848 17224 6860
rect 3476 6820 17224 6848
rect 3476 6808 3482 6820
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 152550 6536 152556 6588
rect 152608 6576 152614 6588
rect 252370 6576 252376 6588
rect 152608 6548 252376 6576
rect 152608 6536 152614 6548
rect 252370 6536 252376 6548
rect 252428 6536 252434 6588
rect 158714 6468 158720 6520
rect 158772 6508 158778 6520
rect 350442 6508 350448 6520
rect 158772 6480 350448 6508
rect 158772 6468 158778 6480
rect 350442 6468 350448 6480
rect 350500 6468 350506 6520
rect 180058 6400 180064 6452
rect 180116 6440 180122 6452
rect 436738 6440 436744 6452
rect 180116 6412 436744 6440
rect 180116 6400 180122 6412
rect 436738 6400 436744 6412
rect 436796 6400 436802 6452
rect 182082 6332 182088 6384
rect 182140 6372 182146 6384
rect 443822 6372 443828 6384
rect 182140 6344 443828 6372
rect 182140 6332 182146 6344
rect 443822 6332 443828 6344
rect 443880 6332 443886 6384
rect 179138 6264 179144 6316
rect 179196 6304 179202 6316
rect 450906 6304 450912 6316
rect 179196 6276 450912 6304
rect 179196 6264 179202 6276
rect 450906 6264 450912 6276
rect 450964 6264 450970 6316
rect 168282 6196 168288 6248
rect 168340 6236 168346 6248
rect 453206 6236 453212 6248
rect 168340 6208 453212 6236
rect 168340 6196 168346 6208
rect 453206 6196 453212 6208
rect 453264 6196 453270 6248
rect 453298 6196 453304 6248
rect 453356 6236 453362 6248
rect 479334 6236 479340 6248
rect 453356 6208 479340 6236
rect 453356 6196 453362 6208
rect 479334 6196 479340 6208
rect 479392 6196 479398 6248
rect 28902 6128 28908 6180
rect 28960 6168 28966 6180
rect 134058 6168 134064 6180
rect 28960 6140 134064 6168
rect 28960 6128 28966 6140
rect 134058 6128 134064 6140
rect 134116 6128 134122 6180
rect 176562 6128 176568 6180
rect 176620 6168 176626 6180
rect 563238 6168 563244 6180
rect 176620 6140 563244 6168
rect 176620 6128 176626 6140
rect 563238 6128 563244 6140
rect 563296 6128 563302 6180
rect 143534 5652 143540 5704
rect 143592 5692 143598 5704
rect 144730 5692 144736 5704
rect 143592 5664 144736 5692
rect 143592 5652 143598 5664
rect 144730 5652 144736 5664
rect 144788 5652 144794 5704
rect 142798 5516 142804 5568
rect 142856 5556 142862 5568
rect 143534 5556 143540 5568
rect 142856 5528 143540 5556
rect 142856 5516 142862 5528
rect 143534 5516 143540 5528
rect 143592 5516 143598 5568
rect 151078 5040 151084 5092
rect 151136 5080 151142 5092
rect 245194 5080 245200 5092
rect 151136 5052 245200 5080
rect 151136 5040 151142 5052
rect 245194 5040 245200 5052
rect 245252 5040 245258 5092
rect 161198 4972 161204 5024
rect 161256 5012 161262 5024
rect 371694 5012 371700 5024
rect 161256 4984 371700 5012
rect 161256 4972 161262 4984
rect 371694 4972 371700 4984
rect 371752 4972 371758 5024
rect 164142 4904 164148 4956
rect 164200 4944 164206 4956
rect 397730 4944 397736 4956
rect 164200 4916 397736 4944
rect 164200 4904 164206 4916
rect 397730 4904 397736 4916
rect 397788 4904 397794 4956
rect 171042 4836 171048 4888
rect 171100 4876 171106 4888
rect 482830 4876 482836 4888
rect 171100 4848 482836 4876
rect 171100 4836 171106 4848
rect 482830 4836 482836 4848
rect 482888 4836 482894 4888
rect 175182 4768 175188 4820
rect 175240 4808 175246 4820
rect 545482 4808 545488 4820
rect 175240 4780 545488 4808
rect 175240 4768 175246 4780
rect 545482 4768 545488 4780
rect 545540 4768 545546 4820
rect 566 4088 572 4140
rect 624 4128 630 4140
rect 7558 4128 7564 4140
rect 624 4100 7564 4128
rect 624 4088 630 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 17310 4128 17316 4140
rect 15988 4100 17316 4128
rect 15988 4088 15994 4100
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 73798 4088 73804 4140
rect 73856 4128 73862 4140
rect 75178 4128 75184 4140
rect 73856 4100 75184 4128
rect 73856 4088 73862 4100
rect 75178 4088 75184 4100
rect 75236 4088 75242 4140
rect 181990 4088 181996 4140
rect 182048 4128 182054 4140
rect 187418 4128 187424 4140
rect 182048 4100 187424 4128
rect 182048 4088 182054 4100
rect 187418 4088 187424 4100
rect 187476 4088 187482 4140
rect 188338 4088 188344 4140
rect 188396 4128 188402 4140
rect 193858 4128 193864 4140
rect 188396 4100 193864 4128
rect 188396 4088 188402 4100
rect 193858 4088 193864 4100
rect 193916 4088 193922 4140
rect 194042 4088 194048 4140
rect 194100 4128 194106 4140
rect 195606 4128 195612 4140
rect 194100 4100 195612 4128
rect 194100 4088 194106 4100
rect 195606 4088 195612 4100
rect 195664 4088 195670 4140
rect 196618 4088 196624 4140
rect 196676 4128 196682 4140
rect 203886 4128 203892 4140
rect 196676 4100 203892 4128
rect 196676 4088 196682 4100
rect 203886 4088 203892 4100
rect 203944 4088 203950 4140
rect 203978 4088 203984 4140
rect 204036 4128 204042 4140
rect 247586 4128 247592 4140
rect 204036 4100 247592 4128
rect 204036 4088 204042 4100
rect 247586 4088 247592 4100
rect 247644 4088 247650 4140
rect 247678 4088 247684 4140
rect 247736 4128 247742 4140
rect 254670 4128 254676 4140
rect 247736 4100 254676 4128
rect 247736 4088 247742 4100
rect 254670 4088 254676 4100
rect 254728 4088 254734 4140
rect 257338 4088 257344 4140
rect 257396 4128 257402 4140
rect 258258 4128 258264 4140
rect 257396 4100 258264 4128
rect 257396 4088 257402 4100
rect 258258 4088 258264 4100
rect 258316 4088 258322 4140
rect 261478 4088 261484 4140
rect 261536 4128 261542 4140
rect 262950 4128 262956 4140
rect 261536 4100 262956 4128
rect 261536 4088 261542 4100
rect 262950 4088 262956 4100
rect 263008 4088 263014 4140
rect 283558 4088 283564 4140
rect 283616 4128 283622 4140
rect 298462 4128 298468 4140
rect 283616 4100 298468 4128
rect 283616 4088 283622 4100
rect 298462 4088 298468 4100
rect 298520 4088 298526 4140
rect 450538 4088 450544 4140
rect 450596 4128 450602 4140
rect 452102 4128 452108 4140
rect 450596 4100 452108 4128
rect 450596 4088 450602 4100
rect 452102 4088 452108 4100
rect 452160 4088 452166 4140
rect 563698 4088 563704 4140
rect 563756 4128 563762 4140
rect 569126 4128 569132 4140
rect 563756 4100 569132 4128
rect 563756 4088 563762 4100
rect 569126 4088 569132 4100
rect 569184 4088 569190 4140
rect 6454 4020 6460 4072
rect 6512 4060 6518 4072
rect 7650 4060 7656 4072
rect 6512 4032 7656 4060
rect 6512 4020 6518 4032
rect 7650 4020 7656 4032
rect 7708 4020 7714 4072
rect 102226 4020 102232 4072
rect 102284 4060 102290 4072
rect 113266 4060 113272 4072
rect 102284 4032 113272 4060
rect 102284 4020 102290 4032
rect 113266 4020 113272 4032
rect 113324 4020 113330 4072
rect 119890 4020 119896 4072
rect 119948 4060 119954 4072
rect 122098 4060 122104 4072
rect 119948 4032 122104 4060
rect 119948 4020 119954 4032
rect 122098 4020 122104 4032
rect 122156 4020 122162 4072
rect 146846 4020 146852 4072
rect 146904 4060 146910 4072
rect 153010 4060 153016 4072
rect 146904 4032 153016 4060
rect 146904 4020 146910 4032
rect 153010 4020 153016 4032
rect 153068 4020 153074 4072
rect 182818 4020 182824 4072
rect 182876 4060 182882 4072
rect 212166 4060 212172 4072
rect 182876 4032 212172 4060
rect 182876 4020 182882 4032
rect 212166 4020 212172 4032
rect 212224 4020 212230 4072
rect 224218 4020 224224 4072
rect 224276 4060 224282 4072
rect 284294 4060 284300 4072
rect 224276 4032 284300 4060
rect 224276 4020 224282 4032
rect 284294 4020 284300 4032
rect 284352 4020 284358 4072
rect 299566 4020 299572 4072
rect 299624 4060 299630 4072
rect 300762 4060 300768 4072
rect 299624 4032 300768 4060
rect 299624 4020 299630 4032
rect 300762 4020 300768 4032
rect 300820 4020 300826 4072
rect 311158 4020 311164 4072
rect 311216 4060 311222 4072
rect 312630 4060 312636 4072
rect 311216 4032 312636 4060
rect 311216 4020 311222 4032
rect 312630 4020 312636 4032
rect 312688 4020 312694 4072
rect 85666 3952 85672 4004
rect 85724 3992 85730 4004
rect 88978 3992 88984 4004
rect 85724 3964 88984 3992
rect 85724 3952 85730 3964
rect 88978 3952 88984 3964
rect 89036 3952 89042 4004
rect 111610 3952 111616 4004
rect 111668 3992 111674 4004
rect 129826 3992 129832 4004
rect 111668 3964 129832 3992
rect 111668 3952 111674 3964
rect 129826 3952 129832 3964
rect 129884 3952 129890 4004
rect 179322 3952 179328 4004
rect 179380 3992 179386 4004
rect 394234 3992 394240 4004
rect 179380 3964 394240 3992
rect 179380 3952 179386 3964
rect 394234 3952 394240 3964
rect 394292 3952 394298 4004
rect 83274 3884 83280 3936
rect 83332 3924 83338 3936
rect 127158 3924 127164 3936
rect 83332 3896 127164 3924
rect 83332 3884 83338 3896
rect 127158 3884 127164 3896
rect 127216 3884 127222 3936
rect 179230 3884 179236 3936
rect 179288 3924 179294 3936
rect 401318 3924 401324 3936
rect 179288 3896 401324 3924
rect 179288 3884 179294 3896
rect 401318 3884 401324 3896
rect 401376 3884 401382 3936
rect 65518 3816 65524 3868
rect 65576 3856 65582 3868
rect 65576 3828 71176 3856
rect 65576 3816 65582 3828
rect 69106 3748 69112 3800
rect 69164 3788 69170 3800
rect 71038 3788 71044 3800
rect 69164 3760 71044 3788
rect 69164 3748 69170 3760
rect 71038 3748 71044 3760
rect 71096 3748 71102 3800
rect 71148 3788 71176 3828
rect 72602 3816 72608 3868
rect 72660 3856 72666 3868
rect 130010 3856 130016 3868
rect 72660 3828 130016 3856
rect 72660 3816 72666 3828
rect 130010 3816 130016 3828
rect 130068 3816 130074 3868
rect 130930 3816 130936 3868
rect 130988 3856 130994 3868
rect 150618 3856 150624 3868
rect 130988 3828 150624 3856
rect 130988 3816 130994 3828
rect 150618 3816 150624 3828
rect 150676 3816 150682 3868
rect 152642 3816 152648 3868
rect 152700 3856 152706 3868
rect 164878 3856 164884 3868
rect 152700 3828 164884 3856
rect 152700 3816 152706 3828
rect 164878 3816 164884 3828
rect 164936 3816 164942 3868
rect 178954 3816 178960 3868
rect 179012 3856 179018 3868
rect 408402 3856 408408 3868
rect 179012 3828 408408 3856
rect 179012 3816 179018 3828
rect 408402 3816 408408 3828
rect 408460 3816 408466 3868
rect 410518 3816 410524 3868
rect 410576 3856 410582 3868
rect 411898 3856 411904 3868
rect 410576 3828 411904 3856
rect 410576 3816 410582 3828
rect 411898 3816 411904 3828
rect 411956 3816 411962 3868
rect 131298 3788 131304 3800
rect 71148 3760 131304 3788
rect 131298 3748 131304 3760
rect 131356 3748 131362 3800
rect 146938 3748 146944 3800
rect 146996 3788 147002 3800
rect 146996 3760 149652 3788
rect 146996 3748 147002 3760
rect 39574 3680 39580 3732
rect 39632 3720 39638 3732
rect 131390 3720 131396 3732
rect 39632 3692 131396 3720
rect 39632 3680 39638 3692
rect 131390 3680 131396 3692
rect 131448 3680 131454 3732
rect 137646 3680 137652 3732
rect 137704 3720 137710 3732
rect 138658 3720 138664 3732
rect 137704 3692 138664 3720
rect 137704 3680 137710 3692
rect 138658 3680 138664 3692
rect 138716 3680 138722 3732
rect 147030 3680 147036 3732
rect 147088 3720 147094 3732
rect 149514 3720 149520 3732
rect 147088 3692 149520 3720
rect 147088 3680 147094 3692
rect 149514 3680 149520 3692
rect 149572 3680 149578 3732
rect 149624 3720 149652 3760
rect 149790 3748 149796 3800
rect 149848 3788 149854 3800
rect 156598 3788 156604 3800
rect 149848 3760 156604 3788
rect 149848 3748 149854 3760
rect 156598 3748 156604 3760
rect 156656 3748 156662 3800
rect 156782 3748 156788 3800
rect 156840 3788 156846 3800
rect 170766 3788 170772 3800
rect 156840 3760 170772 3788
rect 156840 3748 156846 3760
rect 170766 3748 170772 3760
rect 170824 3748 170830 3800
rect 184106 3748 184112 3800
rect 184164 3788 184170 3800
rect 415486 3788 415492 3800
rect 184164 3760 415492 3788
rect 184164 3748 184170 3760
rect 415486 3748 415492 3760
rect 415544 3748 415550 3800
rect 163682 3720 163688 3732
rect 149624 3692 163688 3720
rect 163682 3680 163688 3692
rect 163740 3680 163746 3732
rect 180610 3680 180616 3732
rect 180668 3720 180674 3732
rect 422570 3720 422576 3732
rect 180668 3692 422576 3720
rect 180668 3680 180674 3692
rect 422570 3680 422576 3692
rect 422628 3680 422634 3732
rect 489178 3680 489184 3732
rect 489236 3720 489242 3732
rect 491110 3720 491116 3732
rect 489236 3692 491116 3720
rect 489236 3680 489242 3692
rect 491110 3680 491116 3692
rect 491168 3680 491174 3732
rect 7650 3612 7656 3664
rect 7708 3652 7714 3664
rect 7708 3624 16574 3652
rect 7708 3612 7714 3624
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 13078 3584 13084 3596
rect 11204 3556 13084 3584
rect 11204 3544 11210 3556
rect 13078 3544 13084 3556
rect 13136 3544 13142 3596
rect 16546 3584 16574 3624
rect 21818 3612 21824 3664
rect 21876 3652 21882 3664
rect 124214 3652 124220 3664
rect 21876 3624 124220 3652
rect 21876 3612 21882 3624
rect 124214 3612 124220 3624
rect 124272 3612 124278 3664
rect 124674 3612 124680 3664
rect 124732 3652 124738 3664
rect 129918 3652 129924 3664
rect 124732 3624 129924 3652
rect 124732 3612 124738 3624
rect 129918 3612 129924 3624
rect 129976 3612 129982 3664
rect 131022 3612 131028 3664
rect 131080 3652 131086 3664
rect 162486 3652 162492 3664
rect 131080 3624 162492 3652
rect 131080 3612 131086 3624
rect 162486 3612 162492 3624
rect 162544 3612 162550 3664
rect 180702 3612 180708 3664
rect 180760 3652 180766 3664
rect 429654 3652 429660 3664
rect 180760 3624 429660 3652
rect 180760 3612 180766 3624
rect 429654 3612 429660 3624
rect 429712 3612 429718 3664
rect 431954 3612 431960 3664
rect 432012 3652 432018 3664
rect 433242 3652 433248 3664
rect 432012 3624 433248 3652
rect 432012 3612 432018 3624
rect 433242 3612 433248 3624
rect 433300 3612 433306 3664
rect 454678 3612 454684 3664
rect 454736 3652 454742 3664
rect 497090 3652 497096 3664
rect 454736 3624 497096 3652
rect 454736 3612 454742 3624
rect 497090 3612 497096 3624
rect 497148 3612 497154 3664
rect 127066 3584 127072 3596
rect 16546 3556 127072 3584
rect 127066 3544 127072 3556
rect 127124 3544 127130 3596
rect 128262 3544 128268 3596
rect 128320 3584 128326 3596
rect 166074 3584 166080 3596
rect 128320 3556 166080 3584
rect 128320 3544 128326 3556
rect 166074 3544 166080 3556
rect 166132 3544 166138 3596
rect 176654 3544 176660 3596
rect 176712 3584 176718 3596
rect 179506 3584 179512 3596
rect 176712 3556 179512 3584
rect 176712 3544 176718 3556
rect 179506 3544 179512 3556
rect 179564 3544 179570 3596
rect 185578 3544 185584 3596
rect 185636 3584 185642 3596
rect 187326 3584 187332 3596
rect 185636 3556 187332 3584
rect 185636 3544 185642 3556
rect 187326 3544 187332 3556
rect 187384 3544 187390 3596
rect 187418 3544 187424 3596
rect 187476 3584 187482 3596
rect 461578 3584 461584 3596
rect 187476 3556 461584 3584
rect 187476 3544 187482 3556
rect 461578 3544 461584 3556
rect 461636 3544 461642 3596
rect 525058 3544 525064 3596
rect 525116 3584 525122 3596
rect 527818 3584 527824 3596
rect 525116 3556 527824 3584
rect 525116 3544 525122 3556
rect 527818 3544 527824 3556
rect 527876 3544 527882 3596
rect 574738 3544 574744 3596
rect 574796 3584 574802 3596
rect 576302 3584 576308 3596
rect 574796 3556 576308 3584
rect 574796 3544 574802 3556
rect 576302 3544 576308 3556
rect 576360 3544 576366 3596
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 4798 3516 4804 3528
rect 4120 3488 4804 3516
rect 4120 3476 4126 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 5316 3488 122972 3516
rect 5316 3476 5322 3488
rect 17034 3408 17040 3460
rect 17092 3448 17098 3460
rect 18598 3448 18604 3460
rect 17092 3420 18604 3448
rect 17092 3408 17098 3420
rect 18598 3408 18604 3420
rect 18656 3408 18662 3460
rect 20622 3408 20628 3460
rect 20680 3448 20686 3460
rect 20680 3420 122834 3448
rect 20680 3408 20686 3420
rect 33594 3340 33600 3392
rect 33652 3380 33658 3392
rect 35158 3380 35164 3392
rect 33652 3352 35164 3380
rect 33652 3340 33658 3352
rect 35158 3340 35164 3352
rect 35216 3340 35222 3392
rect 38378 3340 38384 3392
rect 38436 3380 38442 3392
rect 39298 3380 39304 3392
rect 38436 3352 39304 3380
rect 38436 3340 38442 3352
rect 39298 3340 39304 3352
rect 39356 3340 39362 3392
rect 52454 3340 52460 3392
rect 52512 3380 52518 3392
rect 53374 3380 53380 3392
rect 52512 3352 53380 3380
rect 52512 3340 52518 3352
rect 53374 3340 53380 3352
rect 53432 3340 53438 3392
rect 56042 3340 56048 3392
rect 56100 3380 56106 3392
rect 57238 3380 57244 3392
rect 56100 3352 57244 3380
rect 56100 3340 56106 3352
rect 57238 3340 57244 3352
rect 57296 3340 57302 3392
rect 91554 3340 91560 3392
rect 91612 3380 91618 3392
rect 93118 3380 93124 3392
rect 91612 3352 93124 3380
rect 91612 3340 91618 3352
rect 93118 3340 93124 3352
rect 93176 3340 93182 3392
rect 102134 3340 102140 3392
rect 102192 3380 102198 3392
rect 103330 3380 103336 3392
rect 102192 3352 103336 3380
rect 102192 3340 102198 3352
rect 103330 3340 103336 3352
rect 103388 3340 103394 3392
rect 105722 3340 105728 3392
rect 105780 3380 105786 3392
rect 106918 3380 106924 3392
rect 105780 3352 106924 3380
rect 105780 3340 105786 3352
rect 106918 3340 106924 3352
rect 106976 3340 106982 3392
rect 109310 3340 109316 3392
rect 109368 3380 109374 3392
rect 111242 3380 111248 3392
rect 109368 3352 111248 3380
rect 109368 3340 109374 3352
rect 111242 3340 111248 3352
rect 111300 3340 111306 3392
rect 51350 3272 51356 3324
rect 51408 3312 51414 3324
rect 54478 3312 54484 3324
rect 51408 3284 54484 3312
rect 51408 3272 51414 3284
rect 54478 3272 54484 3284
rect 54536 3272 54542 3324
rect 101030 3272 101036 3324
rect 101088 3312 101094 3324
rect 102778 3312 102784 3324
rect 101088 3284 102784 3312
rect 101088 3272 101094 3284
rect 102778 3272 102784 3284
rect 102836 3272 102842 3324
rect 93946 3136 93952 3188
rect 94004 3176 94010 3188
rect 95970 3176 95976 3188
rect 94004 3148 95976 3176
rect 94004 3136 94010 3148
rect 95970 3136 95976 3148
rect 96028 3136 96034 3188
rect 122806 3176 122834 3420
rect 122944 3380 122972 3488
rect 126974 3476 126980 3528
rect 127032 3516 127038 3528
rect 128170 3516 128176 3528
rect 127032 3488 128176 3516
rect 127032 3476 127038 3488
rect 128170 3476 128176 3488
rect 128228 3476 128234 3528
rect 140038 3476 140044 3528
rect 140096 3516 140102 3528
rect 141510 3516 141516 3528
rect 140096 3488 141516 3516
rect 140096 3476 140102 3488
rect 141510 3476 141516 3488
rect 141568 3476 141574 3528
rect 157978 3476 157984 3528
rect 158036 3516 158042 3528
rect 158898 3516 158904 3528
rect 158036 3488 158904 3516
rect 158036 3476 158042 3488
rect 158898 3476 158904 3488
rect 158956 3476 158962 3528
rect 171962 3516 171968 3528
rect 159100 3488 171968 3516
rect 134150 3408 134156 3460
rect 134208 3448 134214 3460
rect 140130 3448 140136 3460
rect 134208 3420 140136 3448
rect 134208 3408 134214 3420
rect 140130 3408 140136 3420
rect 140188 3408 140194 3460
rect 147214 3408 147220 3460
rect 147272 3448 147278 3460
rect 148318 3448 148324 3460
rect 147272 3420 148324 3448
rect 147272 3408 147278 3420
rect 148318 3408 148324 3420
rect 148376 3408 148382 3460
rect 131574 3380 131580 3392
rect 122944 3352 131580 3380
rect 131574 3340 131580 3352
rect 131632 3340 131638 3392
rect 152458 3340 152464 3392
rect 152516 3380 152522 3392
rect 159100 3380 159128 3488
rect 171962 3476 171968 3488
rect 172020 3476 172026 3528
rect 173250 3476 173256 3528
rect 173308 3516 173314 3528
rect 177850 3516 177856 3528
rect 173308 3488 177856 3516
rect 173308 3476 173314 3488
rect 177850 3476 177856 3488
rect 177908 3476 177914 3528
rect 178678 3476 178684 3528
rect 178736 3516 178742 3528
rect 190822 3516 190828 3528
rect 178736 3488 190828 3516
rect 178736 3476 178742 3488
rect 190822 3476 190828 3488
rect 190880 3476 190886 3528
rect 193858 3476 193864 3528
rect 193916 3516 193922 3528
rect 196802 3516 196808 3528
rect 193916 3488 196808 3516
rect 193916 3476 193922 3488
rect 196802 3476 196808 3488
rect 196860 3476 196866 3528
rect 197998 3476 198004 3528
rect 198056 3516 198062 3528
rect 203978 3516 203984 3528
rect 198056 3488 203984 3516
rect 198056 3476 198062 3488
rect 203978 3476 203984 3488
rect 204036 3476 204042 3528
rect 204180 3488 470594 3516
rect 167638 3408 167644 3460
rect 167696 3448 167702 3460
rect 168374 3448 168380 3460
rect 167696 3420 168380 3448
rect 167696 3408 167702 3420
rect 168374 3408 168380 3420
rect 168432 3408 168438 3460
rect 171778 3408 171784 3460
rect 171836 3448 171842 3460
rect 173158 3448 173164 3460
rect 171836 3420 173164 3448
rect 171836 3408 171842 3420
rect 173158 3408 173164 3420
rect 173216 3408 173222 3460
rect 179046 3408 179052 3460
rect 179104 3448 179110 3460
rect 198090 3448 198096 3460
rect 179104 3420 198096 3448
rect 179104 3408 179110 3420
rect 198090 3408 198096 3420
rect 198148 3408 198154 3460
rect 175458 3380 175464 3392
rect 152516 3352 159128 3380
rect 161446 3352 175464 3380
rect 152516 3340 152522 3352
rect 126974 3272 126980 3324
rect 127032 3312 127038 3324
rect 128446 3312 128452 3324
rect 127032 3284 128452 3312
rect 127032 3272 127038 3284
rect 128446 3272 128452 3284
rect 128504 3272 128510 3324
rect 148410 3272 148416 3324
rect 148468 3312 148474 3324
rect 161446 3312 161474 3352
rect 175458 3340 175464 3352
rect 175516 3340 175522 3392
rect 184290 3340 184296 3392
rect 184348 3380 184354 3392
rect 189718 3380 189724 3392
rect 184348 3352 189724 3380
rect 184348 3340 184354 3352
rect 189718 3340 189724 3352
rect 189776 3340 189782 3392
rect 189810 3340 189816 3392
rect 189868 3380 189874 3392
rect 193214 3380 193220 3392
rect 189868 3352 193220 3380
rect 189868 3340 189874 3352
rect 193214 3340 193220 3352
rect 193272 3340 193278 3392
rect 204180 3380 204208 3488
rect 465166 3448 465172 3460
rect 198016 3352 204208 3380
rect 205606 3420 465172 3448
rect 148468 3284 161474 3312
rect 148468 3272 148474 3284
rect 193122 3272 193128 3324
rect 193180 3312 193186 3324
rect 198016 3312 198044 3352
rect 193180 3284 198044 3312
rect 193180 3272 193186 3284
rect 198090 3272 198096 3324
rect 198148 3312 198154 3324
rect 205606 3312 205634 3420
rect 465166 3408 465172 3420
rect 465224 3408 465230 3460
rect 468478 3408 468484 3460
rect 468536 3448 468542 3460
rect 469858 3448 469864 3460
rect 468536 3420 469864 3448
rect 468536 3408 468542 3420
rect 469858 3408 469864 3420
rect 469916 3408 469922 3460
rect 470566 3448 470594 3488
rect 472618 3476 472624 3528
rect 472676 3516 472682 3528
rect 473446 3516 473452 3528
rect 472676 3488 473452 3516
rect 472676 3476 472682 3488
rect 473446 3476 473452 3488
rect 473504 3476 473510 3528
rect 475378 3476 475384 3528
rect 475436 3516 475442 3528
rect 475436 3488 480254 3516
rect 475436 3476 475442 3488
rect 475746 3448 475752 3460
rect 470566 3420 475752 3448
rect 475746 3408 475752 3420
rect 475804 3408 475810 3460
rect 480226 3448 480254 3488
rect 486510 3476 486516 3528
rect 486568 3516 486574 3528
rect 487614 3516 487620 3528
rect 486568 3488 487620 3516
rect 486568 3476 486574 3488
rect 487614 3476 487620 3488
rect 487672 3476 487678 3528
rect 493318 3476 493324 3528
rect 493376 3516 493382 3528
rect 493376 3488 509234 3516
rect 493376 3476 493382 3488
rect 507670 3448 507676 3460
rect 480226 3420 507676 3448
rect 507670 3408 507676 3420
rect 507728 3408 507734 3460
rect 207658 3340 207664 3392
rect 207716 3380 207722 3392
rect 223942 3380 223948 3392
rect 207716 3352 223948 3380
rect 207716 3340 207722 3352
rect 223942 3340 223948 3352
rect 224000 3340 224006 3392
rect 225598 3340 225604 3392
rect 225656 3380 225662 3392
rect 226334 3380 226340 3392
rect 225656 3352 226340 3380
rect 225656 3340 225662 3352
rect 226334 3340 226340 3352
rect 226392 3340 226398 3392
rect 239398 3340 239404 3392
rect 239456 3380 239462 3392
rect 240502 3380 240508 3392
rect 239456 3352 240508 3380
rect 239456 3340 239462 3352
rect 240502 3340 240508 3352
rect 240560 3340 240566 3392
rect 275278 3340 275284 3392
rect 275336 3380 275342 3392
rect 276014 3380 276020 3392
rect 275336 3352 276020 3380
rect 275336 3340 275342 3352
rect 276014 3340 276020 3352
rect 276072 3340 276078 3392
rect 307018 3340 307024 3392
rect 307076 3380 307082 3392
rect 309042 3380 309048 3392
rect 307076 3352 309048 3380
rect 307076 3340 307082 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 329098 3340 329104 3392
rect 329156 3380 329162 3392
rect 330386 3380 330392 3392
rect 329156 3352 330392 3380
rect 329156 3340 329162 3352
rect 330386 3340 330392 3352
rect 330444 3340 330450 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 340966 3340 340972 3392
rect 341024 3380 341030 3392
rect 342162 3380 342168 3392
rect 341024 3352 342168 3380
rect 341024 3340 341030 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 357526 3340 357532 3392
rect 357584 3380 357590 3392
rect 358722 3380 358728 3392
rect 357584 3352 358728 3380
rect 357584 3340 357590 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 364978 3340 364984 3392
rect 365036 3380 365042 3392
rect 367002 3380 367008 3392
rect 365036 3352 367008 3380
rect 365036 3340 365042 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 390554 3340 390560 3392
rect 390612 3380 390618 3392
rect 391842 3380 391848 3392
rect 390612 3352 391848 3380
rect 390612 3340 390618 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 400858 3340 400864 3392
rect 400916 3380 400922 3392
rect 402514 3380 402520 3392
rect 400916 3352 402520 3380
rect 400916 3340 400922 3352
rect 402514 3340 402520 3352
rect 402572 3340 402578 3392
rect 414658 3340 414664 3392
rect 414716 3380 414722 3392
rect 416682 3380 416688 3392
rect 414716 3352 416688 3380
rect 414716 3340 414722 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 418798 3340 418804 3392
rect 418856 3380 418862 3392
rect 420178 3380 420184 3392
rect 418856 3352 420184 3380
rect 418856 3340 418862 3352
rect 420178 3340 420184 3352
rect 420236 3340 420242 3392
rect 422938 3340 422944 3392
rect 422996 3380 423002 3392
rect 424962 3380 424968 3392
rect 422996 3352 424968 3380
rect 422996 3340 423002 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 432598 3340 432604 3392
rect 432656 3380 432662 3392
rect 434438 3380 434444 3392
rect 432656 3352 434444 3380
rect 432656 3340 432662 3352
rect 434438 3340 434444 3352
rect 434496 3340 434502 3392
rect 440234 3340 440240 3392
rect 440292 3380 440298 3392
rect 441522 3380 441528 3392
rect 440292 3352 441528 3380
rect 440292 3340 440298 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 446398 3340 446404 3392
rect 446456 3380 446462 3392
rect 447410 3380 447416 3392
rect 446456 3352 447416 3380
rect 446456 3340 446462 3352
rect 447410 3340 447416 3352
rect 447468 3340 447474 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 456886 3340 456892 3392
rect 456944 3380 456950 3392
rect 458082 3380 458088 3392
rect 456944 3352 458088 3380
rect 456944 3340 456950 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 509206 3380 509234 3488
rect 514018 3476 514024 3528
rect 514076 3516 514082 3528
rect 515950 3516 515956 3528
rect 514076 3488 515956 3516
rect 514076 3476 514082 3488
rect 515950 3476 515956 3488
rect 516008 3476 516014 3528
rect 545758 3476 545764 3528
rect 545816 3516 545822 3528
rect 551462 3516 551468 3528
rect 545816 3488 551468 3516
rect 545816 3476 545822 3488
rect 551462 3476 551468 3488
rect 551520 3476 551526 3528
rect 554038 3476 554044 3528
rect 554096 3516 554102 3528
rect 554958 3516 554964 3528
rect 554096 3488 554964 3516
rect 554096 3476 554102 3488
rect 554958 3476 554964 3488
rect 555016 3476 555022 3528
rect 560938 3476 560944 3528
rect 560996 3516 561002 3528
rect 564434 3516 564440 3528
rect 560996 3488 564440 3516
rect 560996 3476 561002 3488
rect 564434 3476 564440 3488
rect 564492 3476 564498 3528
rect 571978 3476 571984 3528
rect 572036 3516 572042 3528
rect 573910 3516 573916 3528
rect 572036 3488 573916 3516
rect 572036 3476 572042 3488
rect 573910 3476 573916 3488
rect 573968 3476 573974 3528
rect 511350 3408 511356 3460
rect 511408 3448 511414 3460
rect 514754 3448 514760 3460
rect 511408 3420 514760 3448
rect 511408 3408 511414 3420
rect 514754 3408 514760 3420
rect 514812 3408 514818 3460
rect 527910 3408 527916 3460
rect 527968 3448 527974 3460
rect 533706 3448 533712 3460
rect 527968 3420 533712 3448
rect 527968 3408 527974 3420
rect 533706 3408 533712 3420
rect 533764 3408 533770 3460
rect 538950 3408 538956 3460
rect 539008 3448 539014 3460
rect 539594 3448 539600 3460
rect 539008 3420 539600 3448
rect 539008 3408 539014 3420
rect 539594 3408 539600 3420
rect 539652 3408 539658 3460
rect 570598 3408 570604 3460
rect 570656 3448 570662 3460
rect 572714 3448 572720 3460
rect 570656 3420 572720 3448
rect 570656 3408 570662 3420
rect 572714 3408 572720 3420
rect 572772 3408 572778 3460
rect 518342 3380 518348 3392
rect 509206 3352 518348 3380
rect 518342 3340 518348 3352
rect 518400 3340 518406 3392
rect 198148 3284 205634 3312
rect 198148 3272 198154 3284
rect 520918 3272 520924 3324
rect 520976 3312 520982 3324
rect 524230 3312 524236 3324
rect 520976 3284 524236 3312
rect 520976 3272 520982 3284
rect 524230 3272 524236 3284
rect 524288 3272 524294 3324
rect 125870 3204 125876 3256
rect 125928 3244 125934 3256
rect 131482 3244 131488 3256
rect 125928 3216 131488 3244
rect 125928 3204 125934 3216
rect 131482 3204 131488 3216
rect 131540 3204 131546 3256
rect 342990 3204 342996 3256
rect 343048 3244 343054 3256
rect 344554 3244 344560 3256
rect 343048 3216 344560 3244
rect 343048 3204 343054 3216
rect 344554 3204 344560 3216
rect 344612 3204 344618 3256
rect 552750 3204 552756 3256
rect 552808 3244 552814 3256
rect 553762 3244 553768 3256
rect 552808 3216 553768 3244
rect 552808 3204 552814 3216
rect 553762 3204 553768 3216
rect 553820 3204 553826 3256
rect 131114 3176 131120 3188
rect 122806 3148 131120 3176
rect 131114 3136 131120 3148
rect 131172 3136 131178 3188
rect 136450 3136 136456 3188
rect 136508 3176 136514 3188
rect 139946 3176 139952 3188
rect 136508 3148 139952 3176
rect 136508 3136 136514 3148
rect 139946 3136 139952 3148
rect 140004 3136 140010 3188
rect 148502 3136 148508 3188
rect 148560 3176 148566 3188
rect 154206 3176 154212 3188
rect 148560 3148 154212 3176
rect 148560 3136 148566 3148
rect 154206 3136 154212 3148
rect 154264 3136 154270 3188
rect 220078 3136 220084 3188
rect 220136 3176 220142 3188
rect 222746 3176 222752 3188
rect 220136 3148 222752 3176
rect 220136 3136 220142 3148
rect 222746 3136 222752 3148
rect 222804 3136 222810 3188
rect 315298 3136 315304 3188
rect 315356 3176 315362 3188
rect 317322 3176 317328 3188
rect 315356 3148 317328 3176
rect 315356 3136 315362 3148
rect 317322 3136 317328 3148
rect 317380 3136 317386 3188
rect 538858 3136 538864 3188
rect 538916 3176 538922 3188
rect 546678 3176 546684 3188
rect 538916 3148 546684 3176
rect 538916 3136 538922 3148
rect 546678 3136 546684 3148
rect 546736 3136 546742 3188
rect 217318 3068 217324 3120
rect 217376 3108 217382 3120
rect 218054 3108 218060 3120
rect 217376 3080 218060 3108
rect 217376 3068 217382 3080
rect 218054 3068 218060 3080
rect 218112 3068 218118 3120
rect 1670 3000 1676 3052
rect 1728 3040 1734 3052
rect 9030 3040 9036 3052
rect 1728 3012 9036 3040
rect 1728 3000 1734 3012
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 19426 3000 19432 3052
rect 19484 3040 19490 3052
rect 21358 3040 21364 3052
rect 19484 3012 21364 3040
rect 19484 3000 19490 3012
rect 21358 3000 21364 3012
rect 21416 3000 21422 3052
rect 23014 3000 23020 3052
rect 23072 3040 23078 3052
rect 25498 3040 25504 3052
rect 23072 3012 25504 3040
rect 23072 3000 23078 3012
rect 25498 3000 25504 3012
rect 25556 3000 25562 3052
rect 118786 3000 118792 3052
rect 118844 3040 118850 3052
rect 120718 3040 120724 3052
rect 118844 3012 120724 3040
rect 118844 3000 118850 3012
rect 120718 3000 120724 3012
rect 120776 3000 120782 3052
rect 123478 3000 123484 3052
rect 123536 3040 123542 3052
rect 125594 3040 125600 3052
rect 123536 3012 125600 3040
rect 123536 3000 123542 3012
rect 125594 3000 125600 3012
rect 125652 3000 125658 3052
rect 141234 3000 141240 3052
rect 141292 3040 141298 3052
rect 142706 3040 142712 3052
rect 141292 3012 142712 3040
rect 141292 3000 141298 3012
rect 142706 3000 142712 3012
rect 142764 3000 142770 3052
rect 182910 3000 182916 3052
rect 182968 3040 182974 3052
rect 186130 3040 186136 3052
rect 182968 3012 186136 3040
rect 182968 3000 182974 3012
rect 186130 3000 186136 3012
rect 186188 3000 186194 3052
rect 324958 3000 324964 3052
rect 325016 3040 325022 3052
rect 326798 3040 326804 3052
rect 325016 3012 326804 3040
rect 325016 3000 325022 3012
rect 326798 3000 326804 3012
rect 326856 3000 326862 3052
rect 382918 3000 382924 3052
rect 382976 3040 382982 3052
rect 384758 3040 384764 3052
rect 382976 3012 384764 3040
rect 382976 3000 382982 3012
rect 384758 3000 384764 3012
rect 384816 3000 384822 3052
rect 464338 3000 464344 3052
rect 464396 3040 464402 3052
rect 466270 3040 466276 3052
rect 464396 3012 466276 3040
rect 464396 3000 464402 3012
rect 466270 3000 466276 3012
rect 466328 3000 466334 3052
rect 503070 3000 503076 3052
rect 503128 3040 503134 3052
rect 505370 3040 505376 3052
rect 503128 3012 505376 3040
rect 503128 3000 503134 3012
rect 505370 3000 505376 3012
rect 505428 3000 505434 3052
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 14458 2972 14464 2984
rect 12400 2944 14464 2972
rect 12400 2932 12406 2944
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 132954 2932 132960 2984
rect 133012 2972 133018 2984
rect 141418 2972 141424 2984
rect 133012 2944 141424 2972
rect 133012 2932 133018 2944
rect 141418 2932 141424 2944
rect 141476 2932 141482 2984
rect 171870 2932 171876 2984
rect 171928 2972 171934 2984
rect 174262 2972 174268 2984
rect 171928 2944 174268 2972
rect 171928 2932 171934 2944
rect 174262 2932 174268 2944
rect 174320 2932 174326 2984
rect 70302 2864 70308 2916
rect 70360 2904 70366 2916
rect 72418 2904 72424 2916
rect 70360 2876 72424 2904
rect 70360 2864 70366 2876
rect 72418 2864 72424 2876
rect 72476 2864 72482 2916
rect 203518 2864 203524 2916
rect 203576 2904 203582 2916
rect 207382 2904 207388 2916
rect 203576 2876 207388 2904
rect 203576 2864 203582 2876
rect 207382 2864 207388 2876
rect 207440 2864 207446 2916
rect 480898 2864 480904 2916
rect 480956 2904 480962 2916
rect 484026 2904 484032 2916
rect 480956 2876 484032 2904
rect 480956 2864 480962 2876
rect 484026 2864 484032 2876
rect 484084 2864 484090 2916
rect 382274 960 382280 1012
rect 382332 1000 382338 1012
rect 383562 1000 383568 1012
rect 382332 972 383568 1000
rect 382332 960 382338 972
rect 383562 960 383568 972
rect 383620 960 383626 1012
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 137836 700680 137888 700732
rect 157340 700680 157392 700732
rect 155960 700612 156012 700664
rect 202788 700612 202840 700664
rect 157248 700544 157300 700596
rect 218980 700544 219032 700596
rect 89168 700476 89220 700528
rect 160744 700476 160796 700528
rect 24308 700408 24360 700460
rect 162216 700408 162268 700460
rect 8116 700340 8168 700392
rect 162124 700340 162176 700392
rect 148324 700272 148376 700324
rect 543464 700272 543516 700324
rect 543004 700204 543056 700256
rect 559656 700272 559708 700324
rect 105452 699660 105504 699712
rect 106924 699660 106976 699712
rect 265624 699660 265676 699712
rect 267648 699660 267700 699712
rect 347044 699660 347096 699712
rect 348792 699660 348844 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 428464 699660 428516 699712
rect 429844 699660 429896 699712
rect 146300 696940 146352 696992
rect 580172 696940 580224 696992
rect 3424 683204 3476 683256
rect 161480 683204 161532 683256
rect 146944 683136 146996 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 163504 670692 163556 670744
rect 185584 670692 185636 670744
rect 580172 670692 580224 670744
rect 149704 660288 149756 660340
rect 462320 660288 462372 660340
rect 3424 656888 3476 656940
rect 163596 656888 163648 656940
rect 182824 643084 182876 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 164240 632068 164292 632120
rect 198004 630640 198056 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 164884 618264 164936 618316
rect 143540 616836 143592 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 164976 605820 165028 605872
rect 142160 590656 142212 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 165620 579640 165672 579692
rect 144184 576852 144236 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 167644 565836 167696 565888
rect 142436 563048 142488 563100
rect 579804 563048 579856 563100
rect 3424 553392 3476 553444
rect 165712 553392 165764 553444
rect 188344 536800 188396 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 167000 527144 167052 527196
rect 142804 524424 142856 524476
rect 580172 524424 580224 524476
rect 2780 514768 2832 514820
rect 4804 514768 4856 514820
rect 181444 510620 181496 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 167276 500964 167328 501016
rect 139400 484372 139452 484424
rect 580172 484372 580224 484424
rect 140044 470568 140096 470620
rect 579988 470568 580040 470620
rect 3516 462340 3568 462392
rect 170404 462340 170456 462392
rect 180064 456764 180116 456816
rect 580172 456764 580224 456816
rect 3148 448536 3200 448588
rect 170496 448536 170548 448588
rect 157432 447788 157484 447840
rect 169760 447788 169812 447840
rect 138664 430584 138716 430636
rect 580172 430584 580224 430636
rect 3516 422288 3568 422340
rect 169760 422288 169812 422340
rect 138756 418140 138808 418192
rect 580172 418140 580224 418192
rect 2872 409844 2924 409896
rect 171784 409844 171836 409896
rect 184204 404336 184256 404388
rect 580172 404336 580224 404388
rect 3516 397468 3568 397520
rect 171876 397468 171928 397520
rect 178684 378156 178736 378208
rect 580172 378156 580224 378208
rect 3516 371220 3568 371272
rect 152464 371220 152516 371272
rect 3148 357416 3200 357468
rect 113824 357416 113876 357468
rect 135260 351908 135312 351960
rect 580172 351908 580224 351960
rect 3516 345176 3568 345228
rect 7564 345176 7616 345228
rect 134524 324300 134576 324352
rect 580172 324300 580224 324352
rect 3332 318792 3384 318844
rect 173900 318792 173952 318844
rect 135904 311856 135956 311908
rect 579988 311856 580040 311908
rect 3516 304988 3568 305040
rect 175924 304988 175976 305040
rect 134616 298120 134668 298172
rect 580172 298120 580224 298172
rect 3516 292544 3568 292596
rect 174544 292544 174596 292596
rect 113824 291796 113876 291848
rect 173164 291796 173216 291848
rect 4804 289076 4856 289128
rect 169024 289076 169076 289128
rect 151084 287648 151136 287700
rect 477500 287648 477552 287700
rect 145564 286288 145616 286340
rect 198004 286288 198056 286340
rect 189080 284928 189132 284980
rect 265624 284928 265676 284980
rect 154580 284316 154632 284368
rect 189080 284316 189132 284368
rect 207020 283568 207072 283620
rect 364340 283568 364392 283620
rect 151820 282888 151872 282940
rect 207020 282888 207072 282940
rect 147956 280780 148008 280832
rect 527180 280780 527232 280832
rect 144920 279420 144972 279472
rect 182824 279420 182876 279472
rect 141424 277992 141476 278044
rect 188344 277992 188396 278044
rect 137284 276632 137336 276684
rect 184204 276632 184256 276684
rect 40040 275272 40092 275324
rect 160100 275272 160152 275324
rect 187700 275272 187752 275324
rect 331220 275272 331272 275324
rect 153384 274660 153436 274712
rect 187700 274660 187752 274712
rect 71780 273912 71832 273964
rect 159364 273912 159416 273964
rect 189172 273912 189224 273964
rect 234620 273912 234672 273964
rect 156052 273232 156104 273284
rect 189172 273232 189224 273284
rect 132500 271872 132552 271924
rect 580172 271872 580224 271924
rect 137376 271192 137428 271244
rect 178684 271192 178736 271244
rect 149060 271124 149112 271176
rect 494060 271124 494112 271176
rect 7564 269832 7616 269884
rect 172704 269832 172756 269884
rect 147772 269764 147824 269816
rect 543004 269764 543056 269816
rect 3424 268336 3476 268388
rect 120816 268336 120868 268388
rect 146208 268336 146260 268388
rect 185584 268336 185636 268388
rect 120816 267724 120868 267776
rect 168380 267724 168432 267776
rect 207572 266976 207624 267028
rect 299480 266976 299532 267028
rect 154396 266432 154448 266484
rect 207572 266432 207624 266484
rect 3056 266364 3108 266416
rect 175924 266364 175976 266416
rect 152464 265752 152516 265804
rect 173348 265752 173400 265804
rect 141332 265684 141384 265736
rect 181444 265684 181496 265736
rect 106924 265616 106976 265668
rect 158720 265616 158772 265668
rect 174544 265616 174596 265668
rect 194876 265616 194928 265668
rect 172796 265548 172848 265600
rect 196256 265548 196308 265600
rect 173440 265480 173492 265532
rect 197360 265480 197412 265532
rect 164884 265412 164936 265464
rect 165436 265412 165488 265464
rect 170220 265412 170272 265464
rect 170496 265412 170548 265464
rect 196164 265412 196216 265464
rect 171784 265344 171836 265396
rect 199016 265344 199068 265396
rect 170404 265276 170456 265328
rect 170680 265276 170732 265328
rect 199200 265276 199252 265328
rect 118332 265208 118384 265260
rect 138756 265208 138808 265260
rect 168748 265208 168800 265260
rect 169024 265208 169076 265260
rect 198004 265208 198056 265260
rect 114192 265140 114244 265192
rect 135904 265140 135956 265192
rect 160836 265140 160888 265192
rect 194784 265140 194836 265192
rect 119988 265072 120040 265124
rect 146944 265072 146996 265124
rect 163504 265072 163556 265124
rect 197912 265072 197964 265124
rect 119896 265004 119948 265056
rect 148508 265004 148560 265056
rect 157248 265004 157300 265056
rect 192208 265004 192260 265056
rect 120724 264936 120776 264988
rect 150716 264936 150768 264988
rect 151084 264936 151136 264988
rect 165436 264936 165488 264988
rect 203248 264936 203300 264988
rect 139492 264188 139544 264240
rect 180064 264188 180116 264240
rect 204812 264188 204864 264240
rect 428464 264188 428516 264240
rect 172612 263848 172664 263900
rect 173348 263848 173400 263900
rect 190644 263848 190696 263900
rect 175740 263780 175792 263832
rect 199292 263780 199344 263832
rect 115480 263712 115532 263764
rect 134432 263712 134484 263764
rect 134616 263712 134668 263764
rect 158720 263712 158772 263764
rect 159272 263712 159324 263764
rect 190736 263712 190788 263764
rect 115572 263644 115624 263696
rect 137284 263644 137336 263696
rect 137560 263644 137612 263696
rect 153200 263644 153252 263696
rect 158812 263644 158864 263696
rect 193772 263644 193824 263696
rect 111524 263576 111576 263628
rect 137376 263576 137428 263628
rect 150900 263576 150952 263628
rect 204812 263576 204864 263628
rect 137468 263440 137520 263492
rect 580264 263508 580316 263560
rect 153200 263440 153252 263492
rect 153384 263440 153436 263492
rect 171692 263236 171744 263288
rect 171876 263236 171928 263288
rect 177764 263168 177816 263220
rect 193956 263168 194008 263220
rect 3424 263100 3476 263152
rect 178040 263100 178092 263152
rect 118148 263032 118200 263084
rect 125968 263032 126020 263084
rect 131120 263032 131172 263084
rect 131764 263032 131816 263084
rect 580540 263032 580592 263084
rect 113824 262964 113876 263016
rect 130108 262964 130160 263016
rect 580356 262964 580408 263016
rect 112352 262896 112404 262948
rect 128360 262896 128412 262948
rect 164976 262896 165028 262948
rect 192392 262896 192444 262948
rect 114100 262828 114152 262880
rect 134524 262828 134576 262880
rect 134800 262828 134852 262880
rect 155868 262828 155920 262880
rect 189356 262828 189408 262880
rect 282920 262828 282972 262880
rect 112628 262760 112680 262812
rect 131120 262760 131172 262812
rect 159364 262760 159416 262812
rect 159916 262760 159968 262812
rect 194048 262760 194100 262812
rect 113916 262692 113968 262744
rect 133052 262692 133104 262744
rect 171692 262692 171744 262744
rect 206008 262692 206060 262744
rect 109776 262624 109828 262676
rect 138664 262624 138716 262676
rect 162216 262624 162268 262676
rect 204628 262624 204680 262676
rect 3608 262556 3660 262608
rect 176752 262556 176804 262608
rect 182916 262556 182968 262608
rect 190460 262556 190512 262608
rect 3516 262488 3568 262540
rect 178408 262488 178460 262540
rect 115388 262420 115440 262472
rect 123208 262420 123260 262472
rect 178040 262420 178092 262472
rect 194968 262420 195020 262472
rect 116860 262352 116912 262404
rect 127624 262352 127676 262404
rect 132040 262352 132092 262404
rect 580448 262352 580500 262404
rect 121368 262284 121420 262336
rect 128728 262284 128780 262336
rect 183468 262284 183520 262336
rect 190828 262284 190880 262336
rect 181260 262216 181312 262268
rect 190552 262216 190604 262268
rect 4804 261400 4856 261452
rect 177764 261400 177816 261452
rect 115296 261332 115348 261384
rect 137468 261332 137520 261384
rect 176752 261332 176804 261384
rect 197820 261332 197872 261384
rect 133052 261264 133104 261316
rect 472624 261264 472676 261316
rect 116492 261196 116544 261248
rect 134340 261196 134392 261248
rect 180156 261196 180208 261248
rect 193680 261196 193732 261248
rect 121276 261128 121328 261180
rect 132040 261128 132092 261180
rect 180524 261128 180576 261180
rect 195060 261128 195112 261180
rect 118056 261060 118108 261112
rect 131120 261060 131172 261112
rect 181996 261060 182048 261112
rect 199108 261060 199160 261112
rect 119528 260992 119580 261044
rect 125600 260992 125652 261044
rect 178408 260992 178460 261044
rect 196440 260992 196492 261044
rect 119620 260924 119672 260976
rect 127072 260924 127124 260976
rect 181812 260924 181864 260976
rect 192116 260924 192168 260976
rect 119252 260856 119304 260908
rect 130384 260856 130436 260908
rect 184756 260856 184808 260908
rect 196348 260856 196400 260908
rect 119436 260788 119488 260840
rect 124312 260788 124364 260840
rect 167276 260788 167328 260840
rect 168196 260788 168248 260840
rect 117872 260720 117924 260772
rect 122840 260720 122892 260772
rect 173900 260380 173952 260432
rect 181904 260380 181956 260432
rect 134340 260312 134392 260364
rect 187792 260312 187844 260364
rect 166632 260244 166684 260296
rect 206100 260244 206152 260296
rect 7564 260176 7616 260228
rect 176200 260176 176252 260228
rect 184112 260176 184164 260228
rect 192484 260176 192536 260228
rect 157340 260108 157392 260160
rect 158306 260108 158358 260160
rect 165712 260108 165764 260160
rect 166586 260108 166638 260160
rect 169760 260108 169812 260160
rect 171002 260108 171054 260160
rect 200580 260108 200632 260160
rect 116400 260040 116452 260092
rect 147956 260040 148008 260092
rect 167000 260040 167052 260092
rect 167690 260040 167742 260092
rect 116676 259972 116728 260024
rect 139400 259972 139452 260024
rect 181904 260040 181956 260092
rect 193864 260040 193916 260092
rect 189264 259972 189316 260024
rect 119344 259904 119396 259956
rect 132500 259904 132552 259956
rect 133144 259904 133196 259956
rect 166356 259904 166408 259956
rect 190920 259904 190972 259956
rect 117964 259836 118016 259888
rect 140872 259836 140924 259888
rect 176108 259836 176160 259888
rect 203340 259836 203392 259888
rect 115204 259768 115256 259820
rect 139676 259768 139728 259820
rect 168104 259768 168156 259820
rect 196624 259768 196676 259820
rect 116584 259700 116636 259752
rect 142436 259700 142488 259752
rect 158076 259700 158128 259752
rect 189724 259700 189776 259752
rect 112536 259632 112588 259684
rect 142160 259632 142212 259684
rect 143080 259632 143132 259684
rect 158628 259632 158680 259684
rect 184112 259632 184164 259684
rect 184572 259632 184624 259684
rect 192576 259632 192628 259684
rect 112812 259564 112864 259616
rect 124864 259564 124916 259616
rect 179420 259564 179472 259616
rect 189632 259564 189684 259616
rect 113732 259496 113784 259548
rect 129280 259496 129332 259548
rect 184020 259496 184072 259548
rect 207664 259496 207716 259548
rect 112904 259428 112956 259480
rect 126520 259428 126572 259480
rect 176384 259428 176436 259480
rect 196532 259428 196584 259480
rect 187792 259360 187844 259412
rect 580172 259360 580224 259412
rect 472624 245556 472676 245608
rect 579712 245556 579764 245608
rect 3332 241068 3384 241120
rect 7564 241068 7616 241120
rect 2780 215228 2832 215280
rect 4804 215228 4856 215280
rect 471244 206932 471296 206984
rect 580172 206932 580224 206984
rect 123944 200676 123996 200728
rect 120632 200608 120684 200660
rect 131856 200676 131908 200728
rect 132040 200676 132092 200728
rect 108948 200540 109000 200592
rect 132224 200540 132276 200592
rect 123944 200472 123996 200524
rect 129004 200472 129056 200524
rect 132040 200472 132092 200524
rect 107568 200404 107620 200456
rect 120632 200404 120684 200456
rect 118608 200336 118660 200388
rect 131856 200336 131908 200388
rect 118516 200268 118568 200320
rect 117228 200200 117280 200252
rect 129648 200132 129700 200184
rect 119436 200064 119488 200116
rect 125048 200064 125100 200116
rect 126612 199996 126664 200048
rect 130660 199928 130712 199980
rect 129280 199860 129332 199912
rect 132914 199860 132966 199912
rect 133006 199860 133058 199912
rect 133098 199860 133150 199912
rect 133742 199860 133794 199912
rect 133926 199860 133978 199912
rect 134110 199860 134162 199912
rect 134386 199860 134438 199912
rect 134478 199860 134530 199912
rect 134662 199860 134714 199912
rect 134846 199860 134898 199912
rect 127164 199792 127216 199844
rect 132546 199792 132598 199844
rect 126980 199724 127032 199776
rect 133696 199724 133748 199776
rect 133972 199724 134024 199776
rect 134064 199724 134116 199776
rect 134294 199724 134346 199776
rect 134386 199724 134438 199776
rect 134616 199724 134668 199776
rect 134708 199724 134760 199776
rect 132316 199656 132368 199708
rect 135030 199656 135082 199708
rect 104532 199588 104584 199640
rect 135306 199860 135358 199912
rect 135398 199860 135450 199912
rect 135582 199860 135634 199912
rect 135674 199860 135726 199912
rect 135720 199656 135772 199708
rect 135950 199860 136002 199912
rect 136042 199860 136094 199912
rect 136134 199860 136186 199912
rect 136318 199860 136370 199912
rect 136502 199860 136554 199912
rect 136686 199860 136738 199912
rect 135996 199724 136048 199776
rect 136364 199724 136416 199776
rect 136088 199656 136140 199708
rect 136732 199724 136784 199776
rect 135444 199588 135496 199640
rect 135628 199588 135680 199640
rect 135812 199588 135864 199640
rect 136548 199588 136600 199640
rect 136732 199588 136784 199640
rect 137054 199860 137106 199912
rect 137330 199860 137382 199912
rect 137882 199860 137934 199912
rect 137974 199860 138026 199912
rect 137146 199792 137198 199844
rect 137100 199656 137152 199708
rect 136916 199588 136968 199640
rect 137376 199724 137428 199776
rect 137928 199656 137980 199708
rect 138250 199860 138302 199912
rect 138342 199860 138394 199912
rect 138526 199860 138578 199912
rect 138802 199860 138854 199912
rect 137836 199588 137888 199640
rect 138112 199588 138164 199640
rect 138296 199588 138348 199640
rect 138572 199724 138624 199776
rect 139262 199860 139314 199912
rect 139354 199860 139406 199912
rect 139446 199860 139498 199912
rect 139538 199860 139590 199912
rect 139722 199860 139774 199912
rect 139906 199860 139958 199912
rect 139998 199860 140050 199912
rect 140274 199860 140326 199912
rect 139216 199724 139268 199776
rect 139492 199724 139544 199776
rect 139308 199656 139360 199708
rect 139400 199656 139452 199708
rect 139768 199724 139820 199776
rect 139860 199724 139912 199776
rect 139952 199724 140004 199776
rect 138664 199588 138716 199640
rect 138756 199588 138808 199640
rect 140366 199792 140418 199844
rect 140412 199588 140464 199640
rect 140734 199860 140786 199912
rect 140826 199860 140878 199912
rect 141010 199860 141062 199912
rect 140688 199724 140740 199776
rect 140964 199724 141016 199776
rect 140780 199656 140832 199708
rect 140872 199656 140924 199708
rect 141746 199860 141798 199912
rect 141838 199860 141890 199912
rect 142022 199860 142074 199912
rect 142114 199860 142166 199912
rect 142206 199860 142258 199912
rect 142298 199860 142350 199912
rect 142390 199860 142442 199912
rect 141562 199792 141614 199844
rect 141516 199656 141568 199708
rect 141608 199588 141660 199640
rect 141792 199588 141844 199640
rect 141976 199588 142028 199640
rect 97632 199520 97684 199572
rect 142758 199860 142810 199912
rect 142252 199724 142304 199776
rect 142252 199588 142304 199640
rect 142712 199724 142764 199776
rect 142344 199520 142396 199572
rect 143126 199860 143178 199912
rect 143218 199860 143270 199912
rect 143402 199860 143454 199912
rect 143494 199860 143546 199912
rect 143080 199588 143132 199640
rect 143310 199792 143362 199844
rect 143448 199724 143500 199776
rect 143678 199860 143730 199912
rect 143770 199860 143822 199912
rect 143954 199860 144006 199912
rect 144046 199860 144098 199912
rect 144138 199860 144190 199912
rect 144230 199860 144282 199912
rect 144322 199860 144374 199912
rect 143816 199724 143868 199776
rect 143908 199724 143960 199776
rect 144000 199656 144052 199708
rect 143632 199588 143684 199640
rect 143172 199520 143224 199572
rect 143264 199520 143316 199572
rect 97908 199452 97960 199504
rect 144276 199724 144328 199776
rect 144368 199724 144420 199776
rect 144782 199860 144834 199912
rect 144966 199860 145018 199912
rect 144736 199724 144788 199776
rect 116952 199384 117004 199436
rect 123576 199384 123628 199436
rect 127900 199384 127952 199436
rect 115664 199316 115716 199368
rect 143724 199384 143776 199436
rect 145150 199724 145202 199776
rect 145104 199588 145156 199640
rect 144552 199520 144604 199572
rect 145012 199520 145064 199572
rect 145518 199860 145570 199912
rect 145610 199860 145662 199912
rect 145702 199860 145754 199912
rect 145794 199860 145846 199912
rect 146254 199860 146306 199912
rect 146346 199860 146398 199912
rect 146714 199860 146766 199912
rect 146990 199860 147042 199912
rect 145472 199724 145524 199776
rect 145564 199656 145616 199708
rect 145656 199656 145708 199708
rect 145978 199724 146030 199776
rect 146162 199724 146214 199776
rect 145840 199656 145892 199708
rect 145748 199588 145800 199640
rect 145932 199588 145984 199640
rect 146024 199588 146076 199640
rect 146208 199588 146260 199640
rect 144920 199452 144972 199504
rect 145748 199452 145800 199504
rect 146484 199656 146536 199708
rect 146392 199588 146444 199640
rect 146668 199588 146720 199640
rect 147358 199724 147410 199776
rect 146576 199520 146628 199572
rect 147128 199520 147180 199572
rect 146392 199452 146444 199504
rect 146944 199384 146996 199436
rect 147312 199588 147364 199640
rect 147634 199860 147686 199912
rect 147726 199860 147778 199912
rect 147818 199860 147870 199912
rect 147910 199860 147962 199912
rect 148094 199860 148146 199912
rect 148186 199860 148238 199912
rect 148278 199860 148330 199912
rect 148370 199792 148422 199844
rect 148140 199724 148192 199776
rect 148232 199724 148284 199776
rect 147772 199656 147824 199708
rect 147864 199656 147916 199708
rect 147680 199588 147732 199640
rect 147956 199588 148008 199640
rect 148554 199860 148606 199912
rect 147588 199520 147640 199572
rect 148324 199520 148376 199572
rect 148830 199860 148882 199912
rect 148600 199588 148652 199640
rect 148692 199588 148744 199640
rect 149198 199860 149250 199912
rect 149382 199860 149434 199912
rect 149474 199860 149526 199912
rect 149566 199860 149618 199912
rect 149658 199860 149710 199912
rect 149842 199860 149894 199912
rect 150026 199860 150078 199912
rect 150118 199860 150170 199912
rect 150394 199860 150446 199912
rect 150486 199860 150538 199912
rect 149290 199724 149342 199776
rect 148876 199452 148928 199504
rect 149750 199792 149802 199844
rect 149934 199792 149986 199844
rect 149612 199656 149664 199708
rect 149704 199656 149756 199708
rect 149796 199656 149848 199708
rect 149888 199656 149940 199708
rect 149336 199520 149388 199572
rect 149520 199520 149572 199572
rect 149980 199452 150032 199504
rect 149428 199384 149480 199436
rect 150578 199724 150630 199776
rect 150440 199588 150492 199640
rect 150532 199588 150584 199640
rect 150854 199860 150906 199912
rect 150946 199860 150998 199912
rect 151038 199860 151090 199912
rect 151130 199860 151182 199912
rect 151314 199860 151366 199912
rect 151406 199860 151458 199912
rect 150992 199724 151044 199776
rect 151360 199724 151412 199776
rect 151084 199656 151136 199708
rect 150900 199520 150952 199572
rect 151590 199860 151642 199912
rect 151682 199860 151734 199912
rect 151866 199860 151918 199912
rect 152050 199860 152102 199912
rect 152142 199860 152194 199912
rect 152234 199860 152286 199912
rect 151544 199724 151596 199776
rect 151636 199656 151688 199708
rect 152096 199656 152148 199708
rect 152188 199656 152240 199708
rect 151912 199520 151964 199572
rect 152418 199860 152470 199912
rect 152510 199860 152562 199912
rect 152694 199860 152746 199912
rect 152786 199860 152838 199912
rect 152878 199860 152930 199912
rect 153154 199860 153206 199912
rect 153246 199860 153298 199912
rect 153522 199860 153574 199912
rect 154074 199860 154126 199912
rect 154166 199860 154218 199912
rect 154258 199860 154310 199912
rect 154442 199860 154494 199912
rect 154534 199860 154586 199912
rect 154718 199860 154770 199912
rect 154902 199860 154954 199912
rect 154994 199860 155046 199912
rect 155178 199860 155230 199912
rect 155362 199860 155414 199912
rect 152464 199724 152516 199776
rect 152556 199724 152608 199776
rect 152648 199724 152700 199776
rect 152740 199724 152792 199776
rect 152832 199656 152884 199708
rect 154212 199724 154264 199776
rect 154396 199724 154448 199776
rect 154488 199724 154540 199776
rect 154856 199724 154908 199776
rect 154948 199724 155000 199776
rect 155132 199724 155184 199776
rect 155040 199656 155092 199708
rect 153108 199588 153160 199640
rect 153292 199588 153344 199640
rect 153476 199588 153528 199640
rect 154028 199588 154080 199640
rect 154580 199588 154632 199640
rect 154672 199588 154724 199640
rect 155316 199588 155368 199640
rect 153200 199520 153252 199572
rect 153936 199520 153988 199572
rect 155914 199860 155966 199912
rect 156006 199860 156058 199912
rect 156190 199860 156242 199912
rect 156466 199860 156518 199912
rect 155960 199724 156012 199776
rect 150624 199384 150676 199436
rect 151084 199384 151136 199436
rect 153660 199452 153712 199504
rect 154212 199452 154264 199504
rect 155592 199452 155644 199504
rect 180064 200676 180116 200728
rect 180524 200676 180576 200728
rect 187148 200812 187200 200864
rect 180156 200608 180208 200660
rect 156742 199860 156794 199912
rect 156834 199860 156886 199912
rect 156926 199860 156978 199912
rect 157018 199860 157070 199912
rect 156788 199724 156840 199776
rect 156880 199724 156932 199776
rect 156604 199588 156656 199640
rect 156880 199588 156932 199640
rect 156972 199588 157024 199640
rect 157202 199860 157254 199912
rect 157294 199860 157346 199912
rect 157248 199588 157300 199640
rect 157478 199860 157530 199912
rect 157570 199860 157622 199912
rect 157662 199860 157714 199912
rect 157846 199860 157898 199912
rect 157938 199860 157990 199912
rect 158214 199860 158266 199912
rect 158490 199860 158542 199912
rect 158582 199860 158634 199912
rect 157892 199724 157944 199776
rect 157524 199656 157576 199708
rect 157616 199656 157668 199708
rect 158260 199724 158312 199776
rect 158628 199724 158680 199776
rect 157708 199588 157760 199640
rect 158444 199588 158496 199640
rect 158950 199860 159002 199912
rect 159042 199860 159094 199912
rect 159134 199860 159186 199912
rect 159226 199860 159278 199912
rect 159502 199860 159554 199912
rect 159594 199860 159646 199912
rect 159778 199860 159830 199912
rect 159870 199860 159922 199912
rect 160146 199860 160198 199912
rect 158996 199724 159048 199776
rect 159272 199724 159324 199776
rect 159548 199724 159600 199776
rect 159180 199656 159232 199708
rect 159364 199588 159416 199640
rect 159962 199792 160014 199844
rect 159824 199656 159876 199708
rect 159916 199588 159968 199640
rect 157156 199520 157208 199572
rect 159732 199520 159784 199572
rect 160008 199520 160060 199572
rect 160284 199588 160336 199640
rect 160606 199860 160658 199912
rect 160698 199860 160750 199912
rect 160790 199860 160842 199912
rect 160744 199724 160796 199776
rect 160974 199860 161026 199912
rect 161158 199860 161210 199912
rect 161434 199860 161486 199912
rect 161020 199724 161072 199776
rect 161112 199724 161164 199776
rect 161204 199588 161256 199640
rect 160468 199520 160520 199572
rect 160928 199520 160980 199572
rect 161618 199860 161670 199912
rect 161710 199860 161762 199912
rect 162078 199860 162130 199912
rect 162262 199860 162314 199912
rect 162538 199860 162590 199912
rect 162630 199860 162682 199912
rect 162814 199860 162866 199912
rect 162998 199860 163050 199912
rect 163090 199860 163142 199912
rect 161664 199724 161716 199776
rect 161480 199588 161532 199640
rect 161388 199520 161440 199572
rect 161572 199520 161624 199572
rect 162676 199656 162728 199708
rect 163044 199656 163096 199708
rect 162860 199588 162912 199640
rect 162952 199588 163004 199640
rect 163366 199860 163418 199912
rect 182824 200540 182876 200592
rect 163642 199860 163694 199912
rect 163826 199860 163878 199912
rect 163918 199860 163970 199912
rect 164102 199860 164154 199912
rect 164194 199860 164246 199912
rect 163872 199724 163924 199776
rect 163964 199724 164016 199776
rect 164056 199656 164108 199708
rect 163688 199588 163740 199640
rect 160100 199452 160152 199504
rect 151268 199384 151320 199436
rect 151452 199384 151504 199436
rect 163320 199452 163372 199504
rect 163504 199520 163556 199572
rect 163780 199452 163832 199504
rect 161020 199384 161072 199436
rect 177856 200336 177908 200388
rect 202880 200336 202932 200388
rect 181444 200268 181496 200320
rect 191564 200268 191616 200320
rect 193404 200200 193456 200252
rect 164378 199860 164430 199912
rect 164470 199860 164522 199912
rect 164654 199860 164706 199912
rect 164930 199860 164982 199912
rect 165114 199860 165166 199912
rect 164424 199724 164476 199776
rect 164700 199588 164752 199640
rect 164976 199588 165028 199640
rect 164792 199520 164844 199572
rect 165574 199860 165626 199912
rect 165666 199860 165718 199912
rect 165758 199860 165810 199912
rect 166034 199860 166086 199912
rect 166126 199860 166178 199912
rect 166218 199860 166270 199912
rect 166402 199860 166454 199912
rect 166494 199860 166546 199912
rect 166678 199860 166730 199912
rect 165804 199724 165856 199776
rect 165712 199656 165764 199708
rect 165344 199588 165396 199640
rect 165620 199520 165672 199572
rect 164424 199384 164476 199436
rect 114468 199248 114520 199300
rect 142160 199248 142212 199300
rect 151728 199316 151780 199368
rect 153200 199316 153252 199368
rect 153936 199316 153988 199368
rect 146852 199248 146904 199300
rect 115848 199180 115900 199232
rect 148232 199180 148284 199232
rect 151820 199180 151872 199232
rect 159364 199248 159416 199300
rect 164608 199248 164660 199300
rect 156604 199180 156656 199232
rect 164424 199180 164476 199232
rect 165528 199384 165580 199436
rect 166218 199724 166270 199776
rect 166448 199520 166500 199572
rect 166080 199452 166132 199504
rect 166356 199452 166408 199504
rect 167046 199860 167098 199912
rect 167138 199860 167190 199912
rect 167322 199860 167374 199912
rect 167782 199860 167834 199912
rect 167874 199860 167926 199912
rect 168058 199860 168110 199912
rect 166632 199588 166684 199640
rect 166816 199588 166868 199640
rect 167000 199588 167052 199640
rect 167092 199520 167144 199572
rect 167828 199656 167880 199708
rect 168012 199656 168064 199708
rect 167552 199520 167604 199572
rect 168518 199860 168570 199912
rect 168702 199860 168754 199912
rect 168978 199860 169030 199912
rect 169254 199860 169306 199912
rect 169346 199860 169398 199912
rect 168564 199724 168616 199776
rect 168656 199724 168708 199776
rect 167276 199452 167328 199504
rect 168012 199452 168064 199504
rect 168564 199452 168616 199504
rect 169714 199860 169766 199912
rect 169116 199588 169168 199640
rect 169576 199588 169628 199640
rect 169300 199520 169352 199572
rect 169392 199520 169444 199572
rect 169990 199860 170042 199912
rect 170450 199860 170502 199912
rect 170634 199860 170686 199912
rect 170818 199860 170870 199912
rect 170496 199724 170548 199776
rect 170588 199724 170640 199776
rect 181444 200064 181496 200116
rect 178500 199996 178552 200048
rect 171278 199860 171330 199912
rect 171370 199860 171422 199912
rect 171462 199860 171514 199912
rect 170036 199588 170088 199640
rect 170772 199588 170824 199640
rect 171416 199588 171468 199640
rect 171048 199520 171100 199572
rect 171324 199520 171376 199572
rect 171922 199860 171974 199912
rect 172014 199860 172066 199912
rect 172290 199860 172342 199912
rect 172474 199860 172526 199912
rect 172750 199860 172802 199912
rect 172842 199860 172894 199912
rect 173026 199860 173078 199912
rect 173118 199860 173170 199912
rect 173670 199860 173722 199912
rect 173854 199860 173906 199912
rect 174038 199860 174090 199912
rect 171876 199588 171928 199640
rect 172244 199588 172296 199640
rect 172336 199588 172388 199640
rect 172060 199520 172112 199572
rect 172980 199724 173032 199776
rect 172796 199656 172848 199708
rect 173210 199792 173262 199844
rect 173486 199792 173538 199844
rect 172888 199588 172940 199640
rect 173164 199588 173216 199640
rect 173394 199724 173446 199776
rect 173348 199588 173400 199640
rect 173624 199656 173676 199708
rect 174084 199724 174136 199776
rect 173532 199588 173584 199640
rect 173900 199588 173952 199640
rect 173072 199520 173124 199572
rect 173992 199520 174044 199572
rect 174498 199860 174550 199912
rect 174774 199860 174826 199912
rect 175050 199860 175102 199912
rect 174728 199656 174780 199708
rect 175418 199860 175470 199912
rect 175510 199860 175562 199912
rect 175694 199860 175746 199912
rect 175786 199860 175838 199912
rect 175878 199860 175930 199912
rect 176062 199860 176114 199912
rect 176154 199860 176206 199912
rect 175832 199724 175884 199776
rect 175924 199724 175976 199776
rect 176016 199724 176068 199776
rect 176338 199792 176390 199844
rect 176430 199792 176482 199844
rect 175740 199656 175792 199708
rect 176108 199656 176160 199708
rect 176292 199656 176344 199708
rect 175464 199588 175516 199640
rect 175556 199588 175608 199640
rect 176384 199588 176436 199640
rect 174268 199520 174320 199572
rect 174452 199520 174504 199572
rect 175096 199520 175148 199572
rect 175372 199520 175424 199572
rect 176200 199520 176252 199572
rect 176614 199860 176666 199912
rect 176798 199860 176850 199912
rect 177166 199860 177218 199912
rect 181352 199860 181404 199912
rect 177672 199792 177724 199844
rect 216956 200132 217008 200184
rect 179604 199724 179656 199776
rect 215392 199724 215444 199776
rect 176844 199656 176896 199708
rect 177948 199656 178000 199708
rect 215852 199656 215904 199708
rect 176752 199588 176804 199640
rect 169024 199452 169076 199504
rect 169116 199452 169168 199504
rect 217600 199588 217652 199640
rect 168380 199384 168432 199436
rect 217048 199520 217100 199572
rect 182916 199452 182968 199504
rect 190460 199452 190512 199504
rect 180800 199384 180852 199436
rect 190552 199384 190604 199436
rect 165160 199316 165212 199368
rect 165436 199316 165488 199368
rect 166816 199316 166868 199368
rect 192760 199316 192812 199368
rect 190460 199248 190512 199300
rect 165160 199180 165212 199232
rect 165436 199180 165488 199232
rect 219532 199180 219584 199232
rect 112996 199112 113048 199164
rect 145380 199112 145432 199164
rect 156328 199112 156380 199164
rect 215484 199112 215536 199164
rect 114284 199044 114336 199096
rect 146116 199044 146168 199096
rect 154764 199044 154816 199096
rect 215944 199044 215996 199096
rect 113088 198976 113140 199028
rect 146760 198976 146812 199028
rect 154488 198976 154540 199028
rect 215300 198976 215352 199028
rect 115756 198908 115808 198960
rect 149612 198908 149664 198960
rect 165620 198908 165672 198960
rect 177396 198908 177448 198960
rect 117136 198840 117188 198892
rect 118424 198772 118476 198824
rect 123576 198840 123628 198892
rect 147312 198840 147364 198892
rect 165804 198840 165856 198892
rect 183008 198840 183060 198892
rect 146024 198772 146076 198824
rect 157156 198772 157208 198824
rect 157340 198772 157392 198824
rect 162308 198772 162360 198824
rect 180340 198772 180392 198824
rect 145748 198704 145800 198756
rect 155040 198704 155092 198756
rect 181536 198704 181588 198756
rect 142160 198636 142212 198688
rect 153844 198636 153896 198688
rect 155684 198636 155736 198688
rect 177028 198636 177080 198688
rect 177120 198636 177172 198688
rect 181628 198636 181680 198688
rect 132132 198568 132184 198620
rect 135996 198568 136048 198620
rect 136824 198568 136876 198620
rect 138664 198568 138716 198620
rect 143632 198568 143684 198620
rect 150808 198568 150860 198620
rect 165160 198568 165212 198620
rect 168380 198568 168432 198620
rect 121184 198500 121236 198552
rect 144644 198500 144696 198552
rect 154856 198500 154908 198552
rect 173992 198568 174044 198620
rect 200120 198568 200172 198620
rect 186964 198500 187016 198552
rect 123576 198432 123628 198484
rect 139400 198432 139452 198484
rect 170036 198432 170088 198484
rect 181444 198432 181496 198484
rect 181628 198432 181680 198484
rect 211436 198432 211488 198484
rect 121092 198364 121144 198416
rect 144368 198364 144420 198416
rect 169392 198364 169444 198416
rect 171048 198364 171100 198416
rect 173256 198364 173308 198416
rect 212816 198364 212868 198416
rect 118700 198296 118752 198348
rect 143356 198296 143408 198348
rect 151084 198296 151136 198348
rect 154948 198296 155000 198348
rect 119804 198228 119856 198280
rect 138572 198228 138624 198280
rect 170220 198228 170272 198280
rect 211252 198296 211304 198348
rect 177028 198228 177080 198280
rect 180248 198228 180300 198280
rect 181444 198228 181496 198280
rect 211528 198228 211580 198280
rect 105728 198160 105780 198212
rect 132132 198160 132184 198212
rect 176200 198160 176252 198212
rect 178408 198160 178460 198212
rect 178500 198160 178552 198212
rect 212908 198160 212960 198212
rect 110328 198092 110380 198144
rect 142344 198092 142396 198144
rect 158720 198092 158772 198144
rect 105636 198024 105688 198076
rect 136916 198024 136968 198076
rect 143356 198024 143408 198076
rect 145012 198024 145064 198076
rect 108396 197956 108448 198008
rect 142252 197956 142304 198008
rect 167828 198092 167880 198144
rect 170496 198092 170548 198144
rect 171876 198092 171928 198144
rect 214288 198092 214340 198144
rect 175004 198024 175056 198076
rect 214472 198024 214524 198076
rect 167736 197956 167788 198008
rect 168840 197956 168892 198008
rect 176200 197956 176252 198008
rect 120540 197888 120592 197940
rect 144000 197820 144052 197872
rect 158812 197820 158864 197872
rect 170772 197820 170824 197872
rect 138572 197752 138624 197804
rect 144184 197752 144236 197804
rect 162584 197752 162636 197804
rect 171048 197752 171100 197804
rect 178684 197820 178736 197872
rect 214656 197956 214708 198008
rect 176752 197684 176804 197736
rect 179420 197684 179472 197736
rect 166448 197616 166500 197668
rect 178776 197616 178828 197668
rect 166080 197548 166132 197600
rect 170036 197548 170088 197600
rect 135996 197480 136048 197532
rect 141884 197480 141936 197532
rect 163872 197480 163924 197532
rect 172060 197480 172112 197532
rect 173808 197480 173860 197532
rect 179880 197480 179932 197532
rect 133052 197412 133104 197464
rect 137928 197412 137980 197464
rect 170496 197412 170548 197464
rect 174636 197412 174688 197464
rect 134892 197344 134944 197396
rect 138204 197344 138256 197396
rect 163596 197344 163648 197396
rect 173808 197344 173860 197396
rect 176660 197344 176712 197396
rect 176936 197344 176988 197396
rect 121276 197276 121328 197328
rect 124864 197276 124916 197328
rect 127716 197276 127768 197328
rect 151176 197276 151228 197328
rect 168288 197276 168340 197328
rect 185492 197276 185544 197328
rect 121368 197208 121420 197260
rect 127992 197208 128044 197260
rect 128084 197208 128136 197260
rect 141884 197208 141936 197260
rect 142068 197208 142120 197260
rect 144920 197208 144972 197260
rect 163044 197208 163096 197260
rect 197728 197208 197780 197260
rect 119252 197140 119304 197192
rect 124956 197140 125008 197192
rect 126336 197140 126388 197192
rect 151268 197140 151320 197192
rect 155316 197140 155368 197192
rect 163872 197140 163924 197192
rect 168748 197140 168800 197192
rect 198832 197140 198884 197192
rect 121000 197072 121052 197124
rect 128084 197072 128136 197124
rect 128176 197072 128228 197124
rect 149152 197072 149204 197124
rect 150440 197072 150492 197124
rect 151176 197072 151228 197124
rect 154856 197072 154908 197124
rect 156420 197072 156472 197124
rect 158076 197072 158128 197124
rect 192024 197072 192076 197124
rect 107384 197004 107436 197056
rect 137652 197004 137704 197056
rect 141884 197004 141936 197056
rect 145748 197004 145800 197056
rect 161480 197004 161532 197056
rect 167828 197004 167880 197056
rect 168656 197004 168708 197056
rect 203156 197004 203208 197056
rect 111708 196936 111760 196988
rect 132960 196936 133012 196988
rect 160284 196936 160336 196988
rect 193312 196936 193364 196988
rect 123484 196868 123536 196920
rect 148416 196868 148468 196920
rect 159272 196868 159324 196920
rect 193496 196868 193548 196920
rect 114008 196800 114060 196852
rect 145656 196800 145708 196852
rect 150532 196800 150584 196852
rect 150808 196800 150860 196852
rect 153200 196800 153252 196852
rect 153660 196800 153712 196852
rect 163504 196800 163556 196852
rect 197636 196800 197688 196852
rect 111616 196732 111668 196784
rect 133144 196732 133196 196784
rect 135444 196732 135496 196784
rect 135812 196732 135864 196784
rect 139400 196732 139452 196784
rect 139768 196732 139820 196784
rect 149336 196732 149388 196784
rect 149888 196732 149940 196784
rect 150348 196732 150400 196784
rect 154028 196732 154080 196784
rect 161112 196732 161164 196784
rect 161664 196732 161716 196784
rect 161848 196732 161900 196784
rect 162400 196732 162452 196784
rect 164056 196732 164108 196784
rect 197544 196732 197596 196784
rect 107292 196664 107344 196716
rect 139860 196664 139912 196716
rect 140872 196664 140924 196716
rect 141792 196664 141844 196716
rect 146300 196664 146352 196716
rect 146852 196664 146904 196716
rect 147036 196664 147088 196716
rect 149704 196664 149756 196716
rect 153384 196664 153436 196716
rect 104716 196596 104768 196648
rect 136824 196596 136876 196648
rect 137376 196596 137428 196648
rect 137836 196596 137888 196648
rect 140964 196596 141016 196648
rect 142160 196596 142212 196648
rect 147496 196596 147548 196648
rect 153660 196596 153712 196648
rect 157708 196664 157760 196716
rect 158536 196664 158588 196716
rect 161480 196664 161532 196716
rect 162952 196664 163004 196716
rect 165712 196664 165764 196716
rect 166356 196664 166408 196716
rect 167184 196664 167236 196716
rect 201776 196664 201828 196716
rect 220820 196596 220872 196648
rect 119528 196528 119580 196580
rect 126520 196528 126572 196580
rect 129096 196528 129148 196580
rect 150716 196528 150768 196580
rect 165620 196528 165672 196580
rect 166448 196528 166500 196580
rect 117044 196460 117096 196512
rect 123484 196460 123536 196512
rect 129740 196460 129792 196512
rect 132592 196460 132644 196512
rect 157892 196460 157944 196512
rect 163688 196460 163740 196512
rect 165344 196460 165396 196512
rect 165896 196460 165948 196512
rect 127808 196392 127860 196444
rect 140044 196392 140096 196444
rect 120356 196324 120408 196376
rect 128176 196324 128228 196376
rect 150716 196324 150768 196376
rect 151544 196324 151596 196376
rect 119620 196256 119672 196308
rect 128084 196256 128136 196308
rect 133144 196256 133196 196308
rect 138848 196256 138900 196308
rect 141240 196256 141292 196308
rect 142068 196256 142120 196308
rect 144000 196256 144052 196308
rect 144736 196256 144788 196308
rect 132960 196188 133012 196240
rect 143080 196188 143132 196240
rect 157800 196188 157852 196240
rect 157984 196188 158036 196240
rect 174452 196188 174504 196240
rect 180616 196188 180668 196240
rect 177120 196120 177172 196172
rect 177764 196120 177816 196172
rect 131764 196052 131816 196104
rect 138940 196052 138992 196104
rect 157340 196052 157392 196104
rect 126244 195916 126296 195968
rect 145840 195916 145892 195968
rect 154028 195916 154080 195968
rect 154672 195916 154724 195968
rect 154764 195916 154816 195968
rect 155868 195916 155920 195968
rect 157340 195916 157392 195968
rect 157524 195916 157576 195968
rect 122288 195848 122340 195900
rect 140228 195848 140280 195900
rect 108488 195780 108540 195832
rect 133052 195780 133104 195832
rect 135904 195780 135956 195832
rect 136732 195780 136784 195832
rect 143448 195848 143500 195900
rect 152096 195848 152148 195900
rect 152372 195848 152424 195900
rect 162952 196052 163004 196104
rect 163412 196052 163464 196104
rect 165712 195984 165764 196036
rect 166724 195984 166776 196036
rect 171232 195984 171284 196036
rect 171416 195984 171468 196036
rect 176936 195984 176988 196036
rect 177488 195984 177540 196036
rect 164516 195916 164568 195968
rect 164792 195916 164844 195968
rect 165528 195916 165580 195968
rect 166172 195916 166224 195968
rect 168564 195916 168616 195968
rect 185768 195916 185820 195968
rect 180432 195848 180484 195900
rect 118240 195712 118292 195764
rect 135812 195712 135864 195764
rect 110236 195644 110288 195696
rect 140872 195780 140924 195832
rect 147956 195780 148008 195832
rect 157524 195780 157576 195832
rect 158444 195780 158496 195832
rect 161388 195780 161440 195832
rect 138020 195712 138072 195764
rect 149060 195712 149112 195764
rect 154672 195712 154724 195764
rect 155960 195712 156012 195764
rect 156236 195712 156288 195764
rect 157064 195712 157116 195764
rect 140228 195644 140280 195696
rect 146484 195644 146536 195696
rect 170036 195780 170088 195832
rect 200304 195780 200356 195832
rect 171600 195712 171652 195764
rect 192668 195712 192720 195764
rect 196072 195644 196124 195696
rect 109868 195576 109920 195628
rect 142896 195576 142948 195628
rect 162308 195576 162360 195628
rect 171600 195576 171652 195628
rect 105820 195508 105872 195560
rect 133144 195508 133196 195560
rect 135812 195508 135864 195560
rect 138020 195508 138072 195560
rect 159732 195508 159784 195560
rect 174452 195576 174504 195628
rect 174820 195576 174872 195628
rect 179512 195576 179564 195628
rect 211344 195576 211396 195628
rect 193220 195508 193272 195560
rect 112444 195440 112496 195492
rect 145564 195440 145616 195492
rect 151912 195440 151964 195492
rect 152096 195440 152148 195492
rect 158720 195440 158772 195492
rect 159824 195440 159876 195492
rect 165068 195440 165120 195492
rect 198924 195440 198976 195492
rect 114376 195372 114428 195424
rect 148784 195372 148836 195424
rect 149520 195372 149572 195424
rect 149980 195372 150032 195424
rect 161204 195372 161256 195424
rect 194692 195372 194744 195424
rect 111248 195304 111300 195356
rect 145932 195304 145984 195356
rect 149612 195304 149664 195356
rect 150164 195304 150216 195356
rect 156052 195304 156104 195356
rect 156512 195304 156564 195356
rect 160376 195304 160428 195356
rect 111340 195236 111392 195288
rect 144276 195236 144328 195288
rect 146944 195236 146996 195288
rect 152740 195236 152792 195288
rect 158904 195236 158956 195288
rect 159916 195236 159968 195288
rect 175188 195304 175240 195356
rect 175372 195304 175424 195356
rect 180524 195304 180576 195356
rect 210332 195304 210384 195356
rect 214564 195236 214616 195288
rect 129280 195168 129332 195220
rect 140872 195168 140924 195220
rect 166540 195168 166592 195220
rect 181444 195168 181496 195220
rect 140504 195100 140556 195152
rect 143632 195100 143684 195152
rect 160468 195100 160520 195152
rect 161296 195100 161348 195152
rect 168380 195100 168432 195152
rect 169392 195100 169444 195152
rect 171324 195100 171376 195152
rect 172244 195100 172296 195152
rect 132408 195032 132460 195084
rect 144184 195032 144236 195084
rect 152188 195032 152240 195084
rect 152924 195032 152976 195084
rect 160192 194896 160244 194948
rect 160744 194896 160796 194948
rect 166632 194896 166684 194948
rect 183100 194896 183152 194948
rect 156328 194828 156380 194880
rect 156972 194828 157024 194880
rect 133144 194760 133196 194812
rect 139124 194760 139176 194812
rect 164332 194760 164384 194812
rect 164884 194760 164936 194812
rect 132224 194692 132276 194744
rect 138480 194692 138532 194744
rect 151912 194692 151964 194744
rect 152648 194692 152700 194744
rect 117780 194488 117832 194540
rect 120816 194488 120868 194540
rect 141056 194488 141108 194540
rect 143540 194488 143592 194540
rect 165528 194488 165580 194540
rect 167368 194488 167420 194540
rect 147772 194420 147824 194472
rect 148232 194420 148284 194472
rect 130384 194352 130436 194404
rect 147680 194352 147732 194404
rect 173164 194352 173216 194404
rect 207204 194352 207256 194404
rect 108672 194284 108724 194336
rect 140688 194284 140740 194336
rect 175096 194284 175148 194336
rect 208676 194284 208728 194336
rect 109684 194216 109736 194268
rect 108304 194148 108356 194200
rect 140320 194148 140372 194200
rect 147956 194216 148008 194268
rect 148600 194216 148652 194268
rect 175740 194216 175792 194268
rect 210148 194216 210200 194268
rect 141884 194148 141936 194200
rect 179880 194148 179932 194200
rect 207388 194148 207440 194200
rect 100484 194080 100536 194132
rect 126980 194080 127032 194132
rect 174084 194080 174136 194132
rect 208768 194080 208820 194132
rect 103336 194012 103388 194064
rect 135536 194012 135588 194064
rect 158996 194012 159048 194064
rect 176016 194012 176068 194064
rect 177028 194012 177080 194064
rect 177580 194012 177632 194064
rect 179420 194012 179472 194064
rect 211804 194012 211856 194064
rect 108764 193944 108816 193996
rect 143172 193944 143224 193996
rect 158812 193944 158864 193996
rect 159548 193944 159600 193996
rect 162124 193944 162176 193996
rect 174820 193944 174872 193996
rect 175464 193944 175516 193996
rect 210516 193944 210568 193996
rect 104348 193876 104400 193928
rect 139308 193876 139360 193928
rect 151820 193876 151872 193928
rect 171600 193876 171652 193928
rect 174544 193876 174596 193928
rect 214380 193876 214432 193928
rect 96436 193808 96488 193860
rect 135996 193808 136048 193860
rect 141332 193808 141384 193860
rect 143908 193808 143960 193860
rect 169576 193808 169628 193860
rect 221372 193808 221424 193860
rect 156512 193332 156564 193384
rect 157248 193332 157300 193384
rect 119528 193128 119580 193180
rect 143724 193128 143776 193180
rect 157708 193128 157760 193180
rect 158260 193128 158312 193180
rect 166816 193128 166868 193180
rect 200212 193128 200264 193180
rect 119436 193060 119488 193112
rect 145288 193060 145340 193112
rect 163136 193060 163188 193112
rect 163964 193060 164016 193112
rect 167460 193060 167512 193112
rect 201684 193060 201736 193112
rect 123944 192992 123996 193044
rect 153200 192992 153252 193044
rect 170404 192992 170456 193044
rect 204260 192992 204312 193044
rect 112720 192924 112772 192976
rect 146208 192924 146260 192976
rect 153292 192924 153344 192976
rect 153476 192924 153528 192976
rect 169208 192924 169260 192976
rect 203064 192924 203116 192976
rect 101680 192856 101732 192908
rect 135168 192856 135220 192908
rect 169944 192856 169996 192908
rect 204444 192856 204496 192908
rect 101772 192788 101824 192840
rect 134984 192788 135036 192840
rect 171508 192788 171560 192840
rect 205640 192788 205692 192840
rect 108580 192720 108632 192772
rect 142804 192720 142856 192772
rect 170128 192720 170180 192772
rect 204352 192720 204404 192772
rect 108212 192652 108264 192704
rect 142620 192652 142672 192704
rect 170680 192652 170732 192704
rect 204536 192652 204588 192704
rect 112260 192584 112312 192636
rect 146576 192584 146628 192636
rect 172152 192584 172204 192636
rect 205824 192584 205876 192636
rect 97816 192516 97868 192568
rect 143816 192516 143868 192568
rect 162492 192516 162544 192568
rect 171968 192516 172020 192568
rect 172980 192516 173032 192568
rect 207480 192516 207532 192568
rect 97448 192448 97500 192500
rect 150532 192448 150584 192500
rect 155224 192448 155276 192500
rect 216864 192448 216916 192500
rect 129372 192380 129424 192432
rect 150256 192380 150308 192432
rect 164976 192380 165028 192432
rect 174544 192380 174596 192432
rect 174636 192380 174688 192432
rect 202420 192380 202472 192432
rect 130476 192312 130528 192364
rect 149152 192312 149204 192364
rect 171784 192312 171836 192364
rect 183192 192312 183244 192364
rect 130752 192244 130804 192296
rect 147496 192244 147548 192296
rect 108856 191564 108908 191616
rect 141056 191564 141108 191616
rect 104808 191496 104860 191548
rect 137652 191496 137704 191548
rect 153292 191496 153344 191548
rect 154304 191496 154356 191548
rect 107476 191428 107528 191480
rect 139492 191428 139544 191480
rect 116768 191360 116820 191412
rect 149796 191360 149848 191412
rect 99196 191292 99248 191344
rect 132776 191292 132828 191344
rect 160836 191292 160888 191344
rect 167092 191292 167144 191344
rect 103060 191224 103112 191276
rect 137468 191224 137520 191276
rect 167184 191224 167236 191276
rect 168012 191224 168064 191276
rect 171416 191224 171468 191276
rect 172244 191224 172296 191276
rect 175556 191224 175608 191276
rect 176384 191224 176436 191276
rect 188344 191292 188396 191344
rect 201500 191224 201552 191276
rect 99104 191156 99156 191208
rect 146760 191156 146812 191208
rect 166356 191156 166408 191208
rect 200488 191156 200540 191208
rect 99012 191088 99064 191140
rect 133052 191020 133104 191072
rect 133788 191020 133840 191072
rect 135720 191020 135772 191072
rect 136088 191020 136140 191072
rect 138388 191088 138440 191140
rect 139216 191088 139268 191140
rect 140228 191088 140280 191140
rect 140596 191088 140648 191140
rect 163228 191088 163280 191140
rect 211620 191088 211672 191140
rect 146852 191020 146904 191072
rect 167828 191020 167880 191072
rect 168012 191020 168064 191072
rect 169760 191020 169812 191072
rect 170864 191020 170916 191072
rect 171140 191020 171192 191072
rect 171692 191020 171744 191072
rect 172612 191020 172664 191072
rect 173624 191020 173676 191072
rect 175464 191020 175516 191072
rect 176108 191020 176160 191072
rect 167092 190952 167144 191004
rect 168104 190952 168156 191004
rect 142620 190884 142672 190936
rect 142988 190884 143040 190936
rect 167644 190884 167696 190936
rect 168288 190884 168340 190936
rect 174176 190884 174228 190936
rect 174728 190884 174780 190936
rect 132132 190680 132184 190732
rect 132132 190476 132184 190528
rect 155500 190408 155552 190460
rect 185676 190408 185728 190460
rect 132040 190340 132092 190392
rect 132224 190340 132276 190392
rect 132316 190340 132368 190392
rect 132500 190340 132552 190392
rect 173716 190340 173768 190392
rect 205732 190340 205784 190392
rect 120816 190272 120868 190324
rect 151084 190272 151136 190324
rect 174452 190272 174504 190324
rect 208584 190272 208636 190324
rect 106096 190204 106148 190256
rect 137192 190204 137244 190256
rect 176476 190204 176528 190256
rect 210240 190204 210292 190256
rect 103244 190136 103296 190188
rect 136364 190136 136416 190188
rect 177304 190136 177356 190188
rect 211712 190136 211764 190188
rect 110144 190068 110196 190120
rect 144552 190068 144604 190120
rect 157892 190068 157944 190120
rect 202328 190068 202380 190120
rect 110052 190000 110104 190052
rect 144092 190000 144144 190052
rect 158996 190000 159048 190052
rect 207020 190000 207072 190052
rect 101864 189932 101916 189984
rect 135996 189932 136048 189984
rect 137284 189932 137336 189984
rect 137468 189932 137520 189984
rect 157800 189932 157852 189984
rect 219624 189932 219676 189984
rect 108120 189864 108172 189916
rect 143908 189864 143960 189916
rect 157984 189864 158036 189916
rect 221096 189864 221148 189916
rect 97356 189796 97408 189848
rect 144828 189796 144880 189848
rect 156512 189796 156564 189848
rect 221004 189796 221056 189848
rect 96344 189728 96396 189780
rect 149520 189728 149572 189780
rect 156420 189728 156472 189780
rect 221188 189728 221240 189780
rect 159640 189660 159692 189712
rect 185860 189660 185912 189712
rect 137192 188640 137244 188692
rect 137560 188640 137612 188692
rect 132224 188368 132276 188420
rect 132408 188368 132460 188420
rect 142528 188368 142580 188420
rect 143264 188368 143316 188420
rect 168564 188368 168616 188420
rect 168748 188368 168800 188420
rect 168472 188096 168524 188148
rect 169668 188096 169720 188148
rect 135720 187688 135772 187740
rect 136548 187688 136600 187740
rect 172520 187552 172572 187604
rect 173348 187552 173400 187604
rect 101956 187484 102008 187536
rect 135628 187484 135680 187536
rect 166172 187484 166224 187536
rect 212724 187484 212776 187536
rect 100300 187416 100352 187468
rect 133972 187416 134024 187468
rect 161940 187416 161992 187468
rect 210424 187416 210476 187468
rect 105912 187348 105964 187400
rect 139952 187348 140004 187400
rect 160468 187348 160520 187400
rect 208952 187348 209004 187400
rect 100392 187280 100444 187332
rect 134340 187280 134392 187332
rect 160376 187280 160428 187332
rect 208860 187280 208912 187332
rect 104440 187212 104492 187264
rect 138296 187212 138348 187264
rect 163872 187212 163924 187264
rect 215668 187212 215720 187264
rect 98920 187144 98972 187196
rect 133512 187144 133564 187196
rect 168196 187144 168248 187196
rect 219716 187144 219768 187196
rect 98736 187076 98788 187128
rect 133236 187076 133288 187128
rect 156328 187076 156380 187128
rect 210056 187076 210108 187128
rect 106924 187008 106976 187060
rect 141608 187008 141660 187060
rect 158904 187008 158956 187060
rect 218244 187008 218296 187060
rect 98828 186940 98880 186992
rect 145380 186940 145432 186992
rect 152372 186940 152424 186992
rect 217416 186940 217468 186992
rect 134248 186464 134300 186516
rect 135076 186464 135128 186516
rect 189816 165588 189868 165640
rect 580172 165588 580224 165640
rect 164792 158652 164844 158704
rect 197912 158652 197964 158704
rect 177120 158584 177172 158636
rect 210608 158584 210660 158636
rect 165988 158516 166040 158568
rect 201224 158516 201276 158568
rect 168748 158448 168800 158500
rect 203432 158448 203484 158500
rect 168012 158380 168064 158432
rect 216036 158380 216088 158432
rect 166080 158312 166132 158364
rect 217508 158312 217560 158364
rect 152372 158244 152424 158296
rect 204720 158244 204772 158296
rect 164700 158176 164752 158228
rect 219900 158176 219952 158228
rect 164608 158108 164660 158160
rect 219992 158108 220044 158160
rect 163136 158040 163188 158092
rect 219808 158040 219860 158092
rect 152280 157972 152332 158024
rect 218060 157972 218112 158024
rect 168840 157904 168892 157956
rect 198004 157904 198056 157956
rect 168932 157836 168984 157888
rect 196624 157836 196676 157888
rect 177212 157768 177264 157820
rect 203340 157768 203392 157820
rect 163044 155864 163096 155916
rect 184388 155864 184440 155916
rect 161848 155796 161900 155848
rect 184296 155796 184348 155848
rect 162952 155728 163004 155780
rect 186044 155728 186096 155780
rect 164332 155660 164384 155712
rect 188528 155660 188580 155712
rect 171508 155592 171560 155644
rect 200580 155592 200632 155644
rect 158812 155524 158864 155576
rect 188436 155524 188488 155576
rect 157708 155456 157760 155508
rect 188620 155456 188672 155508
rect 165896 155388 165948 155440
rect 200672 155388 200724 155440
rect 165804 155320 165856 155372
rect 200764 155320 200816 155372
rect 165712 155252 165764 155304
rect 211896 155252 211948 155304
rect 164516 155184 164568 155236
rect 213000 155184 213052 155236
rect 164424 155116 164476 155168
rect 184204 155116 184256 155168
rect 119344 154164 119396 154216
rect 133972 154164 134024 154216
rect 96252 154096 96304 154148
rect 134524 154096 134576 154148
rect 97172 154028 97224 154080
rect 140228 154028 140280 154080
rect 96160 153960 96212 154012
rect 140412 153960 140464 154012
rect 165712 153960 165764 154012
rect 203248 153960 203300 154012
rect 96988 153892 97040 153944
rect 145288 153892 145340 153944
rect 162952 153892 163004 153944
rect 204628 153892 204680 153944
rect 120908 153824 120960 153876
rect 170128 153824 170180 153876
rect 173716 153824 173768 153876
rect 214748 153824 214800 153876
rect 95884 153212 95936 153264
rect 184940 153212 184992 153264
rect 192576 153212 192628 153264
rect 158536 153144 158588 153196
rect 187332 153144 187384 153196
rect 156236 153076 156288 153128
rect 187148 153076 187200 153128
rect 157616 153008 157668 153060
rect 188712 153008 188764 153060
rect 160192 152940 160244 152992
rect 184664 152940 184716 152992
rect 186964 152940 187016 152992
rect 218428 152940 218480 152992
rect 175556 152872 175608 152924
rect 207940 152872 207992 152924
rect 176752 152804 176804 152856
rect 209136 152804 209188 152856
rect 176660 152736 176712 152788
rect 209044 152736 209096 152788
rect 157524 152668 157576 152720
rect 191380 152668 191432 152720
rect 160284 152600 160336 152652
rect 209228 152600 209280 152652
rect 158720 152532 158772 152584
rect 218336 152532 218388 152584
rect 111156 152464 111208 152516
rect 142896 152464 142948 152516
rect 154948 152464 155000 152516
rect 218612 152464 218664 152516
rect 157432 152396 157484 152448
rect 187240 152396 187292 152448
rect 183468 152328 183520 152380
rect 207664 152328 207716 152380
rect 187976 151784 188028 151836
rect 580080 151784 580132 151836
rect 114928 151716 114980 151768
rect 140964 151716 141016 151768
rect 101404 151648 101456 151700
rect 134248 151648 134300 151700
rect 102784 151580 102836 151632
rect 135812 151580 135864 151632
rect 98644 151512 98696 151564
rect 133052 151512 133104 151564
rect 102968 151444 103020 151496
rect 137376 151444 137428 151496
rect 100024 151376 100076 151428
rect 134340 151376 134392 151428
rect 174544 151376 174596 151428
rect 199476 151376 199528 151428
rect 100116 151308 100168 151360
rect 134064 151308 134116 151360
rect 171968 151308 172020 151360
rect 206008 151308 206060 151360
rect 101496 151240 101548 151292
rect 136088 151240 136140 151292
rect 168656 151240 168708 151292
rect 203524 151240 203576 151292
rect 98552 151172 98604 151224
rect 133144 151172 133196 151224
rect 167276 151172 167328 151224
rect 206100 151172 206152 151224
rect 101312 151104 101364 151156
rect 135536 151104 135588 151156
rect 154948 151104 155000 151156
rect 207572 151104 207624 151156
rect 96068 151036 96120 151088
rect 139308 151036 139360 151088
rect 153568 151036 153620 151088
rect 207112 151036 207164 151088
rect 118976 150968 119028 151020
rect 144920 150968 144972 151020
rect 124036 150900 124088 150952
rect 141884 150900 141936 150952
rect 125048 150424 125100 150476
rect 580540 150424 580592 150476
rect 182088 150356 182140 150408
rect 195060 150356 195112 150408
rect 171876 150288 171928 150340
rect 191288 150288 191340 150340
rect 175372 150220 175424 150272
rect 204904 150220 204956 150272
rect 172888 150152 172940 150204
rect 206192 150152 206244 150204
rect 174176 150084 174228 150136
rect 207572 150084 207624 150136
rect 172704 150016 172756 150068
rect 206284 150016 206336 150068
rect 173900 149948 173952 150000
rect 207756 149948 207808 150000
rect 173992 149880 174044 149932
rect 207664 149880 207716 149932
rect 171324 149812 171376 149864
rect 204996 149812 205048 149864
rect 175188 149744 175240 149796
rect 207848 149744 207900 149796
rect 99840 149676 99892 149728
rect 148048 149676 148100 149728
rect 171416 149676 171468 149728
rect 206100 149676 206152 149728
rect 3148 149132 3200 149184
rect 180892 149132 180944 149184
rect 182088 149132 182140 149184
rect 125692 149064 125744 149116
rect 126520 149064 126572 149116
rect 580632 149064 580684 149116
rect 118884 148996 118936 149048
rect 147036 148996 147088 149048
rect 171048 148996 171100 149048
rect 195060 148996 195112 149048
rect 104164 148928 104216 148980
rect 131948 148928 132000 148980
rect 161756 148928 161808 148980
rect 188804 148928 188856 148980
rect 110788 148860 110840 148912
rect 142528 148860 142580 148912
rect 162768 148860 162820 148912
rect 198372 148860 198424 148912
rect 122472 148792 122524 148844
rect 153476 148792 153528 148844
rect 161020 148792 161072 148844
rect 195612 148792 195664 148844
rect 111064 148724 111116 148776
rect 142620 148724 142672 148776
rect 161296 148724 161348 148776
rect 196900 148724 196952 148776
rect 98460 148656 98512 148708
rect 130660 148656 130712 148708
rect 164240 148656 164292 148708
rect 199752 148656 199804 148708
rect 118792 148588 118844 148640
rect 152188 148588 152240 148640
rect 168288 148588 168340 148640
rect 202052 148588 202104 148640
rect 99932 148520 99984 148572
rect 132316 148520 132368 148572
rect 169668 148520 169720 148572
rect 203708 148520 203760 148572
rect 114836 148452 114888 148504
rect 149336 148452 149388 148504
rect 160008 148452 160060 148504
rect 195152 148452 195204 148504
rect 97080 148384 97132 148436
rect 152096 148384 152148 148436
rect 165620 148384 165672 148436
rect 200856 148384 200908 148436
rect 112352 148316 112404 148368
rect 128912 148316 128964 148368
rect 187976 148316 188028 148368
rect 120908 148248 120960 148300
rect 147956 148248 148008 148300
rect 177672 148248 177724 148300
rect 199660 148248 199712 148300
rect 106740 148180 106792 148232
rect 131856 148180 131908 148232
rect 179604 147568 179656 147620
rect 196440 147568 196492 147620
rect 179788 147500 179840 147552
rect 199200 147500 199252 147552
rect 178592 147432 178644 147484
rect 199292 147432 199344 147484
rect 176660 147364 176712 147416
rect 197820 147364 197872 147416
rect 109592 147296 109644 147348
rect 138572 147296 138624 147348
rect 170036 147296 170088 147348
rect 195704 147296 195756 147348
rect 105360 147228 105412 147280
rect 137192 147228 137244 147280
rect 169852 147228 169904 147280
rect 199292 147228 199344 147280
rect 110696 147160 110748 147212
rect 144000 147160 144052 147212
rect 157340 147160 157392 147212
rect 182732 147160 182784 147212
rect 182916 147160 182968 147212
rect 183192 147160 183244 147212
rect 102876 147092 102928 147144
rect 135720 147092 135772 147144
rect 172520 147092 172572 147144
rect 104072 147024 104124 147076
rect 137284 147024 137336 147076
rect 156144 147024 156196 147076
rect 182640 147024 182692 147076
rect 206376 147092 206428 147144
rect 109408 146956 109460 147008
rect 143632 146956 143684 147008
rect 171140 146956 171192 147008
rect 205088 146956 205140 147008
rect 105452 146888 105504 146940
rect 140136 146888 140188 146940
rect 161388 146888 161440 146940
rect 197912 146888 197964 146940
rect 179512 146820 179564 146872
rect 197360 146820 197412 146872
rect 181536 146752 181588 146804
rect 190092 146752 190144 146804
rect 182732 146684 182784 146736
rect 189724 146684 189776 146736
rect 182640 146616 182692 146668
rect 190000 146616 190052 146668
rect 113824 146208 113876 146260
rect 129740 146208 129792 146260
rect 180156 146208 180208 146260
rect 193588 146208 193640 146260
rect 112628 146140 112680 146192
rect 130016 146140 130068 146192
rect 178132 146140 178184 146192
rect 193956 146140 194008 146192
rect 110972 146072 111024 146124
rect 132224 146072 132276 146124
rect 178040 146072 178092 146124
rect 194968 146072 195020 146124
rect 119896 146004 119948 146056
rect 149244 146004 149296 146056
rect 167920 146004 167972 146056
rect 194232 146004 194284 146056
rect 111432 145936 111484 145988
rect 142160 145936 142212 145988
rect 165528 145936 165580 145988
rect 192576 145936 192628 145988
rect 116400 145868 116452 145920
rect 149060 145868 149112 145920
rect 161664 145868 161716 145920
rect 196992 145868 197044 145920
rect 116216 145800 116268 145852
rect 149704 145800 149756 145852
rect 157616 145800 157668 145852
rect 192208 145800 192260 145852
rect 117780 145732 117832 145784
rect 151820 145732 151872 145784
rect 161572 145732 161624 145784
rect 197084 145732 197136 145784
rect 116308 145664 116360 145716
rect 150716 145664 150768 145716
rect 157248 145664 157300 145716
rect 192208 145664 192260 145716
rect 113824 145596 113876 145648
rect 148416 145596 148468 145648
rect 150348 145596 150400 145648
rect 190184 145596 190236 145648
rect 3516 145528 3568 145580
rect 116492 145460 116544 145512
rect 130108 145460 130160 145512
rect 179420 145528 179472 145580
rect 196532 145528 196584 145580
rect 179696 145460 179748 145512
rect 189632 145460 189684 145512
rect 115480 144848 115532 144900
rect 135352 144848 135404 144900
rect 174360 144848 174412 144900
rect 196256 144848 196308 144900
rect 114192 144780 114244 144832
rect 136180 144780 136232 144832
rect 168472 144780 168524 144832
rect 194508 144780 194560 144832
rect 110880 144712 110932 144764
rect 132040 144712 132092 144764
rect 171048 144712 171100 144764
rect 196164 144712 196216 144764
rect 115296 144644 115348 144696
rect 138020 144644 138072 144696
rect 165804 144644 165856 144696
rect 192392 144644 192444 144696
rect 111524 144576 111576 144628
rect 137284 144576 137336 144628
rect 156696 144576 156748 144628
rect 189356 144576 189408 144628
rect 119988 144508 120040 144560
rect 147772 144508 147824 144560
rect 159456 144508 159508 144560
rect 192484 144508 192536 144560
rect 109776 144440 109828 144492
rect 138940 144440 138992 144492
rect 155684 144440 155736 144492
rect 189080 144440 189132 144492
rect 119712 144372 119764 144424
rect 150532 144372 150584 144424
rect 155868 144372 155920 144424
rect 191472 144372 191524 144424
rect 112536 144304 112588 144356
rect 143908 144304 143960 144356
rect 160008 144304 160060 144356
rect 193772 144304 193824 144356
rect 119344 144236 119396 144288
rect 129188 144236 129240 144288
rect 130292 144236 130344 144288
rect 189816 144236 189868 144288
rect 124956 144168 125008 144220
rect 131488 144168 131540 144220
rect 580356 144168 580408 144220
rect 117688 144100 117740 144152
rect 127900 144100 127952 144152
rect 175924 144100 175976 144152
rect 194876 144100 194928 144152
rect 113732 144032 113784 144084
rect 130292 144032 130344 144084
rect 180248 144032 180300 144084
rect 189356 144032 189408 144084
rect 185860 143760 185912 143812
rect 192392 143760 192444 143812
rect 115388 143488 115440 143540
rect 124220 143488 124272 143540
rect 174912 143488 174964 143540
rect 179512 143488 179564 143540
rect 185676 143488 185728 143540
rect 189632 143488 189684 143540
rect 124864 143420 124916 143472
rect 132868 143420 132920 143472
rect 176568 143420 176620 143472
rect 178592 143420 178644 143472
rect 186228 143420 186280 143472
rect 187792 143420 187844 143472
rect 118148 143352 118200 143404
rect 127440 143352 127492 143404
rect 177488 143352 177540 143404
rect 179420 143352 179472 143404
rect 116860 143284 116912 143336
rect 128728 143284 128780 143336
rect 171416 143284 171468 143336
rect 179788 143284 179840 143336
rect 114192 143216 114244 143268
rect 129280 143216 129332 143268
rect 185584 143216 185636 143268
rect 196348 143216 196400 143268
rect 118056 143148 118108 143200
rect 131764 143148 131816 143200
rect 131856 143148 131908 143200
rect 141148 143148 141200 143200
rect 165528 143148 165580 143200
rect 189540 143148 189592 143200
rect 113916 143080 113968 143132
rect 133420 143080 133472 143132
rect 160560 143080 160612 143132
rect 190736 143080 190788 143132
rect 117964 143012 118016 143064
rect 141700 143012 141752 143064
rect 156052 143012 156104 143064
rect 191840 143012 191892 143064
rect 116676 142944 116728 142996
rect 140044 142944 140096 142996
rect 154856 142944 154908 142996
rect 191104 142944 191156 142996
rect 115204 142876 115256 142928
rect 140780 142876 140832 142928
rect 168380 142876 168432 142928
rect 211988 142876 212040 142928
rect 116584 142808 116636 142860
rect 143540 142808 143592 142860
rect 150624 142808 150676 142860
rect 213092 142808 213144 142860
rect 183468 142672 183520 142724
rect 184480 142672 184532 142724
rect 128728 142468 128780 142520
rect 137008 142468 137060 142520
rect 184848 142468 184900 142520
rect 190828 142468 190880 142520
rect 129924 142400 129976 142452
rect 133512 142400 133564 142452
rect 120632 142332 120684 142384
rect 186228 142332 186280 142384
rect 128084 142264 128136 142316
rect 549904 142264 549956 142316
rect 130108 142196 130160 142248
rect 127992 142128 128044 142180
rect 129832 142128 129884 142180
rect 130016 142128 130068 142180
rect 132500 142128 132552 142180
rect 133512 142196 133564 142248
rect 579804 142196 579856 142248
rect 134524 142128 134576 142180
rect 137008 142128 137060 142180
rect 580816 142128 580868 142180
rect 112812 142060 112864 142112
rect 125508 142060 125560 142112
rect 182732 142060 182784 142112
rect 199108 142060 199160 142112
rect 112904 141992 112956 142044
rect 127532 141992 127584 142044
rect 176016 141992 176068 142044
rect 193956 141992 194008 142044
rect 115480 141924 115532 141976
rect 130476 141924 130528 141976
rect 173808 141924 173860 141976
rect 190644 141924 190696 141976
rect 114100 141856 114152 141908
rect 135628 141856 135680 141908
rect 175096 141856 175148 141908
rect 193864 141856 193916 141908
rect 115572 141788 115624 141840
rect 138388 141788 138440 141840
rect 168748 141788 168800 141840
rect 189264 141788 189316 141840
rect 112628 141720 112680 141772
rect 141608 141720 141660 141772
rect 166816 141720 166868 141772
rect 190920 141720 190972 141772
rect 116400 141652 116452 141704
rect 147220 141652 147272 141704
rect 156972 141652 157024 141704
rect 189908 141652 189960 141704
rect 115112 141584 115164 141636
rect 146852 141584 146904 141636
rect 157432 141584 157484 141636
rect 192300 141584 192352 141636
rect 116860 141516 116912 141568
rect 149612 141516 149664 141568
rect 154764 141516 154816 141568
rect 190828 141516 190880 141568
rect 113732 141448 113784 141500
rect 148232 141448 148284 141500
rect 163780 141448 163832 141500
rect 204628 141448 204680 141500
rect 112812 141380 112864 141432
rect 153660 141380 153712 141432
rect 154672 141380 154724 141432
rect 213184 141380 213236 141432
rect 118332 141312 118384 141364
rect 129372 141312 129424 141364
rect 179512 141312 179564 141364
rect 180616 141312 180668 141364
rect 193680 141312 193732 141364
rect 184296 141244 184348 141296
rect 196532 141244 196584 141296
rect 186044 141176 186096 141228
rect 198004 141176 198056 141228
rect 119068 140836 119120 140888
rect 179512 140836 179564 140888
rect 8944 140768 8996 140820
rect 183192 140768 183244 140820
rect 129740 140700 129792 140752
rect 130660 140700 130712 140752
rect 142160 140700 142212 140752
rect 142804 140700 142856 140752
rect 149244 140700 149296 140752
rect 149520 140700 149572 140752
rect 151820 140700 151872 140752
rect 152740 140700 152792 140752
rect 157340 140700 157392 140752
rect 158260 140700 158312 140752
rect 167000 140700 167052 140752
rect 167644 140700 167696 140752
rect 168840 140700 168892 140752
rect 169300 140700 169352 140752
rect 169760 140700 169812 140752
rect 193680 140700 193732 140752
rect 117964 140632 118016 140684
rect 127716 140632 127768 140684
rect 176660 140632 176712 140684
rect 177580 140632 177632 140684
rect 178040 140632 178092 140684
rect 178684 140632 178736 140684
rect 118056 140564 118108 140616
rect 127808 140564 127860 140616
rect 112904 140496 112956 140548
rect 123392 140496 123444 140548
rect 117872 140428 117924 140480
rect 129096 140428 129148 140480
rect 116676 140360 116728 140412
rect 129004 140360 129056 140412
rect 114100 140292 114152 140344
rect 130384 140292 130436 140344
rect 180064 140292 180116 140344
rect 189172 140292 189224 140344
rect 120724 140224 120776 140276
rect 151176 140224 151228 140276
rect 183100 140224 183152 140276
rect 193772 140224 193824 140276
rect 115296 140156 115348 140208
rect 148140 140156 148192 140208
rect 176200 140156 176252 140208
rect 188160 140156 188212 140208
rect 188712 140156 188764 140208
rect 191012 140156 191064 140208
rect 117780 140088 117832 140140
rect 151268 140088 151320 140140
rect 155776 140088 155828 140140
rect 178592 140088 178644 140140
rect 206008 140088 206060 140140
rect 104256 140020 104308 140072
rect 138296 140020 138348 140072
rect 119252 139952 119304 140004
rect 126428 139952 126480 140004
rect 190000 140020 190052 140072
rect 190920 140020 190972 140072
rect 191196 139952 191248 140004
rect 125692 139884 125744 139936
rect 126336 139884 126388 139936
rect 187332 139884 187384 139936
rect 192300 139884 192352 139936
rect 187148 139816 187200 139868
rect 189448 139816 189500 139868
rect 187240 139748 187292 139800
rect 192852 139816 192904 139868
rect 173256 139680 173308 139732
rect 199016 139680 199068 139732
rect 161480 139612 161532 139664
rect 194784 139612 194836 139664
rect 95976 139544 96028 139596
rect 182180 139544 182232 139596
rect 4804 139476 4856 139528
rect 180800 139476 180852 139528
rect 181444 139476 181496 139528
rect 182640 139476 182692 139528
rect 192116 139476 192168 139528
rect 113640 139408 113692 139460
rect 122196 139408 122248 139460
rect 126152 139408 126204 139460
rect 327724 139408 327776 139460
rect 184664 139340 184716 139392
rect 186504 139340 186556 139392
rect 188436 139272 188488 139324
rect 192484 139272 192536 139324
rect 188252 138864 188304 138916
rect 195336 138864 195388 138916
rect 188804 138796 188856 138848
rect 196440 138796 196492 138848
rect 188528 138728 188580 138780
rect 199384 138728 199436 138780
rect 3424 138660 3476 138712
rect 120632 138660 120684 138712
rect 188160 138660 188212 138712
rect 203616 138660 203668 138712
rect 191288 138116 191340 138168
rect 198188 138116 198240 138168
rect 188620 137980 188672 138032
rect 190000 137980 190052 138032
rect 3240 137912 3292 137964
rect 119068 137912 119120 137964
rect 188160 137776 188212 137828
rect 202144 137776 202196 137828
rect 188896 136688 188948 136740
rect 202236 136688 202288 136740
rect 202328 136552 202380 136604
rect 206468 136552 206520 136604
rect 195428 124856 195480 124908
rect 204812 124856 204864 124908
rect 192576 122068 192628 122120
rect 202328 122068 202380 122120
rect 191196 118668 191248 118720
rect 191932 118668 191984 118720
rect 189724 114520 189776 114572
rect 191104 114520 191156 114572
rect 190000 114384 190052 114436
rect 192576 114384 192628 114436
rect 189908 113840 189960 113892
rect 191196 113840 191248 113892
rect 189816 113704 189868 113756
rect 191932 113704 191984 113756
rect 2780 110780 2832 110832
rect 4804 110780 4856 110832
rect 115020 110440 115072 110492
rect 120724 110440 120776 110492
rect 549904 100648 549956 100700
rect 579620 100648 579672 100700
rect 105636 89088 105688 89140
rect 105728 88884 105780 88936
rect 482284 86912 482336 86964
rect 579620 86912 579672 86964
rect 197912 86776 197964 86828
rect 198004 86572 198056 86624
rect 3516 85484 3568 85536
rect 95976 85484 96028 85536
rect 188896 82764 188948 82816
rect 203708 82764 203760 82816
rect 188988 82084 189040 82136
rect 196164 82084 196216 82136
rect 215852 81064 215904 81116
rect 216128 81064 216180 81116
rect 114928 80996 114980 81048
rect 120724 80996 120776 81048
rect 109500 80860 109552 80912
rect 120816 80860 120868 80912
rect 105176 80792 105228 80844
rect 120080 80792 120132 80844
rect 121000 80792 121052 80844
rect 112444 80724 112496 80776
rect 112352 80656 112404 80708
rect 118700 80588 118752 80640
rect 121092 80520 121144 80572
rect 121184 80452 121236 80504
rect 102784 80384 102836 80436
rect 124864 80384 124916 80436
rect 131948 80384 132000 80436
rect 131764 80316 131816 80368
rect 131672 80112 131724 80164
rect 130384 80044 130436 80096
rect 130476 79976 130528 80028
rect 133006 79908 133058 79960
rect 132638 79840 132690 79892
rect 133650 79908 133702 79960
rect 134110 79908 134162 79960
rect 133282 79840 133334 79892
rect 133374 79840 133426 79892
rect 133466 79840 133518 79892
rect 113732 79772 113784 79824
rect 99840 79704 99892 79756
rect 132316 79704 132368 79756
rect 120540 79636 120592 79688
rect 130568 79636 130620 79688
rect 131028 79636 131080 79688
rect 133098 79772 133150 79824
rect 132592 79704 132644 79756
rect 132776 79636 132828 79688
rect 109684 79568 109736 79620
rect 123760 79568 123812 79620
rect 127072 79568 127124 79620
rect 132960 79636 133012 79688
rect 133052 79636 133104 79688
rect 133512 79636 133564 79688
rect 133420 79568 133472 79620
rect 106924 79500 106976 79552
rect 122840 79500 122892 79552
rect 124128 79500 124180 79552
rect 128636 79500 128688 79552
rect 133144 79500 133196 79552
rect 108028 79432 108080 79484
rect 108672 79432 108724 79484
rect 113640 79432 113692 79484
rect 108396 79364 108448 79416
rect 126980 79364 127032 79416
rect 132500 79432 132552 79484
rect 133834 79840 133886 79892
rect 133926 79840 133978 79892
rect 133880 79704 133932 79756
rect 133788 79636 133840 79688
rect 133972 79568 134024 79620
rect 134478 79908 134530 79960
rect 134846 79908 134898 79960
rect 134938 79908 134990 79960
rect 134662 79840 134714 79892
rect 136042 79908 136094 79960
rect 135674 79840 135726 79892
rect 135766 79840 135818 79892
rect 135214 79772 135266 79824
rect 135398 79772 135450 79824
rect 135490 79772 135542 79824
rect 134892 79636 134944 79688
rect 135076 79636 135128 79688
rect 135536 79636 135588 79688
rect 134524 79568 134576 79620
rect 134616 79568 134668 79620
rect 135168 79568 135220 79620
rect 135352 79568 135404 79620
rect 134800 79500 134852 79552
rect 130844 79364 130896 79416
rect 131028 79364 131080 79416
rect 96068 79296 96120 79348
rect 108212 79296 108264 79348
rect 131212 79296 131264 79348
rect 132316 79296 132368 79348
rect 132776 79364 132828 79416
rect 134248 79364 134300 79416
rect 135444 79364 135496 79416
rect 135858 79772 135910 79824
rect 135812 79568 135864 79620
rect 136594 79908 136646 79960
rect 136870 79908 136922 79960
rect 137330 79908 137382 79960
rect 136410 79840 136462 79892
rect 136502 79840 136554 79892
rect 136456 79704 136508 79756
rect 136180 79500 136232 79552
rect 135996 79432 136048 79484
rect 136456 79432 136508 79484
rect 137054 79840 137106 79892
rect 137606 79908 137658 79960
rect 137974 79908 138026 79960
rect 138066 79908 138118 79960
rect 138526 79908 138578 79960
rect 136916 79772 136968 79824
rect 137100 79704 137152 79756
rect 137008 79636 137060 79688
rect 137422 79840 137474 79892
rect 137928 79704 137980 79756
rect 137560 79636 137612 79688
rect 138250 79840 138302 79892
rect 138112 79636 138164 79688
rect 137836 79500 137888 79552
rect 138572 79568 138624 79620
rect 138388 79432 138440 79484
rect 138894 79908 138946 79960
rect 138986 79908 139038 79960
rect 139170 79908 139222 79960
rect 139262 79908 139314 79960
rect 139124 79636 139176 79688
rect 139722 79908 139774 79960
rect 139814 79908 139866 79960
rect 139768 79704 139820 79756
rect 139998 79908 140050 79960
rect 140090 79840 140142 79892
rect 140274 79840 140326 79892
rect 139032 79500 139084 79552
rect 139952 79636 140004 79688
rect 139400 79568 139452 79620
rect 139308 79432 139360 79484
rect 139676 79500 139728 79552
rect 140458 79908 140510 79960
rect 140550 79908 140602 79960
rect 140642 79908 140694 79960
rect 140826 79908 140878 79960
rect 140320 79704 140372 79756
rect 140412 79704 140464 79756
rect 140688 79636 140740 79688
rect 141010 79840 141062 79892
rect 139860 79432 139912 79484
rect 140228 79432 140280 79484
rect 140872 79568 140924 79620
rect 141562 79908 141614 79960
rect 141746 79908 141798 79960
rect 141838 79908 141890 79960
rect 141930 79908 141982 79960
rect 142206 79908 142258 79960
rect 141286 79840 141338 79892
rect 141608 79636 141660 79688
rect 142114 79840 142166 79892
rect 142482 79840 142534 79892
rect 142574 79840 142626 79892
rect 141700 79568 141752 79620
rect 142252 79636 142304 79688
rect 142160 79568 142212 79620
rect 142620 79704 142672 79756
rect 141148 79500 141200 79552
rect 141240 79500 141292 79552
rect 141792 79500 141844 79552
rect 140596 79432 140648 79484
rect 141424 79432 141476 79484
rect 141516 79432 141568 79484
rect 142528 79432 142580 79484
rect 143126 79908 143178 79960
rect 143218 79908 143270 79960
rect 143402 79908 143454 79960
rect 143494 79908 143546 79960
rect 143264 79704 143316 79756
rect 143356 79636 143408 79688
rect 143080 79568 143132 79620
rect 143632 79500 143684 79552
rect 144414 79908 144466 79960
rect 144506 79908 144558 79960
rect 143862 79840 143914 79892
rect 143954 79840 144006 79892
rect 144138 79840 144190 79892
rect 144322 79840 144374 79892
rect 144092 79704 144144 79756
rect 144184 79636 144236 79688
rect 143816 79568 143868 79620
rect 144414 79772 144466 79824
rect 144874 79908 144926 79960
rect 145150 79908 145202 79960
rect 145242 79908 145294 79960
rect 145334 79908 145386 79960
rect 144598 79840 144650 79892
rect 144690 79840 144742 79892
rect 144460 79636 144512 79688
rect 143908 79500 143960 79552
rect 136916 79364 136968 79416
rect 142712 79364 142764 79416
rect 142804 79364 142856 79416
rect 142896 79364 142948 79416
rect 144552 79364 144604 79416
rect 145196 79704 145248 79756
rect 145380 79636 145432 79688
rect 145610 79908 145662 79960
rect 145886 79908 145938 79960
rect 145978 79908 146030 79960
rect 146346 79908 146398 79960
rect 146438 79908 146490 79960
rect 146622 79908 146674 79960
rect 146714 79908 146766 79960
rect 146806 79908 146858 79960
rect 146990 79908 147042 79960
rect 147082 79908 147134 79960
rect 147174 79908 147226 79960
rect 145794 79840 145846 79892
rect 145656 79500 145708 79552
rect 145472 79432 145524 79484
rect 145840 79704 145892 79756
rect 146070 79840 146122 79892
rect 146162 79840 146214 79892
rect 146116 79704 146168 79756
rect 145932 79636 145984 79688
rect 146208 79636 146260 79688
rect 146530 79840 146582 79892
rect 146576 79636 146628 79688
rect 146668 79636 146720 79688
rect 146300 79568 146352 79620
rect 146392 79568 146444 79620
rect 146898 79772 146950 79824
rect 146760 79500 146812 79552
rect 146852 79432 146904 79484
rect 148094 79908 148146 79960
rect 149106 79908 149158 79960
rect 149290 79908 149342 79960
rect 149474 79908 149526 79960
rect 149566 79908 149618 79960
rect 149842 79908 149894 79960
rect 150026 79908 150078 79960
rect 150118 79908 150170 79960
rect 150670 79908 150722 79960
rect 150762 79908 150814 79960
rect 147542 79772 147594 79824
rect 148462 79840 148514 79892
rect 148830 79840 148882 79892
rect 148278 79772 148330 79824
rect 147496 79636 147548 79688
rect 147588 79636 147640 79688
rect 148048 79636 148100 79688
rect 147220 79568 147272 79620
rect 147864 79568 147916 79620
rect 148232 79568 148284 79620
rect 147404 79500 147456 79552
rect 145748 79364 145800 79416
rect 147036 79364 147088 79416
rect 149198 79772 149250 79824
rect 148968 79568 149020 79620
rect 149152 79568 149204 79620
rect 149244 79500 149296 79552
rect 149520 79772 149572 79824
rect 150072 79704 150124 79756
rect 149796 79500 149848 79552
rect 148508 79432 148560 79484
rect 149336 79432 149388 79484
rect 149612 79432 149664 79484
rect 148876 79364 148928 79416
rect 149428 79364 149480 79416
rect 150578 79840 150630 79892
rect 150532 79636 150584 79688
rect 150808 79568 150860 79620
rect 151084 79500 151136 79552
rect 151406 79908 151458 79960
rect 152142 79908 152194 79960
rect 152418 79908 152470 79960
rect 152510 79908 152562 79960
rect 153338 79908 153390 79960
rect 153430 79908 153482 79960
rect 153522 79908 153574 79960
rect 153798 79908 153850 79960
rect 154074 79908 154126 79960
rect 154166 79908 154218 79960
rect 154350 79908 154402 79960
rect 151590 79840 151642 79892
rect 151958 79840 152010 79892
rect 152234 79840 152286 79892
rect 151636 79704 151688 79756
rect 151544 79568 151596 79620
rect 152372 79704 152424 79756
rect 152970 79840 153022 79892
rect 153154 79840 153206 79892
rect 153246 79840 153298 79892
rect 152694 79772 152746 79824
rect 152188 79636 152240 79688
rect 152464 79636 152516 79688
rect 152648 79636 152700 79688
rect 152004 79568 152056 79620
rect 152832 79568 152884 79620
rect 151452 79500 151504 79552
rect 151360 79432 151412 79484
rect 151820 79432 151872 79484
rect 153384 79704 153436 79756
rect 153844 79704 153896 79756
rect 153476 79636 153528 79688
rect 153568 79636 153620 79688
rect 153936 79568 153988 79620
rect 153752 79500 153804 79552
rect 154304 79704 154356 79756
rect 205088 80792 205140 80844
rect 178224 80588 178276 80640
rect 213184 80724 213236 80776
rect 302240 80724 302292 80776
rect 177764 80452 177816 80504
rect 196716 80656 196768 80708
rect 380900 80656 380952 80708
rect 192484 80588 192536 80640
rect 177764 80316 177816 80368
rect 178316 80316 178368 80368
rect 191012 80520 191064 80572
rect 188344 80452 188396 80504
rect 192392 80452 192444 80504
rect 188436 80384 188488 80436
rect 195336 80384 195388 80436
rect 187056 80316 187108 80368
rect 195152 80316 195204 80368
rect 178408 80248 178460 80300
rect 154626 79908 154678 79960
rect 154488 79636 154540 79688
rect 154580 79568 154632 79620
rect 154212 79432 154264 79484
rect 154994 79908 155046 79960
rect 155086 79908 155138 79960
rect 155178 79908 155230 79960
rect 155454 79908 155506 79960
rect 155546 79908 155598 79960
rect 155730 79908 155782 79960
rect 155822 79908 155874 79960
rect 155914 79908 155966 79960
rect 158030 79908 158082 79960
rect 154902 79840 154954 79892
rect 155040 79500 155092 79552
rect 155408 79568 155460 79620
rect 155638 79772 155690 79824
rect 155224 79500 155276 79552
rect 155500 79500 155552 79552
rect 155316 79432 155368 79484
rect 156834 79840 156886 79892
rect 156926 79840 156978 79892
rect 157478 79840 157530 79892
rect 157846 79840 157898 79892
rect 156282 79772 156334 79824
rect 155868 79500 155920 79552
rect 155776 79432 155828 79484
rect 156972 79704 157024 79756
rect 156788 79568 156840 79620
rect 157616 79568 157668 79620
rect 156696 79500 156748 79552
rect 157432 79500 157484 79552
rect 158214 79908 158266 79960
rect 158306 79908 158358 79960
rect 158306 79772 158358 79824
rect 158260 79636 158312 79688
rect 158490 79908 158542 79960
rect 158582 79908 158634 79960
rect 158674 79908 158726 79960
rect 158628 79772 158680 79824
rect 159134 79908 159186 79960
rect 159226 79908 159278 79960
rect 159318 79908 159370 79960
rect 159502 79908 159554 79960
rect 159594 79908 159646 79960
rect 159962 79908 160014 79960
rect 160146 79908 160198 79960
rect 160514 79908 160566 79960
rect 158950 79772 159002 79824
rect 159042 79772 159094 79824
rect 159180 79772 159232 79824
rect 158720 79636 158772 79688
rect 158812 79636 158864 79688
rect 158168 79568 158220 79620
rect 158536 79568 158588 79620
rect 158076 79432 158128 79484
rect 158904 79568 158956 79620
rect 158904 79432 158956 79484
rect 154856 79364 154908 79416
rect 155132 79364 155184 79416
rect 159272 79704 159324 79756
rect 159778 79772 159830 79824
rect 159548 79704 159600 79756
rect 160606 79840 160658 79892
rect 160790 79840 160842 79892
rect 161066 79840 161118 79892
rect 160468 79772 160520 79824
rect 160560 79704 160612 79756
rect 159824 79636 159876 79688
rect 160100 79636 160152 79688
rect 161342 79840 161394 79892
rect 161986 79908 162038 79960
rect 162078 79908 162130 79960
rect 162170 79908 162222 79960
rect 162354 79908 162406 79960
rect 162446 79908 162498 79960
rect 162538 79908 162590 79960
rect 162722 79908 162774 79960
rect 163090 79908 163142 79960
rect 163274 79908 163326 79960
rect 163366 79908 163418 79960
rect 163458 79908 163510 79960
rect 161618 79840 161670 79892
rect 161710 79840 161762 79892
rect 161020 79568 161072 79620
rect 161204 79568 161256 79620
rect 161480 79568 161532 79620
rect 161848 79500 161900 79552
rect 162032 79772 162084 79824
rect 162308 79772 162360 79824
rect 162446 79772 162498 79824
rect 162124 79704 162176 79756
rect 162492 79636 162544 79688
rect 162998 79772 163050 79824
rect 162676 79568 162728 79620
rect 163136 79636 163188 79688
rect 163228 79636 163280 79688
rect 163320 79636 163372 79688
rect 163044 79568 163096 79620
rect 162492 79500 162544 79552
rect 162860 79500 162912 79552
rect 164378 79908 164430 79960
rect 164562 79908 164614 79960
rect 165022 79908 165074 79960
rect 165574 79908 165626 79960
rect 165758 79908 165810 79960
rect 165942 79908 165994 79960
rect 166034 79908 166086 79960
rect 163734 79840 163786 79892
rect 164102 79772 164154 79824
rect 164654 79840 164706 79892
rect 164516 79704 164568 79756
rect 164608 79704 164660 79756
rect 164332 79636 164384 79688
rect 164884 79636 164936 79688
rect 164056 79568 164108 79620
rect 161940 79432 161992 79484
rect 159548 79364 159600 79416
rect 160744 79364 160796 79416
rect 143172 79296 143224 79348
rect 164424 79364 164476 79416
rect 165206 79840 165258 79892
rect 165298 79772 165350 79824
rect 165390 79772 165442 79824
rect 165804 79704 165856 79756
rect 165436 79636 165488 79688
rect 165528 79636 165580 79688
rect 165344 79568 165396 79620
rect 166034 79772 166086 79824
rect 166310 79908 166362 79960
rect 166402 79908 166454 79960
rect 166494 79908 166546 79960
rect 166862 79908 166914 79960
rect 166448 79636 166500 79688
rect 178132 80180 178184 80232
rect 191288 80180 191340 80232
rect 191932 80180 191984 80232
rect 178040 80112 178092 80164
rect 167046 79908 167098 79960
rect 167000 79636 167052 79688
rect 166080 79568 166132 79620
rect 166172 79568 166224 79620
rect 166632 79568 166684 79620
rect 166908 79568 166960 79620
rect 166356 79500 166408 79552
rect 167092 79500 167144 79552
rect 167414 79908 167466 79960
rect 167506 79908 167558 79960
rect 168334 79908 168386 79960
rect 168426 79908 168478 79960
rect 168702 79908 168754 79960
rect 168978 79908 169030 79960
rect 169070 79908 169122 79960
rect 169162 79908 169214 79960
rect 167966 79840 168018 79892
rect 168150 79840 168202 79892
rect 168104 79704 168156 79756
rect 168012 79636 168064 79688
rect 168196 79636 168248 79688
rect 167920 79500 167972 79552
rect 167552 79432 167604 79484
rect 168518 79840 168570 79892
rect 168886 79840 168938 79892
rect 168656 79772 168708 79824
rect 168748 79772 168800 79824
rect 168840 79704 168892 79756
rect 168472 79568 168524 79620
rect 169254 79840 169306 79892
rect 169116 79704 169168 79756
rect 169208 79704 169260 79756
rect 169530 79908 169582 79960
rect 169714 79840 169766 79892
rect 169484 79704 169536 79756
rect 169392 79636 169444 79688
rect 167092 79364 167144 79416
rect 168932 79432 168984 79484
rect 169576 79500 169628 79552
rect 169898 79772 169950 79824
rect 169990 79772 170042 79824
rect 170174 79772 170226 79824
rect 170266 79772 170318 79824
rect 170036 79636 170088 79688
rect 169852 79568 169904 79620
rect 169944 79568 169996 79620
rect 170128 79568 170180 79620
rect 169760 79432 169812 79484
rect 170910 79908 170962 79960
rect 171278 79908 171330 79960
rect 171370 79908 171422 79960
rect 171554 79908 171606 79960
rect 171646 79908 171698 79960
rect 171830 79908 171882 79960
rect 171922 79908 171974 79960
rect 170726 79840 170778 79892
rect 170818 79840 170870 79892
rect 170864 79636 170916 79688
rect 170680 79568 170732 79620
rect 171416 79704 171468 79756
rect 171508 79704 171560 79756
rect 171738 79840 171790 79892
rect 171600 79636 171652 79688
rect 171232 79568 171284 79620
rect 172106 79908 172158 79960
rect 172290 79908 172342 79960
rect 172658 79908 172710 79960
rect 171968 79636 172020 79688
rect 172198 79840 172250 79892
rect 172750 79840 172802 79892
rect 174038 79908 174090 79960
rect 173026 79840 173078 79892
rect 172382 79772 172434 79824
rect 172566 79772 172618 79824
rect 173302 79772 173354 79824
rect 172244 79704 172296 79756
rect 171876 79568 171928 79620
rect 172060 79568 172112 79620
rect 172152 79568 172204 79620
rect 172612 79636 172664 79688
rect 173348 79636 173400 79688
rect 172428 79500 172480 79552
rect 169300 79364 169352 79416
rect 171140 79364 171192 79416
rect 171784 79364 171836 79416
rect 172888 79364 172940 79416
rect 172980 79364 173032 79416
rect 173256 79364 173308 79416
rect 173072 79296 173124 79348
rect 111340 79228 111392 79280
rect 145012 79228 145064 79280
rect 147864 79228 147916 79280
rect 172980 79228 173032 79280
rect 173946 79772 173998 79824
rect 173900 79636 173952 79688
rect 174222 79840 174274 79892
rect 174268 79636 174320 79688
rect 174498 79908 174550 79960
rect 174590 79908 174642 79960
rect 174682 79908 174734 79960
rect 174544 79772 174596 79824
rect 175326 79908 175378 79960
rect 178224 80044 178276 80096
rect 186964 80044 187016 80096
rect 190092 80044 190144 80096
rect 215852 80044 215904 80096
rect 288440 80044 288492 80096
rect 178776 79976 178828 80028
rect 175878 79908 175930 79960
rect 175970 79908 176022 79960
rect 176154 79908 176206 79960
rect 176338 79908 176390 79960
rect 176430 79908 176482 79960
rect 176890 79908 176942 79960
rect 177074 79908 177126 79960
rect 177764 79908 177816 79960
rect 175694 79840 175746 79892
rect 175510 79772 175562 79824
rect 174728 79636 174780 79688
rect 175188 79636 175240 79688
rect 175280 79636 175332 79688
rect 175464 79636 175516 79688
rect 175832 79704 175884 79756
rect 176614 79840 176666 79892
rect 176798 79840 176850 79892
rect 176016 79704 176068 79756
rect 176200 79704 176252 79756
rect 176384 79704 176436 79756
rect 176292 79636 176344 79688
rect 173532 79500 173584 79552
rect 175924 79568 175976 79620
rect 176108 79568 176160 79620
rect 177166 79840 177218 79892
rect 213092 79840 213144 79892
rect 238760 79840 238812 79892
rect 216772 79772 216824 79824
rect 217416 79772 217468 79824
rect 252560 79772 252612 79824
rect 177120 79704 177172 79756
rect 183744 79704 183796 79756
rect 219992 79704 220044 79756
rect 180432 79636 180484 79688
rect 217508 79636 217560 79688
rect 176936 79568 176988 79620
rect 177028 79568 177080 79620
rect 178960 79568 179012 79620
rect 216036 79568 216088 79620
rect 376760 79568 376812 79620
rect 176660 79500 176712 79552
rect 176844 79500 176896 79552
rect 212172 79500 212224 79552
rect 480260 79500 480312 79552
rect 173992 79432 174044 79484
rect 179420 79432 179472 79484
rect 201408 79432 201460 79484
rect 212908 79432 212960 79484
rect 500960 79432 501012 79484
rect 174912 79364 174964 79416
rect 197268 79364 197320 79416
rect 197360 79364 197412 79416
rect 211988 79364 212040 79416
rect 212172 79364 212224 79416
rect 213736 79364 213788 79416
rect 525800 79364 525852 79416
rect 174452 79296 174504 79348
rect 179512 79296 179564 79348
rect 191288 79296 191340 79348
rect 198188 79296 198240 79348
rect 523132 79296 523184 79348
rect 200028 79228 200080 79280
rect 221188 79228 221240 79280
rect 221372 79228 221424 79280
rect 116400 79160 116452 79212
rect 146852 79160 146904 79212
rect 96160 79092 96212 79144
rect 119804 79092 119856 79144
rect 147220 79092 147272 79144
rect 112536 79024 112588 79076
rect 146116 79024 146168 79076
rect 161940 79092 161992 79144
rect 164884 79092 164936 79144
rect 172520 79092 172572 79144
rect 173072 79160 173124 79212
rect 173992 79160 174044 79212
rect 174084 79160 174136 79212
rect 174544 79160 174596 79212
rect 207664 79160 207716 79212
rect 174452 79092 174504 79144
rect 174636 79092 174688 79144
rect 201316 79092 201368 79144
rect 115112 78956 115164 79008
rect 146300 78956 146352 79008
rect 162860 79024 162912 79076
rect 197912 79024 197964 79076
rect 163412 78956 163464 79008
rect 165252 78956 165304 79008
rect 170496 78956 170548 79008
rect 170772 78956 170824 79008
rect 173348 78956 173400 79008
rect 212816 78956 212868 79008
rect 213736 78956 213788 79008
rect 111248 78888 111300 78940
rect 145840 78888 145892 78940
rect 146024 78888 146076 78940
rect 156052 78888 156104 78940
rect 157064 78888 157116 78940
rect 157524 78888 157576 78940
rect 157892 78888 157944 78940
rect 161204 78888 161256 78940
rect 208952 78888 209004 78940
rect 124128 78820 124180 78872
rect 140596 78820 140648 78872
rect 150716 78820 150768 78872
rect 213092 78820 213144 78872
rect 134248 78752 134300 78804
rect 147864 78752 147916 78804
rect 152096 78752 152148 78804
rect 216772 78752 216824 78804
rect 130844 78684 130896 78736
rect 137008 78684 137060 78736
rect 99932 78616 99984 78668
rect 125508 78616 125560 78668
rect 134064 78616 134116 78668
rect 130292 78548 130344 78600
rect 132316 78548 132368 78600
rect 142436 78684 142488 78736
rect 155960 78684 156012 78736
rect 157248 78684 157300 78736
rect 159088 78684 159140 78736
rect 160100 78684 160152 78736
rect 162584 78684 162636 78736
rect 138480 78616 138532 78668
rect 138756 78616 138808 78668
rect 140228 78616 140280 78668
rect 140688 78616 140740 78668
rect 141240 78616 141292 78668
rect 141608 78616 141660 78668
rect 147036 78616 147088 78668
rect 147404 78616 147456 78668
rect 156052 78616 156104 78668
rect 156880 78616 156932 78668
rect 165988 78616 166040 78668
rect 166724 78616 166776 78668
rect 168012 78684 168064 78736
rect 179328 78684 179380 78736
rect 201316 78684 201368 78736
rect 539692 78684 539744 78736
rect 171876 78616 171928 78668
rect 172704 78616 172756 78668
rect 172888 78616 172940 78668
rect 172980 78616 173032 78668
rect 174912 78616 174964 78668
rect 176660 78616 176712 78668
rect 177212 78616 177264 78668
rect 156236 78548 156288 78600
rect 119436 78480 119488 78532
rect 145380 78480 145432 78532
rect 158904 78480 158956 78532
rect 159732 78480 159784 78532
rect 165436 78548 165488 78600
rect 215852 78548 215904 78600
rect 191564 78480 191616 78532
rect 191748 78480 191800 78532
rect 119528 78344 119580 78396
rect 133144 78412 133196 78464
rect 163044 78412 163096 78464
rect 167460 78412 167512 78464
rect 168104 78412 168156 78464
rect 197912 78412 197964 78464
rect 129464 78344 129516 78396
rect 142344 78344 142396 78396
rect 161020 78344 161072 78396
rect 168012 78344 168064 78396
rect 168656 78344 168708 78396
rect 168840 78344 168892 78396
rect 169668 78344 169720 78396
rect 199016 78344 199068 78396
rect 108304 78276 108356 78328
rect 131948 78276 132000 78328
rect 132224 78276 132276 78328
rect 137560 78276 137612 78328
rect 168748 78276 168800 78328
rect 169300 78276 169352 78328
rect 173900 78276 173952 78328
rect 174636 78276 174688 78328
rect 175372 78276 175424 78328
rect 178224 78276 178276 78328
rect 179328 78276 179380 78328
rect 202328 78276 202380 78328
rect 104532 78208 104584 78260
rect 127164 78208 127216 78260
rect 129648 78208 129700 78260
rect 142252 78208 142304 78260
rect 158812 78208 158864 78260
rect 159824 78208 159876 78260
rect 167920 78208 167972 78260
rect 169668 78208 169720 78260
rect 172520 78208 172572 78260
rect 183744 78208 183796 78260
rect 184204 78208 184256 78260
rect 107016 78140 107068 78192
rect 129832 78140 129884 78192
rect 130752 78140 130804 78192
rect 138204 78140 138256 78192
rect 139032 78140 139084 78192
rect 154948 78140 155000 78192
rect 165436 78140 165488 78192
rect 166448 78140 166500 78192
rect 180156 78140 180208 78192
rect 180432 78140 180484 78192
rect 180616 78140 180668 78192
rect 200488 78140 200540 78192
rect 104072 78072 104124 78124
rect 127716 78072 127768 78124
rect 101312 78004 101364 78056
rect 128268 78004 128320 78056
rect 131028 78004 131080 78056
rect 141792 78072 141844 78124
rect 157432 78072 157484 78124
rect 163044 78072 163096 78124
rect 163596 78072 163648 78124
rect 179236 78072 179288 78124
rect 168656 78004 168708 78056
rect 169392 78004 169444 78056
rect 46940 77936 46992 77988
rect 105636 77936 105688 77988
rect 106740 77936 106792 77988
rect 131304 77936 131356 77988
rect 131672 77936 131724 77988
rect 132316 77936 132368 77988
rect 141424 77936 141476 77988
rect 164332 77936 164384 77988
rect 178868 78004 178920 78056
rect 180708 78072 180760 78124
rect 202052 78072 202104 78124
rect 214748 78004 214800 78056
rect 215852 78004 215904 78056
rect 216128 78004 216180 78056
rect 270500 78004 270552 78056
rect 173900 77936 173952 77988
rect 174268 77936 174320 77988
rect 103152 77868 103204 77920
rect 124220 77868 124272 77920
rect 125508 77868 125560 77920
rect 133972 77868 134024 77920
rect 134616 77868 134668 77920
rect 109592 77800 109644 77852
rect 127624 77800 127676 77852
rect 130844 77800 130896 77852
rect 141884 77868 141936 77920
rect 166908 77868 166960 77920
rect 181628 77936 181680 77988
rect 182088 77936 182140 77988
rect 191748 77936 191800 77988
rect 306380 77936 306432 77988
rect 179328 77868 179380 77920
rect 198004 77868 198056 77920
rect 137008 77800 137060 77852
rect 144920 77800 144972 77852
rect 160468 77800 160520 77852
rect 162124 77800 162176 77852
rect 172520 77800 172572 77852
rect 172796 77800 172848 77852
rect 175924 77800 175976 77852
rect 177212 77800 177264 77852
rect 180432 77800 180484 77852
rect 195244 77800 195296 77852
rect 129556 77732 129608 77784
rect 142160 77732 142212 77784
rect 166356 77732 166408 77784
rect 180340 77732 180392 77784
rect 123760 77664 123812 77716
rect 141700 77664 141752 77716
rect 162492 77664 162544 77716
rect 178960 77664 179012 77716
rect 180064 77664 180116 77716
rect 194048 77664 194100 77716
rect 105728 77596 105780 77648
rect 137192 77596 137244 77648
rect 153476 77596 153528 77648
rect 215852 77596 215904 77648
rect 105636 77528 105688 77580
rect 135076 77528 135128 77580
rect 142252 77528 142304 77580
rect 142988 77528 143040 77580
rect 152464 77528 152516 77580
rect 152740 77528 152792 77580
rect 157156 77528 157208 77580
rect 162584 77528 162636 77580
rect 165804 77528 165856 77580
rect 126980 77460 127032 77512
rect 129648 77460 129700 77512
rect 130936 77460 130988 77512
rect 140044 77460 140096 77512
rect 142712 77460 142764 77512
rect 142896 77460 142948 77512
rect 161848 77460 161900 77512
rect 166908 77460 166960 77512
rect 167460 77528 167512 77580
rect 179328 77528 179380 77580
rect 180616 77460 180668 77512
rect 133144 77392 133196 77444
rect 143540 77392 143592 77444
rect 144000 77392 144052 77444
rect 144092 77324 144144 77376
rect 161480 77324 161532 77376
rect 161848 77324 161900 77376
rect 197912 77324 197964 77376
rect 287704 77324 287756 77376
rect 135720 77256 135772 77308
rect 136088 77256 136140 77308
rect 137008 77256 137060 77308
rect 137284 77256 137336 77308
rect 142620 77256 142672 77308
rect 143356 77256 143408 77308
rect 153476 77256 153528 77308
rect 153844 77256 153896 77308
rect 164240 77256 164292 77308
rect 165528 77256 165580 77308
rect 199016 77256 199068 77308
rect 453304 77256 453356 77308
rect 101220 77188 101272 77240
rect 99012 77120 99064 77172
rect 146392 77120 146444 77172
rect 96160 77052 96212 77104
rect 138572 77052 138624 77104
rect 114284 76984 114336 77036
rect 146576 76984 146628 77036
rect 111616 76916 111668 76968
rect 143356 76916 143408 76968
rect 105360 76848 105412 76900
rect 132224 76848 132276 76900
rect 134524 76848 134576 76900
rect 134800 76848 134852 76900
rect 144184 76848 144236 76900
rect 144368 76848 144420 76900
rect 115664 76780 115716 76832
rect 147036 76780 147088 76832
rect 114008 76712 114060 76764
rect 143448 76712 143500 76764
rect 116952 76644 117004 76696
rect 147312 76644 147364 76696
rect 96436 76576 96488 76628
rect 125600 76576 125652 76628
rect 128268 76576 128320 76628
rect 131396 76576 131448 76628
rect 135352 76576 135404 76628
rect 136640 76576 136692 76628
rect 137468 76576 137520 76628
rect 144920 76576 144972 76628
rect 146024 76576 146076 76628
rect 155408 77188 155460 77240
rect 218060 77188 218112 77240
rect 218336 77188 218388 77240
rect 155132 76984 155184 77036
rect 218428 77120 218480 77172
rect 157340 76916 157392 76968
rect 157708 76916 157760 76968
rect 159916 76916 159968 76968
rect 218888 77052 218940 77104
rect 164332 76984 164384 77036
rect 164792 76984 164844 77036
rect 164608 76916 164660 76968
rect 165528 76916 165580 76968
rect 153200 76848 153252 76900
rect 154304 76848 154356 76900
rect 154764 76848 154816 76900
rect 154948 76848 155000 76900
rect 160744 76848 160796 76900
rect 208860 76984 208912 77036
rect 167460 76916 167512 76968
rect 168196 76916 168248 76968
rect 171784 76916 171836 76968
rect 196164 76916 196216 76968
rect 168840 76848 168892 76900
rect 169208 76848 169260 76900
rect 173532 76848 173584 76900
rect 174268 76848 174320 76900
rect 175372 76848 175424 76900
rect 176568 76848 176620 76900
rect 177948 76848 178000 76900
rect 211804 76848 211856 76900
rect 157340 76780 157392 76832
rect 157984 76780 158036 76832
rect 168196 76780 168248 76832
rect 169668 76780 169720 76832
rect 201960 76780 202012 76832
rect 154764 76712 154816 76764
rect 155040 76712 155092 76764
rect 170220 76712 170272 76764
rect 171968 76712 172020 76764
rect 172612 76712 172664 76764
rect 173532 76712 173584 76764
rect 206284 76712 206336 76764
rect 218428 76712 218480 76764
rect 289820 76712 289872 76764
rect 148968 76644 149020 76696
rect 182824 76644 182876 76696
rect 218060 76644 218112 76696
rect 218612 76644 218664 76696
rect 296720 76644 296772 76696
rect 149244 76576 149296 76628
rect 150348 76576 150400 76628
rect 151452 76576 151504 76628
rect 198004 76576 198056 76628
rect 218888 76576 218940 76628
rect 353300 76576 353352 76628
rect 67640 76508 67692 76560
rect 105360 76508 105412 76560
rect 111248 76508 111300 76560
rect 113272 76440 113324 76492
rect 112628 76372 112680 76424
rect 129924 76372 129976 76424
rect 130844 76372 130896 76424
rect 125600 76304 125652 76356
rect 134432 76508 134484 76560
rect 134892 76508 134944 76560
rect 143356 76508 143408 76560
rect 146300 76508 146352 76560
rect 146576 76508 146628 76560
rect 182180 76508 182232 76560
rect 196164 76508 196216 76560
rect 196808 76508 196860 76560
rect 389180 76508 389232 76560
rect 145564 76440 145616 76492
rect 146024 76440 146076 76492
rect 147220 76440 147272 76492
rect 178684 76440 178736 76492
rect 140688 76372 140740 76424
rect 163688 76372 163740 76424
rect 171784 76372 171836 76424
rect 173440 76372 173492 76424
rect 173716 76372 173768 76424
rect 174176 76372 174228 76424
rect 177672 76372 177724 76424
rect 177856 76372 177908 76424
rect 199292 76372 199344 76424
rect 139676 76304 139728 76356
rect 145380 76304 145432 76356
rect 145564 76304 145616 76356
rect 152372 76304 152424 76356
rect 152832 76304 152884 76356
rect 170588 76304 170640 76356
rect 170772 76304 170824 76356
rect 176384 76304 176436 76356
rect 180432 76304 180484 76356
rect 170128 76236 170180 76288
rect 177856 76236 177908 76288
rect 131028 76168 131080 76220
rect 150624 76168 150676 76220
rect 150992 76168 151044 76220
rect 172704 76168 172756 76220
rect 173624 76168 173676 76220
rect 174176 76168 174228 76220
rect 175188 76168 175240 76220
rect 195704 76304 195756 76356
rect 163228 76100 163280 76152
rect 163412 76100 163464 76152
rect 170772 76100 170824 76152
rect 175832 76100 175884 76152
rect 176108 76100 176160 76152
rect 101312 76032 101364 76084
rect 101496 76032 101548 76084
rect 136640 76032 136692 76084
rect 137376 76032 137428 76084
rect 132776 75964 132828 76016
rect 133512 75964 133564 76016
rect 138020 75964 138072 76016
rect 138756 75964 138808 76016
rect 165988 75964 166040 76016
rect 166724 75964 166776 76016
rect 88984 75896 89036 75948
rect 96160 75896 96212 75948
rect 99932 75896 99984 75948
rect 100484 75896 100536 75948
rect 121460 75896 121512 75948
rect 123760 75896 123812 75948
rect 135536 75896 135588 75948
rect 136456 75896 136508 75948
rect 138480 75896 138532 75948
rect 138848 75896 138900 75948
rect 143448 75896 143500 75948
rect 145380 75896 145432 75948
rect 152464 75896 152516 75948
rect 160744 75896 160796 75948
rect 161388 75896 161440 75948
rect 164792 75896 164844 75948
rect 165068 75896 165120 75948
rect 168472 75896 168524 75948
rect 168840 75896 168892 75948
rect 172244 75896 172296 75948
rect 172428 75896 172480 75948
rect 176936 75896 176988 75948
rect 177948 75896 178000 75948
rect 97356 75828 97408 75880
rect 132040 75828 132092 75880
rect 137376 75828 137428 75880
rect 137744 75828 137796 75880
rect 158076 75828 158128 75880
rect 206468 75828 206520 75880
rect 98828 75760 98880 75812
rect 145840 75760 145892 75812
rect 163136 75760 163188 75812
rect 163320 75760 163372 75812
rect 170956 75760 171008 75812
rect 202236 75760 202288 75812
rect 202788 75760 202840 75812
rect 96068 75692 96120 75744
rect 99380 75692 99432 75744
rect 100484 75692 100536 75744
rect 104164 75692 104216 75744
rect 137836 75692 137888 75744
rect 172336 75692 172388 75744
rect 205548 75692 205600 75744
rect 206376 75692 206428 75744
rect 113088 75624 113140 75676
rect 147496 75624 147548 75676
rect 157892 75624 157944 75676
rect 89720 75420 89772 75472
rect 104348 75420 104400 75472
rect 139216 75556 139268 75608
rect 163320 75556 163372 75608
rect 163780 75556 163832 75608
rect 168748 75624 168800 75676
rect 169576 75624 169628 75676
rect 171876 75624 171928 75676
rect 206284 75624 206336 75676
rect 192300 75556 192352 75608
rect 119344 75488 119396 75540
rect 152280 75488 152332 75540
rect 152648 75488 152700 75540
rect 161480 75488 161532 75540
rect 162400 75488 162452 75540
rect 170864 75488 170916 75540
rect 204536 75488 204588 75540
rect 112996 75420 113048 75472
rect 145748 75420 145800 75472
rect 150900 75420 150952 75472
rect 151268 75420 151320 75472
rect 168748 75420 168800 75472
rect 169484 75420 169536 75472
rect 169852 75420 169904 75472
rect 171048 75420 171100 75472
rect 171416 75420 171468 75472
rect 172060 75420 172112 75472
rect 172796 75420 172848 75472
rect 173808 75420 173860 75472
rect 174636 75420 174688 75472
rect 207296 75420 207348 75472
rect 52460 75148 52512 75200
rect 100300 75352 100352 75404
rect 100484 75284 100536 75336
rect 107752 75352 107804 75404
rect 136548 75352 136600 75404
rect 150348 75352 150400 75404
rect 107016 75216 107068 75268
rect 107476 75216 107528 75268
rect 131120 75284 131172 75336
rect 133788 75284 133840 75336
rect 139952 75284 140004 75336
rect 140780 75284 140832 75336
rect 141976 75284 142028 75336
rect 150808 75284 150860 75336
rect 151268 75284 151320 75336
rect 158904 75352 158956 75404
rect 159456 75352 159508 75404
rect 160192 75352 160244 75404
rect 160928 75352 160980 75404
rect 178132 75352 178184 75404
rect 205916 75352 205968 75404
rect 216772 75284 216824 75336
rect 138296 75216 138348 75268
rect 138848 75216 138900 75268
rect 139768 75216 139820 75268
rect 140320 75216 140372 75268
rect 142896 75216 142948 75268
rect 143264 75216 143316 75268
rect 146668 75216 146720 75268
rect 176292 75216 176344 75268
rect 202788 75216 202840 75268
rect 454684 75216 454736 75268
rect 102876 75148 102928 75200
rect 107752 75148 107804 75200
rect 117136 75148 117188 75200
rect 145932 75148 145984 75200
rect 123116 75080 123168 75132
rect 108488 75012 108540 75064
rect 130016 75012 130068 75064
rect 137928 75012 137980 75064
rect 135996 74944 136048 74996
rect 136272 74944 136324 74996
rect 148048 75080 148100 75132
rect 176200 75148 176252 75200
rect 177304 75148 177356 75200
rect 201960 75148 202012 75200
rect 205916 75148 205968 75200
rect 499580 75148 499632 75200
rect 157432 75080 157484 75132
rect 158628 75080 158680 75132
rect 159088 75080 159140 75132
rect 159640 75080 159692 75132
rect 160192 75080 160244 75132
rect 160560 75080 160612 75132
rect 160652 75080 160704 75132
rect 161204 75080 161256 75132
rect 169024 75080 169076 75132
rect 176384 75080 176436 75132
rect 180340 75080 180392 75132
rect 219900 75080 219952 75132
rect 153752 74944 153804 74996
rect 146392 74808 146444 74860
rect 166724 75012 166776 75064
rect 172888 75012 172940 75064
rect 173808 75012 173860 75064
rect 176292 75012 176344 75064
rect 157892 74944 157944 74996
rect 158628 74944 158680 74996
rect 168472 74944 168524 74996
rect 169392 74944 169444 74996
rect 183560 75012 183612 75064
rect 184848 75012 184900 75064
rect 210608 75012 210660 75064
rect 185032 74944 185084 74996
rect 161204 74876 161256 74928
rect 169024 74876 169076 74928
rect 175556 74876 175608 74928
rect 176292 74876 176344 74928
rect 162308 74808 162360 74860
rect 162676 74808 162728 74860
rect 154672 74672 154724 74724
rect 155316 74672 155368 74724
rect 166724 74672 166776 74724
rect 180800 74672 180852 74724
rect 149704 74604 149756 74656
rect 150256 74604 150308 74656
rect 206284 74604 206336 74656
rect 475384 74604 475436 74656
rect 165712 74536 165764 74588
rect 166172 74536 166224 74588
rect 206376 74536 206428 74588
rect 511264 74536 511316 74588
rect 96344 74468 96396 74520
rect 149704 74468 149756 74520
rect 150072 74468 150124 74520
rect 153384 74468 153436 74520
rect 220820 74468 220872 74520
rect 114836 74400 114888 74452
rect 149980 74400 150032 74452
rect 159272 74400 159324 74452
rect 159916 74400 159968 74452
rect 161848 74400 161900 74452
rect 218244 74400 218296 74452
rect 122380 74332 122432 74384
rect 151544 74332 151596 74384
rect 155868 74332 155920 74384
rect 189816 74332 189868 74384
rect 98920 74264 98972 74316
rect 132960 74264 133012 74316
rect 166264 74264 166316 74316
rect 166908 74264 166960 74316
rect 200764 74264 200816 74316
rect 119252 74196 119304 74248
rect 151820 74196 151872 74248
rect 172428 74196 172480 74248
rect 206100 74196 206152 74248
rect 117964 74128 118016 74180
rect 150900 74128 150952 74180
rect 151636 74128 151688 74180
rect 155592 74128 155644 74180
rect 155868 74128 155920 74180
rect 171048 74128 171100 74180
rect 204444 74128 204496 74180
rect 101496 74060 101548 74112
rect 134984 74060 135036 74112
rect 173808 74060 173860 74112
rect 206192 74060 206244 74112
rect 116768 73992 116820 74044
rect 95976 73856 96028 73908
rect 107108 73856 107160 73908
rect 139400 73924 139452 73976
rect 159916 73992 159968 74044
rect 180064 73992 180116 74044
rect 181996 73992 182048 74044
rect 219716 73992 219768 74044
rect 220820 73992 220872 74044
rect 269120 73992 269172 74044
rect 163044 73924 163096 73976
rect 192208 73924 192260 73976
rect 322940 73924 322992 73976
rect 149888 73856 149940 73908
rect 207664 73856 207716 73908
rect 218244 73856 218296 73908
rect 354680 73856 354732 73908
rect 35900 73788 35952 73840
rect 101496 73788 101548 73840
rect 106280 73788 106332 73840
rect 136364 73788 136416 73840
rect 151544 73788 151596 73840
rect 248420 73788 248472 73840
rect 268384 73788 268436 73840
rect 581000 73788 581052 73840
rect 118056 73720 118108 73772
rect 141516 73720 141568 73772
rect 151820 73720 151872 73772
rect 152924 73720 152976 73772
rect 163044 73720 163096 73772
rect 164148 73720 164200 73772
rect 175188 73720 175240 73772
rect 207572 73720 207624 73772
rect 158076 73652 158128 73704
rect 158444 73652 158496 73704
rect 169208 73652 169260 73704
rect 179052 73652 179104 73704
rect 203156 73652 203208 73704
rect 97632 73584 97684 73636
rect 131488 73584 131540 73636
rect 132316 73584 132368 73636
rect 164056 73584 164108 73636
rect 166264 73584 166316 73636
rect 168288 73584 168340 73636
rect 181996 73584 182048 73636
rect 118516 73516 118568 73568
rect 149796 73516 149848 73568
rect 135812 73380 135864 73432
rect 136180 73380 136232 73432
rect 122104 73176 122156 73228
rect 122840 73176 122892 73228
rect 127716 73108 127768 73160
rect 136640 73108 136692 73160
rect 167644 73108 167696 73160
rect 168288 73108 168340 73160
rect 180708 73108 180760 73160
rect 327724 73108 327776 73160
rect 580172 73108 580224 73160
rect 115756 73040 115808 73092
rect 149152 73040 149204 73092
rect 149612 73040 149664 73092
rect 157800 73040 157852 73092
rect 221096 73040 221148 73092
rect 222108 73040 222160 73092
rect 129004 72972 129056 73024
rect 152832 72972 152884 73024
rect 161296 72972 161348 73024
rect 209228 72972 209280 73024
rect 114376 72904 114428 72956
rect 147864 72904 147916 72956
rect 148784 72904 148836 72956
rect 155776 72904 155828 72956
rect 190828 72904 190880 72956
rect 117228 72836 117280 72888
rect 149336 72836 149388 72888
rect 150164 72836 150216 72888
rect 166540 72836 166592 72888
rect 200948 72836 201000 72888
rect 115848 72768 115900 72820
rect 148140 72768 148192 72820
rect 148416 72768 148468 72820
rect 155224 72768 155276 72820
rect 189724 72768 189776 72820
rect 221372 72768 221424 72820
rect 311164 72768 311216 72820
rect 109868 72700 109920 72752
rect 142252 72700 142304 72752
rect 155776 72700 155828 72752
rect 189080 72700 189132 72752
rect 189632 72700 189684 72752
rect 283564 72700 283616 72752
rect 96620 72428 96672 72480
rect 107292 72428 107344 72480
rect 139124 72632 139176 72684
rect 145656 72632 145708 72684
rect 156880 72632 156932 72684
rect 162676 72632 162728 72684
rect 196532 72632 196584 72684
rect 222108 72632 222160 72684
rect 324964 72632 325016 72684
rect 117044 72564 117096 72616
rect 147956 72564 148008 72616
rect 148508 72564 148560 72616
rect 155684 72564 155736 72616
rect 118608 72496 118660 72548
rect 148048 72496 148100 72548
rect 148968 72496 149020 72548
rect 176936 72564 176988 72616
rect 177396 72564 177448 72616
rect 189080 72496 189132 72548
rect 111800 72428 111852 72480
rect 112444 72428 112496 72480
rect 140964 72428 141016 72480
rect 157064 72428 157116 72480
rect 191472 72564 191524 72616
rect 305000 72564 305052 72616
rect 110880 72360 110932 72412
rect 138204 72360 138256 72412
rect 160100 72360 160152 72412
rect 193956 72496 194008 72548
rect 340880 72496 340932 72548
rect 109960 72292 110012 72344
rect 128360 72292 128412 72344
rect 129464 72292 129516 72344
rect 162216 72292 162268 72344
rect 196624 72292 196676 72344
rect 382280 72428 382332 72480
rect 105544 72224 105596 72276
rect 140136 72224 140188 72276
rect 156604 72224 156656 72276
rect 221372 72224 221424 72276
rect 114192 72156 114244 72208
rect 148324 72156 148376 72208
rect 148508 72156 148560 72208
rect 156696 72156 156748 72208
rect 157248 72156 157300 72208
rect 190920 72156 190972 72208
rect 160100 72088 160152 72140
rect 161112 72088 161164 72140
rect 159732 72020 159784 72072
rect 194232 72088 194284 72140
rect 176292 72020 176344 72072
rect 176476 72020 176528 72072
rect 108672 71680 108724 71732
rect 114560 71680 114612 71732
rect 127624 71680 127676 71732
rect 138020 71680 138072 71732
rect 138296 71680 138348 71732
rect 157708 71680 157760 71732
rect 158352 71680 158404 71732
rect 159548 71680 159600 71732
rect 160008 71680 160060 71732
rect 169944 71680 169996 71732
rect 211528 71680 211580 71732
rect 212448 71680 212500 71732
rect 3516 71612 3568 71664
rect 8944 71612 8996 71664
rect 102600 71612 102652 71664
rect 151360 71612 151412 71664
rect 192852 71612 192904 71664
rect 99104 71544 99156 71596
rect 101496 71476 101548 71528
rect 135444 71476 135496 71528
rect 156788 71544 156840 71596
rect 157156 71544 157208 71596
rect 191196 71544 191248 71596
rect 192484 71544 192536 71596
rect 193128 71544 193180 71596
rect 202144 71544 202196 71596
rect 146944 71476 146996 71528
rect 156512 71476 156564 71528
rect 157064 71476 157116 71528
rect 191656 71476 191708 71528
rect 115296 71408 115348 71460
rect 148232 71408 148284 71460
rect 148692 71408 148744 71460
rect 160008 71408 160060 71460
rect 193864 71408 193916 71460
rect 122196 71340 122248 71392
rect 107660 71272 107712 71324
rect 108028 71272 108080 71324
rect 140504 71272 140556 71324
rect 170036 71340 170088 71392
rect 170864 71340 170916 71392
rect 171784 71340 171836 71392
rect 199568 71340 199620 71392
rect 153660 71272 153712 71324
rect 154304 71272 154356 71324
rect 169576 71272 169628 71324
rect 203524 71272 203576 71324
rect 111064 71204 111116 71256
rect 142344 71204 142396 71256
rect 161020 71204 161072 71256
rect 195612 71204 195664 71256
rect 118884 71136 118936 71188
rect 150256 71136 150308 71188
rect 160928 71136 160980 71188
rect 195520 71136 195572 71188
rect 71044 71068 71096 71120
rect 107384 71068 107436 71120
rect 137652 71068 137704 71120
rect 147036 71068 147088 71120
rect 184296 71068 184348 71120
rect 42800 71000 42852 71052
rect 101496 71000 101548 71052
rect 104900 71000 104952 71052
rect 132408 71000 132460 71052
rect 148968 71000 149020 71052
rect 200120 71000 200172 71052
rect 212448 71000 212500 71052
rect 480904 71000 480956 71052
rect 120356 70932 120408 70984
rect 149244 70932 149296 70984
rect 170864 70932 170916 70984
rect 204352 70932 204404 70984
rect 97448 70864 97500 70916
rect 151176 70864 151228 70916
rect 158536 70864 158588 70916
rect 191380 70864 191432 70916
rect 113548 70796 113600 70848
rect 128452 70796 128504 70848
rect 129556 70796 129608 70848
rect 165528 70796 165580 70848
rect 171784 70796 171836 70848
rect 178868 70796 178920 70848
rect 219808 70796 219860 70848
rect 149244 70728 149296 70780
rect 150072 70728 150124 70780
rect 97080 70320 97132 70372
rect 151912 70320 151964 70372
rect 168104 70320 168156 70372
rect 195060 70320 195112 70372
rect 97540 70184 97592 70236
rect 151084 70252 151136 70304
rect 165252 70252 165304 70304
rect 213000 70252 213052 70304
rect 115020 70184 115072 70236
rect 150716 70184 150768 70236
rect 162400 70184 162452 70236
rect 196440 70184 196492 70236
rect 98552 70116 98604 70168
rect 132776 70116 132828 70168
rect 162308 70116 162360 70168
rect 197084 70116 197136 70168
rect 108580 70048 108632 70100
rect 142436 70048 142488 70100
rect 164608 70048 164660 70100
rect 199752 70048 199804 70100
rect 108948 69980 109000 70032
rect 142528 69980 142580 70032
rect 164792 69980 164844 70032
rect 165252 69980 165304 70032
rect 199384 69980 199436 70032
rect 110972 69912 111024 69964
rect 144000 69912 144052 69964
rect 146944 69912 146996 69964
rect 161572 69912 161624 69964
rect 162308 69912 162360 69964
rect 164884 69912 164936 69964
rect 165436 69912 165488 69964
rect 166172 69912 166224 69964
rect 196992 69912 197044 69964
rect 101680 69844 101732 69896
rect 85580 69776 85632 69828
rect 105820 69776 105872 69828
rect 35992 69640 36044 69692
rect 101680 69640 101732 69692
rect 110236 69844 110288 69896
rect 142804 69844 142856 69896
rect 148416 69844 148468 69896
rect 196624 69844 196676 69896
rect 118792 69776 118844 69828
rect 152740 69776 152792 69828
rect 161664 69776 161716 69828
rect 162400 69776 162452 69828
rect 162584 69776 162636 69828
rect 189448 69776 189500 69828
rect 317420 69776 317472 69828
rect 134984 69708 135036 69760
rect 159180 69708 159232 69760
rect 193496 69708 193548 69760
rect 345020 69708 345072 69760
rect 138756 69640 138808 69692
rect 147496 69640 147548 69692
rect 182916 69640 182968 69692
rect 195060 69640 195112 69692
rect 368480 69640 368532 69692
rect 111708 69572 111760 69624
rect 142160 69572 142212 69624
rect 143080 69572 143132 69624
rect 161848 69572 161900 69624
rect 162584 69572 162636 69624
rect 163504 69572 163556 69624
rect 163964 69572 164016 69624
rect 102784 69504 102836 69556
rect 132500 69504 132552 69556
rect 166172 69504 166224 69556
rect 174268 69572 174320 69624
rect 175096 69572 175148 69624
rect 208676 69572 208728 69624
rect 198372 69504 198424 69556
rect 107200 69436 107252 69488
rect 120080 69436 120132 69488
rect 161756 69436 161808 69488
rect 162768 69436 162820 69488
rect 210424 69436 210476 69488
rect 120172 69368 120224 69420
rect 120724 69368 120776 69420
rect 141240 69300 141292 69352
rect 102784 69028 102836 69080
rect 105544 69028 105596 69080
rect 150716 69028 150768 69080
rect 151544 69028 151596 69080
rect 99288 68960 99340 69012
rect 153476 68960 153528 69012
rect 160376 68960 160428 69012
rect 214564 68960 214616 69012
rect 114100 68892 114152 68944
rect 115480 68824 115532 68876
rect 145104 68892 145156 68944
rect 147036 68892 147088 68944
rect 166080 68892 166132 68944
rect 166816 68892 166868 68944
rect 60740 68620 60792 68672
rect 102968 68756 103020 68808
rect 137100 68756 137152 68808
rect 148600 68824 148652 68876
rect 148876 68824 148928 68876
rect 165988 68824 166040 68876
rect 211896 68892 211948 68944
rect 171508 68824 171560 68876
rect 172152 68824 172204 68876
rect 172888 68824 172940 68876
rect 173716 68824 173768 68876
rect 177672 68824 177724 68876
rect 209964 68824 210016 68876
rect 211068 68824 211120 68876
rect 149520 68756 149572 68808
rect 165804 68756 165856 68808
rect 166448 68756 166500 68808
rect 171416 68756 171468 68808
rect 172336 68756 172388 68808
rect 175924 68756 175976 68808
rect 200672 68756 200724 68808
rect 108764 68688 108816 68740
rect 142712 68688 142764 68740
rect 142896 68688 142948 68740
rect 165712 68688 165764 68740
rect 166356 68688 166408 68740
rect 168840 68688 168892 68740
rect 169392 68688 169444 68740
rect 203432 68688 203484 68740
rect 103336 68620 103388 68672
rect 135628 68620 135680 68672
rect 166816 68620 166868 68672
rect 201224 68620 201276 68672
rect 34520 68552 34572 68604
rect 99840 68552 99892 68604
rect 112904 68552 112956 68604
rect 99196 68484 99248 68536
rect 131580 68484 131632 68536
rect 132684 68484 132736 68536
rect 140044 68552 140096 68604
rect 142252 68552 142304 68604
rect 149152 68552 149204 68604
rect 220820 68552 220872 68604
rect 144368 68484 144420 68536
rect 172336 68484 172388 68536
rect 205824 68484 205876 68536
rect 214564 68484 214616 68536
rect 358820 68484 358872 68536
rect 103152 68416 103204 68468
rect 134248 68416 134300 68468
rect 165344 68416 165396 68468
rect 197820 68416 197872 68468
rect 396080 68416 396132 68468
rect 40040 68348 40092 68400
rect 103336 68348 103388 68400
rect 110788 68348 110840 68400
rect 142712 68348 142764 68400
rect 142988 68348 143040 68400
rect 165896 68348 165948 68400
rect 193772 68348 193824 68400
rect 440240 68348 440292 68400
rect 97172 68280 97224 68332
rect 106280 68280 106332 68332
rect 139676 68280 139728 68332
rect 147312 68280 147364 68332
rect 189724 68280 189776 68332
rect 211068 68280 211120 68332
rect 536840 68280 536892 68332
rect 118976 68212 119028 68264
rect 141976 68212 142028 68264
rect 173716 68212 173768 68264
rect 207204 68212 207256 68264
rect 172152 68144 172204 68196
rect 205640 68144 205692 68196
rect 166448 68076 166500 68128
rect 175924 68076 175976 68128
rect 166356 68008 166408 68060
rect 200856 68076 200908 68128
rect 149520 67600 149572 67652
rect 149888 67600 149940 67652
rect 153476 67600 153528 67652
rect 154212 67600 154264 67652
rect 124864 67532 124916 67584
rect 135352 67532 135404 67584
rect 135904 67532 135956 67584
rect 96988 67464 97040 67516
rect 145656 67532 145708 67584
rect 146024 67532 146076 67584
rect 163412 67532 163464 67584
rect 164148 67532 164200 67584
rect 164516 67532 164568 67584
rect 165160 67532 165212 67584
rect 211620 67532 211672 67584
rect 166172 67464 166224 67516
rect 212724 67464 212776 67516
rect 119804 67396 119856 67448
rect 153292 67396 153344 67448
rect 157708 67396 157760 67448
rect 192576 67396 192628 67448
rect 193036 67396 193088 67448
rect 100024 67328 100076 67380
rect 133972 67328 134024 67380
rect 134524 67328 134576 67380
rect 165160 67328 165212 67380
rect 199660 67328 199712 67380
rect 100116 67260 100168 67312
rect 134064 67260 134116 67312
rect 134616 67260 134668 67312
rect 165620 67260 165672 67312
rect 166172 67260 166224 67312
rect 177028 67260 177080 67312
rect 177856 67260 177908 67312
rect 211344 67260 211396 67312
rect 100392 67192 100444 67244
rect 134156 67192 134208 67244
rect 166724 67192 166776 67244
rect 196164 67192 196216 67244
rect 104440 67124 104492 67176
rect 138848 67124 138900 67176
rect 175464 67124 175516 67176
rect 204904 67124 204956 67176
rect 77300 66920 77352 66972
rect 104440 66920 104492 66972
rect 44180 66852 44232 66904
rect 101772 66852 101824 66904
rect 136180 67056 136232 67108
rect 147956 67056 148008 67108
rect 203524 67056 203576 67108
rect 106924 66988 106976 67040
rect 109408 66988 109460 67040
rect 140136 66988 140188 67040
rect 154304 66988 154356 67040
rect 274640 66988 274692 67040
rect 107568 66920 107620 66972
rect 135536 66920 135588 66972
rect 159088 66920 159140 66972
rect 159732 66920 159784 66972
rect 188344 66920 188396 66972
rect 193036 66920 193088 66972
rect 332692 66920 332744 66972
rect 120080 66852 120132 66904
rect 120724 66852 120776 66904
rect 141148 66852 141200 66904
rect 165988 66852 166040 66904
rect 166816 66852 166868 66904
rect 120264 66784 120316 66836
rect 120816 66784 120868 66836
rect 141056 66784 141108 66836
rect 162124 66784 162176 66836
rect 188436 66852 188488 66904
rect 196164 66852 196216 66904
rect 196900 66852 196952 66904
rect 375380 66852 375432 66904
rect 97724 66716 97776 66768
rect 151268 66716 151320 66768
rect 153292 66240 153344 66292
rect 154028 66240 154080 66292
rect 110052 66172 110104 66224
rect 143908 66172 143960 66224
rect 147128 66172 147180 66224
rect 163320 66172 163372 66224
rect 164056 66172 164108 66224
rect 172796 66172 172848 66224
rect 173624 66172 173676 66224
rect 175372 66172 175424 66224
rect 176292 66172 176344 66224
rect 176936 66172 176988 66224
rect 177672 66172 177724 66224
rect 204904 66240 204956 66292
rect 554044 66240 554096 66292
rect 210240 66172 210292 66224
rect 104440 66104 104492 66156
rect 136916 66104 136968 66156
rect 211712 66104 211764 66156
rect 103244 66036 103296 66088
rect 103428 66036 103480 66088
rect 135812 66036 135864 66088
rect 164424 66036 164476 66088
rect 198924 66036 198976 66088
rect 93124 65900 93176 65952
rect 107016 65900 107068 65952
rect 139860 65968 139912 66020
rect 173624 65968 173676 66020
rect 205732 65968 205784 66020
rect 110328 65900 110380 65952
rect 142160 65900 142212 65952
rect 142620 65900 142672 65952
rect 154948 65900 155000 65952
rect 155684 65900 155736 65952
rect 186964 65900 187016 65952
rect 78680 65764 78732 65816
rect 104716 65764 104768 65816
rect 75920 65696 75972 65748
rect 104164 65696 104216 65748
rect 60832 65628 60884 65680
rect 105728 65628 105780 65680
rect 52552 65560 52604 65612
rect 103428 65560 103480 65612
rect 35164 65492 35216 65544
rect 103336 65492 103388 65544
rect 134432 65832 134484 65884
rect 164056 65832 164108 65884
rect 191288 65832 191340 65884
rect 113180 65764 113232 65816
rect 120264 65764 120316 65816
rect 160284 65764 160336 65816
rect 161020 65764 161072 65816
rect 187056 65764 187108 65816
rect 147864 65560 147916 65612
rect 209964 65560 210016 65612
rect 198924 65492 198976 65544
rect 418804 65492 418856 65544
rect 141516 64880 141568 64932
rect 142252 64880 142304 64932
rect 97816 64812 97868 64864
rect 144092 64812 144144 64864
rect 174176 64812 174228 64864
rect 214380 64812 214432 64864
rect 104164 64744 104216 64796
rect 138480 64744 138532 64796
rect 158996 64744 159048 64796
rect 193404 64744 193456 64796
rect 103796 64676 103848 64728
rect 137468 64676 137520 64728
rect 168656 64676 168708 64728
rect 203064 64676 203116 64728
rect 103980 64608 104032 64660
rect 132592 64608 132644 64660
rect 149796 64404 149848 64456
rect 224960 64404 225012 64456
rect 152648 64336 152700 64388
rect 256700 64336 256752 64388
rect 193404 64268 193456 64320
rect 340972 64268 341024 64320
rect 203064 64200 203116 64252
rect 472624 64200 472676 64252
rect 88340 64132 88392 64184
rect 104164 64132 104216 64184
rect 147404 64132 147456 64184
rect 183560 64132 183612 64184
rect 214380 64132 214432 64184
rect 543740 64132 543792 64184
rect 144368 63996 144420 64048
rect 147220 63996 147272 64048
rect 144092 63520 144144 63572
rect 144276 63520 144328 63572
rect 100576 63452 100628 63504
rect 134340 63452 134392 63504
rect 154764 63452 154816 63504
rect 215484 63452 215536 63504
rect 104348 63384 104400 63436
rect 104808 63384 104860 63436
rect 137192 63384 137244 63436
rect 168564 63384 168616 63436
rect 169300 63384 169352 63436
rect 203616 63384 203668 63436
rect 157616 63316 157668 63368
rect 192024 63316 192076 63368
rect 193036 63316 193088 63368
rect 168104 63248 168156 63300
rect 201500 63248 201552 63300
rect 167460 62908 167512 62960
rect 168104 62908 168156 62960
rect 72424 62840 72476 62892
rect 104348 62840 104400 62892
rect 197636 62840 197688 62892
rect 197820 62840 197872 62892
rect 215484 62840 215536 62892
rect 292580 62840 292632 62892
rect 27620 62772 27672 62824
rect 100576 62772 100628 62824
rect 108856 62772 108908 62824
rect 115940 62772 115992 62824
rect 116952 62772 117004 62824
rect 138664 62772 138716 62824
rect 142344 62772 142396 62824
rect 193036 62772 193088 62824
rect 331220 62772 331272 62824
rect 103520 62704 103572 62756
rect 108304 62704 108356 62756
rect 145932 62228 145984 62280
rect 148324 62228 148376 62280
rect 106832 62024 106884 62076
rect 117228 62024 117280 62076
rect 172704 62024 172756 62076
rect 212540 62024 212592 62076
rect 213828 62024 213880 62076
rect 163228 61956 163280 62008
rect 197636 61956 197688 62008
rect 151912 61548 151964 61600
rect 251180 61548 251232 61600
rect 154488 61480 154540 61532
rect 277400 61480 277452 61532
rect 197636 61412 197688 61464
rect 394700 61412 394752 61464
rect 146392 61344 146444 61396
rect 185584 61344 185636 61396
rect 213828 61344 213880 61396
rect 529940 61344 529992 61396
rect 98644 60664 98696 60716
rect 132960 60664 133012 60716
rect 145840 60664 145892 60716
rect 152648 60664 152700 60716
rect 154672 60664 154724 60716
rect 189080 60664 189132 60716
rect 189356 60664 189408 60716
rect 98000 60596 98052 60648
rect 105912 60596 105964 60648
rect 139768 60596 139820 60648
rect 158904 60596 158956 60648
rect 193312 60596 193364 60648
rect 194508 60596 194560 60648
rect 105820 60528 105872 60580
rect 106096 60528 106148 60580
rect 137008 60528 137060 60580
rect 167368 60528 167420 60580
rect 193680 60528 193732 60580
rect 194416 60528 194468 60580
rect 153108 60120 153160 60172
rect 259460 60120 259512 60172
rect 62120 60052 62172 60104
rect 105820 60052 105872 60104
rect 189080 60052 189132 60104
rect 299480 60052 299532 60104
rect 21364 59984 21416 60036
rect 98644 59984 98696 60036
rect 147312 59984 147364 60036
rect 187700 59984 187752 60036
rect 194508 59984 194560 60036
rect 349160 59984 349212 60036
rect 140136 59780 140188 59832
rect 142528 59780 142580 59832
rect 194416 59372 194468 59424
rect 459560 59372 459612 59424
rect 100760 59304 100812 59356
rect 101864 59304 101916 59356
rect 135720 59304 135772 59356
rect 167184 59304 167236 59356
rect 201776 59304 201828 59356
rect 202788 59304 202840 59356
rect 157524 59236 157576 59288
rect 192760 59236 192812 59288
rect 193036 59236 193088 59288
rect 193036 58692 193088 58744
rect 327080 58692 327132 58744
rect 48320 58624 48372 58676
rect 100760 58624 100812 58676
rect 202788 58624 202840 58676
rect 448520 58624 448572 58676
rect 168472 57876 168524 57928
rect 203248 57876 203300 57928
rect 204168 57876 204220 57928
rect 160192 57808 160244 57860
rect 194692 57808 194744 57860
rect 195060 57808 195112 57860
rect 156144 57740 156196 57792
rect 190460 57740 190512 57792
rect 191748 57740 191800 57792
rect 153016 57400 153068 57452
rect 263600 57400 263652 57452
rect 191748 57332 191800 57384
rect 309140 57332 309192 57384
rect 195060 57264 195112 57316
rect 362960 57264 363012 57316
rect 204168 57196 204220 57248
rect 473452 57196 473504 57248
rect 178776 56516 178828 56568
rect 217048 56516 217100 56568
rect 167000 56448 167052 56500
rect 201868 56448 201920 56500
rect 202788 56448 202840 56500
rect 163136 56380 163188 56432
rect 197636 56380 197688 56432
rect 158812 56312 158864 56364
rect 193220 56312 193272 56364
rect 194508 56312 194560 56364
rect 156052 56244 156104 56296
rect 189080 56244 189132 56296
rect 150256 56176 150308 56228
rect 220084 56176 220136 56228
rect 189080 56108 189132 56160
rect 313280 56108 313332 56160
rect 194508 56040 194560 56092
rect 351920 56040 351972 56092
rect 197636 55972 197688 56024
rect 398840 55972 398892 56024
rect 202788 55904 202840 55956
rect 448612 55904 448664 55956
rect 217048 55836 217100 55888
rect 564532 55836 564584 55888
rect 109592 55156 109644 55208
rect 138388 55156 138440 55208
rect 164332 55156 164384 55208
rect 198832 55156 198884 55208
rect 168380 55088 168432 55140
rect 202880 55088 202932 55140
rect 198832 54544 198884 54596
rect 414664 54544 414716 54596
rect 202880 54476 202932 54528
rect 464344 54476 464396 54528
rect 172060 53728 172112 53780
rect 204260 53728 204312 53780
rect 166264 53660 166316 53712
rect 198096 53660 198148 53712
rect 151636 53184 151688 53236
rect 242900 53184 242952 53236
rect 198096 53116 198148 53168
rect 402980 53116 403032 53168
rect 204260 53048 204312 53100
rect 490012 53048 490064 53100
rect 197452 52504 197504 52556
rect 197636 52504 197688 52556
rect 155960 52368 156012 52420
rect 189632 52368 189684 52420
rect 150164 51688 150216 51740
rect 217324 51688 217376 51740
rect 189632 51076 189684 51128
rect 320180 51076 320232 51128
rect 157432 51008 157484 51060
rect 192668 51008 192720 51060
rect 193036 51008 193088 51060
rect 176844 50940 176896 50992
rect 208492 50940 208544 50992
rect 193036 50396 193088 50448
rect 338120 50396 338172 50448
rect 110420 50328 110472 50380
rect 119344 50328 119396 50380
rect 145748 50328 145800 50380
rect 167644 50328 167696 50380
rect 208492 50328 208544 50380
rect 209136 50328 209188 50380
rect 569960 50328 570012 50380
rect 143816 49648 143868 49700
rect 148416 49648 148468 49700
rect 154580 49648 154632 49700
rect 189448 49648 189500 49700
rect 147680 49104 147732 49156
rect 201592 49104 201644 49156
rect 189448 48968 189500 49020
rect 190184 48968 190236 49020
rect 285680 48968 285732 49020
rect 148692 47608 148744 47660
rect 204260 47608 204312 47660
rect 150072 47540 150124 47592
rect 215300 47540 215352 47592
rect 135260 46928 135312 46980
rect 142436 46928 142488 46980
rect 176752 46860 176804 46912
rect 208492 46860 208544 46912
rect 209044 46860 209096 46912
rect 151544 46248 151596 46300
rect 233240 46248 233292 46300
rect 208492 46180 208544 46232
rect 571984 46180 572036 46232
rect 172612 45500 172664 45552
rect 205916 45500 205968 45552
rect 148600 44820 148652 44872
rect 198740 44820 198792 44872
rect 205916 44140 205968 44192
rect 520924 44140 520976 44192
rect 176660 44072 176712 44124
rect 210148 44072 210200 44124
rect 211068 44072 211120 44124
rect 152924 43528 152976 43580
rect 267740 43528 267792 43580
rect 163044 43460 163096 43512
rect 408500 43460 408552 43512
rect 167276 43392 167328 43444
rect 458180 43392 458232 43444
rect 211068 42780 211120 42832
rect 576860 42780 576912 42832
rect 151452 42304 151504 42356
rect 239404 42304 239456 42356
rect 159732 42236 159784 42288
rect 350540 42236 350592 42288
rect 164240 42168 164292 42220
rect 426440 42168 426492 42220
rect 166356 42100 166408 42152
rect 438860 42100 438912 42152
rect 70400 42032 70452 42084
rect 136640 42032 136692 42084
rect 145564 42032 145616 42084
rect 167000 42032 167052 42084
rect 169760 42032 169812 42084
rect 495440 42032 495492 42084
rect 156604 40876 156656 40928
rect 307024 40876 307076 40928
rect 167092 40808 167144 40860
rect 462320 40808 462372 40860
rect 172244 40740 172296 40792
rect 498292 40740 498344 40792
rect 174912 40672 174964 40724
rect 535460 40672 535512 40724
rect 177488 39992 177540 40044
rect 213920 39992 213972 40044
rect 214380 39992 214432 40044
rect 151360 39584 151412 39636
rect 236000 39584 236052 39636
rect 165068 39516 165120 39568
rect 409880 39516 409932 39568
rect 214380 39448 214432 39500
rect 518900 39448 518952 39500
rect 173532 39380 173584 39432
rect 516140 39380 516192 39432
rect 77392 39312 77444 39364
rect 138296 39312 138348 39364
rect 176108 39312 176160 39364
rect 558920 39312 558972 39364
rect 138020 38972 138072 39024
rect 142896 38972 142948 39024
rect 152832 38088 152884 38140
rect 257344 38088 257396 38140
rect 169392 38020 169444 38072
rect 463700 38020 463752 38072
rect 169484 37952 169536 38004
rect 476120 37952 476172 38004
rect 13820 37884 13872 37936
rect 132776 37884 132828 37936
rect 145656 37884 145708 37936
rect 168472 37884 168524 37936
rect 172520 37884 172572 37936
rect 525064 37884 525116 37936
rect 148508 36864 148560 36916
rect 205640 36864 205692 36916
rect 154396 36796 154448 36848
rect 267832 36796 267884 36848
rect 162216 36728 162268 36780
rect 361580 36728 361632 36780
rect 170496 36660 170548 36712
rect 481640 36660 481692 36712
rect 172152 36592 172204 36644
rect 503720 36592 503772 36644
rect 175004 36524 175056 36576
rect 534080 36524 534132 36576
rect 169300 35232 169352 35284
rect 467840 35232 467892 35284
rect 31760 35164 31812 35216
rect 133972 35164 134024 35216
rect 175280 35164 175332 35216
rect 552020 35164 552072 35216
rect 159916 34008 159968 34060
rect 346400 34008 346452 34060
rect 168104 33940 168156 33992
rect 446404 33940 446456 33992
rect 170680 33872 170732 33924
rect 488540 33872 488592 33924
rect 144276 33804 144328 33856
rect 145012 33804 145064 33856
rect 176200 33804 176252 33856
rect 565820 33804 565872 33856
rect 45560 33736 45612 33788
rect 135352 33736 135404 33788
rect 145472 33736 145524 33788
rect 171784 33736 171836 33788
rect 177672 33736 177724 33788
rect 578240 33736 578292 33788
rect 3516 33056 3568 33108
rect 95884 33056 95936 33108
rect 149980 32512 150032 32564
rect 225604 32512 225656 32564
rect 151728 32444 151780 32496
rect 242992 32444 243044 32496
rect 159824 32376 159876 32428
rect 339500 32376 339552 32428
rect 152740 31152 152792 31204
rect 264980 31152 265032 31204
rect 160928 31084 160980 31136
rect 357440 31084 357492 31136
rect 17316 31016 17368 31068
rect 132868 31016 132920 31068
rect 169576 31016 169628 31068
rect 470600 31016 470652 31068
rect 155592 29792 155644 29844
rect 299572 29792 299624 29844
rect 162952 29724 163004 29776
rect 407212 29724 407264 29776
rect 170772 29656 170824 29708
rect 491300 29656 491352 29708
rect 24860 29588 24912 29640
rect 134156 29588 134208 29640
rect 177764 29588 177816 29640
rect 574100 29588 574152 29640
rect 158352 28432 158404 28484
rect 321560 28432 321612 28484
rect 166448 28364 166500 28416
rect 427820 28364 427872 28416
rect 171324 28296 171376 28348
rect 502340 28296 502392 28348
rect 184848 28228 184900 28280
rect 582380 28228 582432 28280
rect 154212 27140 154264 27192
rect 275284 27140 275336 27192
rect 162308 27072 162360 27124
rect 374092 27072 374144 27124
rect 165160 27004 165212 27056
rect 410524 27004 410576 27056
rect 171232 26936 171284 26988
rect 506572 26936 506624 26988
rect 144920 26868 144972 26920
rect 171876 26868 171928 26920
rect 172336 26868 172388 26920
rect 510620 26868 510672 26920
rect 154120 25780 154172 25832
rect 278780 25780 278832 25832
rect 162400 25712 162452 25764
rect 378140 25712 378192 25764
rect 165252 25644 165304 25696
rect 418160 25644 418212 25696
rect 171140 25576 171192 25628
rect 509240 25576 509292 25628
rect 173716 25508 173768 25560
rect 524420 25508 524472 25560
rect 154304 24284 154356 24336
rect 282920 24284 282972 24336
rect 163964 24216 164016 24268
rect 391940 24216 391992 24268
rect 172428 24148 172480 24200
rect 513380 24148 513432 24200
rect 173624 24080 173676 24132
rect 531412 24080 531464 24132
rect 157064 22992 157116 23044
rect 310520 22992 310572 23044
rect 162860 22924 162912 22976
rect 398932 22924 398984 22976
rect 166632 22856 166684 22908
rect 440332 22856 440384 22908
rect 173808 22788 173860 22840
rect 520280 22788 520332 22840
rect 175096 22720 175148 22772
rect 538956 22720 539008 22772
rect 143724 21360 143776 21412
rect 157984 21360 158036 21412
rect 158444 21360 158496 21412
rect 329104 21360 329156 21412
rect 342904 21360 342956 21412
rect 471980 21360 472032 21412
rect 153844 20136 153896 20188
rect 280160 20136 280212 20188
rect 155224 20068 155276 20120
rect 291200 20068 291252 20120
rect 155684 20000 155736 20052
rect 287060 20000 287112 20052
rect 287704 20000 287756 20052
rect 456892 20000 456944 20052
rect 161020 19932 161072 19984
rect 357532 19932 357584 19984
rect 154028 18776 154080 18828
rect 273260 18776 273312 18828
rect 166172 18708 166224 18760
rect 431960 18708 432012 18760
rect 176292 18640 176344 18692
rect 567200 18640 567252 18692
rect 177948 18572 178000 18624
rect 571340 18572 571392 18624
rect 149888 17416 149940 17468
rect 219440 17416 219492 17468
rect 168196 17348 168248 17400
rect 445760 17348 445812 17400
rect 169668 17280 169720 17332
rect 477500 17280 477552 17332
rect 177856 17212 177908 17264
rect 570604 17212 570656 17264
rect 149704 16124 149756 16176
rect 227536 16124 227588 16176
rect 161112 16056 161164 16108
rect 361120 16056 361172 16108
rect 161204 15988 161256 16040
rect 364616 15988 364668 16040
rect 165344 15920 165396 15972
rect 420920 15920 420972 15972
rect 176384 15852 176436 15904
rect 560392 15852 560444 15904
rect 155776 14696 155828 14748
rect 293224 14696 293276 14748
rect 157156 14628 157208 14680
rect 314660 14628 314712 14680
rect 162676 14560 162728 14612
rect 385960 14560 386012 14612
rect 164056 14492 164108 14544
rect 404360 14492 404412 14544
rect 30104 14424 30156 14476
rect 133880 14424 133932 14476
rect 170956 14424 171008 14476
rect 493048 14424 493100 14476
rect 153936 13336 153988 13388
rect 272432 13336 272484 13388
rect 157248 13268 157300 13320
rect 307944 13268 307996 13320
rect 162584 13200 162636 13252
rect 382372 13200 382424 13252
rect 162492 13132 162544 13184
rect 386696 13132 386748 13184
rect 144184 13064 144236 13116
rect 155408 13064 155460 13116
rect 170864 13064 170916 13116
rect 486332 13064 486384 13116
rect 486424 13064 486476 13116
rect 581736 13064 581788 13116
rect 151176 11976 151228 12028
rect 241704 11976 241756 12028
rect 157340 11908 157392 11960
rect 328736 11908 328788 11960
rect 162768 11840 162820 11892
rect 379520 11840 379572 11892
rect 165436 11772 165488 11824
rect 417424 11772 417476 11824
rect 174084 11704 174136 11756
rect 541992 11704 542044 11756
rect 209964 11636 210016 11688
rect 210976 11636 211028 11688
rect 234620 11636 234672 11688
rect 235816 11636 235868 11688
rect 259460 11636 259512 11688
rect 260656 11636 260708 11688
rect 151268 10548 151320 10600
rect 234620 10548 234672 10600
rect 158536 10480 158588 10532
rect 336280 10480 336332 10532
rect 160100 10412 160152 10464
rect 372896 10412 372948 10464
rect 166724 10344 166776 10396
rect 432052 10344 432104 10396
rect 87512 10276 87564 10328
rect 138112 10276 138164 10328
rect 173992 10276 174044 10328
rect 548616 10276 548668 10328
rect 155868 9120 155920 9172
rect 301964 9120 302016 9172
rect 158628 9052 158680 9104
rect 325608 9052 325660 9104
rect 165528 8984 165580 9036
rect 414296 8984 414348 9036
rect 143632 8916 143684 8968
rect 157800 8916 157852 8968
rect 176476 8916 176528 8968
rect 556160 8916 556212 8968
rect 160008 7828 160060 7880
rect 343364 7828 343416 7880
rect 161388 7760 161440 7812
rect 365812 7760 365864 7812
rect 166908 7692 166960 7744
rect 435548 7692 435600 7744
rect 166816 7624 166868 7676
rect 442632 7624 442684 7676
rect 54944 7556 54996 7608
rect 135536 7556 135588 7608
rect 173900 7556 173952 7608
rect 538404 7556 538456 7608
rect 3424 6808 3476 6860
rect 17224 6808 17276 6860
rect 152556 6536 152608 6588
rect 252376 6536 252428 6588
rect 158720 6468 158772 6520
rect 350448 6468 350500 6520
rect 180064 6400 180116 6452
rect 436744 6400 436796 6452
rect 182088 6332 182140 6384
rect 443828 6332 443880 6384
rect 179144 6264 179196 6316
rect 450912 6264 450964 6316
rect 168288 6196 168340 6248
rect 453212 6196 453264 6248
rect 453304 6196 453356 6248
rect 479340 6196 479392 6248
rect 28908 6128 28960 6180
rect 134064 6128 134116 6180
rect 176568 6128 176620 6180
rect 563244 6128 563296 6180
rect 143540 5652 143592 5704
rect 144736 5652 144788 5704
rect 142804 5516 142856 5568
rect 143540 5516 143592 5568
rect 151084 5040 151136 5092
rect 245200 5040 245252 5092
rect 161204 4972 161256 5024
rect 371700 4972 371752 5024
rect 164148 4904 164200 4956
rect 397736 4904 397788 4956
rect 171048 4836 171100 4888
rect 482836 4836 482888 4888
rect 175188 4768 175240 4820
rect 545488 4768 545540 4820
rect 572 4088 624 4140
rect 7564 4088 7616 4140
rect 15936 4088 15988 4140
rect 17316 4088 17368 4140
rect 73804 4088 73856 4140
rect 75184 4088 75236 4140
rect 181996 4088 182048 4140
rect 187424 4088 187476 4140
rect 188344 4088 188396 4140
rect 193864 4088 193916 4140
rect 194048 4088 194100 4140
rect 195612 4088 195664 4140
rect 196624 4088 196676 4140
rect 203892 4088 203944 4140
rect 203984 4088 204036 4140
rect 247592 4088 247644 4140
rect 247684 4088 247736 4140
rect 254676 4088 254728 4140
rect 257344 4088 257396 4140
rect 258264 4088 258316 4140
rect 261484 4088 261536 4140
rect 262956 4088 263008 4140
rect 283564 4088 283616 4140
rect 298468 4088 298520 4140
rect 450544 4088 450596 4140
rect 452108 4088 452160 4140
rect 563704 4088 563756 4140
rect 569132 4088 569184 4140
rect 6460 4020 6512 4072
rect 7656 4020 7708 4072
rect 102232 4020 102284 4072
rect 113272 4020 113324 4072
rect 119896 4020 119948 4072
rect 122104 4020 122156 4072
rect 146852 4020 146904 4072
rect 153016 4020 153068 4072
rect 182824 4020 182876 4072
rect 212172 4020 212224 4072
rect 224224 4020 224276 4072
rect 284300 4020 284352 4072
rect 299572 4020 299624 4072
rect 300768 4020 300820 4072
rect 311164 4020 311216 4072
rect 312636 4020 312688 4072
rect 85672 3952 85724 4004
rect 88984 3952 89036 4004
rect 111616 3952 111668 4004
rect 129832 3952 129884 4004
rect 179328 3952 179380 4004
rect 394240 3952 394292 4004
rect 83280 3884 83332 3936
rect 127164 3884 127216 3936
rect 179236 3884 179288 3936
rect 401324 3884 401376 3936
rect 65524 3816 65576 3868
rect 69112 3748 69164 3800
rect 71044 3748 71096 3800
rect 72608 3816 72660 3868
rect 130016 3816 130068 3868
rect 130936 3816 130988 3868
rect 150624 3816 150676 3868
rect 152648 3816 152700 3868
rect 164884 3816 164936 3868
rect 178960 3816 179012 3868
rect 408408 3816 408460 3868
rect 410524 3816 410576 3868
rect 411904 3816 411956 3868
rect 131304 3748 131356 3800
rect 146944 3748 146996 3800
rect 39580 3680 39632 3732
rect 131396 3680 131448 3732
rect 137652 3680 137704 3732
rect 138664 3680 138716 3732
rect 147036 3680 147088 3732
rect 149520 3680 149572 3732
rect 149796 3748 149848 3800
rect 156604 3748 156656 3800
rect 156788 3748 156840 3800
rect 170772 3748 170824 3800
rect 184112 3748 184164 3800
rect 415492 3748 415544 3800
rect 163688 3680 163740 3732
rect 180616 3680 180668 3732
rect 422576 3680 422628 3732
rect 489184 3680 489236 3732
rect 491116 3680 491168 3732
rect 7656 3612 7708 3664
rect 11152 3544 11204 3596
rect 13084 3544 13136 3596
rect 21824 3612 21876 3664
rect 124220 3612 124272 3664
rect 124680 3612 124732 3664
rect 129924 3612 129976 3664
rect 131028 3612 131080 3664
rect 162492 3612 162544 3664
rect 180708 3612 180760 3664
rect 429660 3612 429712 3664
rect 431960 3612 432012 3664
rect 433248 3612 433300 3664
rect 454684 3612 454736 3664
rect 497096 3612 497148 3664
rect 127072 3544 127124 3596
rect 128268 3544 128320 3596
rect 166080 3544 166132 3596
rect 176660 3544 176712 3596
rect 179512 3544 179564 3596
rect 185584 3544 185636 3596
rect 187332 3544 187384 3596
rect 187424 3544 187476 3596
rect 461584 3544 461636 3596
rect 525064 3544 525116 3596
rect 527824 3544 527876 3596
rect 574744 3544 574796 3596
rect 576308 3544 576360 3596
rect 4068 3476 4120 3528
rect 4804 3476 4856 3528
rect 5264 3476 5316 3528
rect 17040 3408 17092 3460
rect 18604 3408 18656 3460
rect 20628 3408 20680 3460
rect 33600 3340 33652 3392
rect 35164 3340 35216 3392
rect 38384 3340 38436 3392
rect 39304 3340 39356 3392
rect 52460 3340 52512 3392
rect 53380 3340 53432 3392
rect 56048 3340 56100 3392
rect 57244 3340 57296 3392
rect 91560 3340 91612 3392
rect 93124 3340 93176 3392
rect 102140 3340 102192 3392
rect 103336 3340 103388 3392
rect 105728 3340 105780 3392
rect 106924 3340 106976 3392
rect 109316 3340 109368 3392
rect 111248 3340 111300 3392
rect 51356 3272 51408 3324
rect 54484 3272 54536 3324
rect 101036 3272 101088 3324
rect 102784 3272 102836 3324
rect 93952 3136 94004 3188
rect 95976 3136 96028 3188
rect 126980 3476 127032 3528
rect 128176 3476 128228 3528
rect 140044 3476 140096 3528
rect 141516 3476 141568 3528
rect 157984 3476 158036 3528
rect 158904 3476 158956 3528
rect 134156 3408 134208 3460
rect 140136 3408 140188 3460
rect 147220 3408 147272 3460
rect 148324 3408 148376 3460
rect 131580 3340 131632 3392
rect 152464 3340 152516 3392
rect 171968 3476 172020 3528
rect 173256 3476 173308 3528
rect 177856 3476 177908 3528
rect 178684 3476 178736 3528
rect 190828 3476 190880 3528
rect 193864 3476 193916 3528
rect 196808 3476 196860 3528
rect 198004 3476 198056 3528
rect 203984 3476 204036 3528
rect 167644 3408 167696 3460
rect 168380 3408 168432 3460
rect 171784 3408 171836 3460
rect 173164 3408 173216 3460
rect 179052 3408 179104 3460
rect 198096 3408 198148 3460
rect 126980 3272 127032 3324
rect 128452 3272 128504 3324
rect 148416 3272 148468 3324
rect 175464 3340 175516 3392
rect 184296 3340 184348 3392
rect 189724 3340 189776 3392
rect 189816 3340 189868 3392
rect 193220 3340 193272 3392
rect 193128 3272 193180 3324
rect 198096 3272 198148 3324
rect 465172 3408 465224 3460
rect 468484 3408 468536 3460
rect 469864 3408 469916 3460
rect 472624 3476 472676 3528
rect 473452 3476 473504 3528
rect 475384 3476 475436 3528
rect 475752 3408 475804 3460
rect 486516 3476 486568 3528
rect 487620 3476 487672 3528
rect 493324 3476 493376 3528
rect 507676 3408 507728 3460
rect 207664 3340 207716 3392
rect 223948 3340 224000 3392
rect 225604 3340 225656 3392
rect 226340 3340 226392 3392
rect 239404 3340 239456 3392
rect 240508 3340 240560 3392
rect 275284 3340 275336 3392
rect 276020 3340 276072 3392
rect 307024 3340 307076 3392
rect 309048 3340 309100 3392
rect 329104 3340 329156 3392
rect 330392 3340 330444 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 340972 3340 341024 3392
rect 342168 3340 342220 3392
rect 357532 3340 357584 3392
rect 358728 3340 358780 3392
rect 364984 3340 365036 3392
rect 367008 3340 367060 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 390560 3340 390612 3392
rect 391848 3340 391900 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 400864 3340 400916 3392
rect 402520 3340 402572 3392
rect 414664 3340 414716 3392
rect 416688 3340 416740 3392
rect 418804 3340 418856 3392
rect 420184 3340 420236 3392
rect 422944 3340 422996 3392
rect 424968 3340 425020 3392
rect 432604 3340 432656 3392
rect 434444 3340 434496 3392
rect 440240 3340 440292 3392
rect 441528 3340 441580 3392
rect 446404 3340 446456 3392
rect 447416 3340 447468 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 456892 3340 456944 3392
rect 458088 3340 458140 3392
rect 514024 3476 514076 3528
rect 515956 3476 516008 3528
rect 545764 3476 545816 3528
rect 551468 3476 551520 3528
rect 554044 3476 554096 3528
rect 554964 3476 555016 3528
rect 560944 3476 560996 3528
rect 564440 3476 564492 3528
rect 571984 3476 572036 3528
rect 573916 3476 573968 3528
rect 511356 3408 511408 3460
rect 514760 3408 514812 3460
rect 527916 3408 527968 3460
rect 533712 3408 533764 3460
rect 538956 3408 539008 3460
rect 539600 3408 539652 3460
rect 570604 3408 570656 3460
rect 572720 3408 572772 3460
rect 518348 3340 518400 3392
rect 520924 3272 520976 3324
rect 524236 3272 524288 3324
rect 125876 3204 125928 3256
rect 131488 3204 131540 3256
rect 342996 3204 343048 3256
rect 344560 3204 344612 3256
rect 552756 3204 552808 3256
rect 553768 3204 553820 3256
rect 131120 3136 131172 3188
rect 136456 3136 136508 3188
rect 139952 3136 140004 3188
rect 148508 3136 148560 3188
rect 154212 3136 154264 3188
rect 220084 3136 220136 3188
rect 222752 3136 222804 3188
rect 315304 3136 315356 3188
rect 317328 3136 317380 3188
rect 538864 3136 538916 3188
rect 546684 3136 546736 3188
rect 217324 3068 217376 3120
rect 218060 3068 218112 3120
rect 1676 3000 1728 3052
rect 9036 3000 9088 3052
rect 19432 3000 19484 3052
rect 21364 3000 21416 3052
rect 23020 3000 23072 3052
rect 25504 3000 25556 3052
rect 118792 3000 118844 3052
rect 120724 3000 120776 3052
rect 123484 3000 123536 3052
rect 125600 3000 125652 3052
rect 141240 3000 141292 3052
rect 142712 3000 142764 3052
rect 182916 3000 182968 3052
rect 186136 3000 186188 3052
rect 324964 3000 325016 3052
rect 326804 3000 326856 3052
rect 382924 3000 382976 3052
rect 384764 3000 384816 3052
rect 464344 3000 464396 3052
rect 466276 3000 466328 3052
rect 503076 3000 503128 3052
rect 505376 3000 505428 3052
rect 12348 2932 12400 2984
rect 14464 2932 14516 2984
rect 132960 2932 133012 2984
rect 141424 2932 141476 2984
rect 171876 2932 171928 2984
rect 174268 2932 174320 2984
rect 70308 2864 70360 2916
rect 72424 2864 72476 2916
rect 203524 2864 203576 2916
rect 207388 2864 207440 2916
rect 480904 2864 480956 2916
rect 484032 2864 484084 2916
rect 382280 960 382332 1012
rect 383568 960 383620 1012
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700398 8156 703520
rect 24320 700466 24348 703520
rect 24308 700460 24360 700466
rect 24308 700402 24360 700408
rect 8116 700392 8168 700398
rect 8116 700334 8168 700340
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 2778 514856 2834 514865
rect 2778 514791 2780 514800
rect 2832 514791 2834 514800
rect 4804 514820 4856 514826
rect 2780 514762 2832 514768
rect 4804 514762 4856 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 409902 2912 410479
rect 2872 409896 2924 409902
rect 2872 409838 2924 409844
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3436 268394 3464 475623
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3516 397520 3568 397526
rect 3514 397488 3516 397497
rect 3568 397488 3570 397497
rect 3514 397423 3570 397432
rect 3514 371376 3570 371385
rect 3514 371311 3570 371320
rect 3528 371278 3556 371311
rect 3516 371272 3568 371278
rect 3516 371214 3568 371220
rect 3514 345400 3570 345409
rect 3514 345335 3570 345344
rect 3528 345234 3556 345335
rect 3516 345228 3568 345234
rect 3516 345170 3568 345176
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3528 305046 3556 306167
rect 3516 305040 3568 305046
rect 3516 304982 3568 304988
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3528 292602 3556 293111
rect 3516 292596 3568 292602
rect 3516 292538 3568 292544
rect 4816 289134 4844 514762
rect 7564 345228 7616 345234
rect 7564 345170 7616 345176
rect 4804 289128 4856 289134
rect 4804 289070 4856 289076
rect 7576 269890 7604 345170
rect 40052 275330 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 40040 275324 40092 275330
rect 40040 275266 40092 275272
rect 71792 273970 71820 702986
rect 89180 700534 89208 703520
rect 89168 700528 89220 700534
rect 89168 700470 89220 700476
rect 105464 699718 105492 703520
rect 137848 700738 137876 703520
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 137836 700732 137888 700738
rect 137836 700674 137888 700680
rect 148324 700324 148376 700330
rect 148324 700266 148376 700272
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106924 699712 106976 699718
rect 106924 699654 106976 699660
rect 71780 273964 71832 273970
rect 71780 273906 71832 273912
rect 7564 269884 7616 269890
rect 7564 269826 7616 269832
rect 3424 268388 3476 268394
rect 3424 268330 3476 268336
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 106936 265674 106964 699654
rect 146300 696992 146352 696998
rect 146300 696934 146352 696940
rect 143540 616888 143592 616894
rect 143540 616830 143592 616836
rect 142160 590708 142212 590714
rect 142160 590650 142212 590656
rect 139400 484424 139452 484430
rect 139400 484366 139452 484372
rect 138664 430636 138716 430642
rect 138664 430578 138716 430584
rect 113824 357468 113876 357474
rect 113824 357410 113876 357416
rect 113836 291854 113864 357410
rect 135260 351960 135312 351966
rect 135260 351902 135312 351908
rect 134524 324352 134576 324358
rect 134524 324294 134576 324300
rect 113824 291848 113876 291854
rect 113824 291790 113876 291796
rect 132500 271924 132552 271930
rect 132500 271866 132552 271872
rect 120816 268388 120868 268394
rect 120816 268330 120868 268336
rect 120828 267782 120856 268330
rect 120816 267776 120868 267782
rect 120868 267724 120948 267734
rect 120816 267718 120948 267724
rect 120828 267706 120948 267718
rect 106924 265668 106976 265674
rect 106924 265610 106976 265616
rect 118332 265260 118384 265266
rect 118332 265202 118384 265208
rect 114192 265192 114244 265198
rect 114192 265134 114244 265140
rect 111524 263628 111576 263634
rect 111524 263570 111576 263576
rect 3424 263152 3476 263158
rect 3424 263094 3476 263100
rect 3332 241120 3384 241126
rect 3330 241088 3332 241097
rect 3384 241088 3386 241097
rect 3330 241023 3386 241032
rect 2780 215280 2832 215286
rect 2780 215222 2832 215228
rect 2792 214985 2820 215222
rect 2778 214976 2834 214985
rect 2778 214911 2834 214920
rect 3436 188873 3464 263094
rect 111430 262848 111486 262857
rect 111430 262783 111486 262792
rect 109776 262676 109828 262682
rect 109776 262618 109828 262624
rect 3608 262608 3660 262614
rect 3608 262550 3660 262556
rect 3516 262540 3568 262546
rect 3516 262482 3568 262488
rect 3528 201929 3556 262482
rect 3620 254153 3648 262550
rect 4804 261452 4856 261458
rect 4804 261394 4856 261400
rect 3606 254144 3662 254153
rect 3606 254079 3662 254088
rect 4816 215286 4844 261394
rect 7564 260228 7616 260234
rect 7564 260170 7616 260176
rect 7576 241126 7604 260170
rect 7564 241120 7616 241126
rect 7564 241062 7616 241068
rect 4804 215280 4856 215286
rect 4804 215222 4856 215228
rect 3514 201920 3570 201929
rect 3514 201855 3570 201864
rect 108948 200592 109000 200598
rect 108948 200534 109000 200540
rect 107568 200456 107620 200462
rect 107568 200398 107620 200404
rect 104532 199640 104584 199646
rect 104532 199582 104584 199588
rect 97632 199572 97684 199578
rect 97632 199514 97684 199520
rect 96436 193860 96488 193866
rect 96436 193802 96488 193808
rect 96344 189780 96396 189786
rect 96344 189722 96396 189728
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3514 162888 3570 162897
rect 3514 162823 3570 162832
rect 3146 149832 3202 149841
rect 3146 149767 3202 149776
rect 3160 149190 3188 149767
rect 3148 149184 3200 149190
rect 3148 149126 3200 149132
rect 3528 145586 3556 162823
rect 96252 154148 96304 154154
rect 96252 154090 96304 154096
rect 96160 154012 96212 154018
rect 96160 153954 96212 153960
rect 95884 153264 95936 153270
rect 95884 153206 95936 153212
rect 3516 145580 3568 145586
rect 3516 145522 3568 145528
rect 8944 140820 8996 140826
rect 8944 140762 8996 140768
rect 4804 139528 4856 139534
rect 4804 139470 4856 139476
rect 3424 138712 3476 138718
rect 3424 138654 3476 138660
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 2780 110832 2832 110838
rect 2780 110774 2832 110780
rect 2792 110673 2820 110774
rect 2778 110664 2834 110673
rect 2778 110599 2834 110608
rect 2778 77888 2834 77897
rect 2778 77823 2834 77832
rect 2792 16574 2820 77823
rect 3436 19417 3464 138654
rect 4816 110838 4844 139470
rect 4804 110832 4856 110838
rect 4804 110774 4856 110780
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 7562 75168 7618 75177
rect 7562 75103 7618 75112
rect 3516 71664 3568 71670
rect 3514 71632 3516 71641
rect 3568 71632 3570 71641
rect 3514 71567 3570 71576
rect 4802 64152 4858 64161
rect 4802 64087 4858 64096
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 2792 16546 2912 16574
rect 572 4140 624 4146
rect 572 4082 624 4088
rect 584 480 612 4082
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1688 480 1716 2994
rect 2884 480 2912 16546
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4816 3534 4844 64087
rect 7576 4146 7604 75103
rect 8298 72448 8354 72457
rect 8298 72383 8354 72392
rect 7654 66872 7710 66881
rect 7654 66807 7710 66816
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7668 4078 7696 66807
rect 8312 16574 8340 72383
rect 8956 71670 8984 140762
rect 17222 139496 17278 139505
rect 17222 139431 17278 139440
rect 13082 76528 13138 76537
rect 13082 76463 13138 76472
rect 8944 71664 8996 71670
rect 8944 71606 8996 71612
rect 9678 71224 9734 71233
rect 9678 71159 9734 71168
rect 9034 71088 9090 71097
rect 9034 71023 9090 71032
rect 8312 16546 8800 16574
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 4080 480 4108 3470
rect 5276 480 5304 3470
rect 6472 480 6500 4014
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7668 480 7696 3606
rect 8772 480 8800 16546
rect 9048 3058 9076 71023
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 71159
rect 12438 55856 12494 55865
rect 12438 55791 12494 55800
rect 12452 16574 12480 55791
rect 12452 16546 13032 16574
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11164 480 11192 3538
rect 13004 3482 13032 16546
rect 13096 3602 13124 76463
rect 14462 73808 14518 73817
rect 14462 73743 14518 73752
rect 13820 37936 13872 37942
rect 13820 37878 13872 37884
rect 13832 16574 13860 37878
rect 13832 16546 14320 16574
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 13004 3454 13584 3482
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12360 480 12388 2926
rect 13556 480 13584 3454
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 14476 2990 14504 73743
rect 17236 6866 17264 139431
rect 46940 77988 46992 77994
rect 46940 77930 46992 77936
rect 35900 73840 35952 73846
rect 35900 73782 35952 73788
rect 18602 69592 18658 69601
rect 18602 69527 18658 69536
rect 17958 53136 18014 53145
rect 17958 53071 18014 53080
rect 17316 31068 17368 31074
rect 17316 31010 17368 31016
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17328 4146 17356 31010
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 15948 480 15976 4082
rect 17040 3460 17092 3466
rect 17040 3402 17092 3408
rect 17052 480 17080 3402
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 53071
rect 18616 3466 18644 69527
rect 34520 68604 34572 68610
rect 34520 68546 34572 68552
rect 26238 68232 26294 68241
rect 26238 68167 26294 68176
rect 23478 61432 23534 61441
rect 23478 61367 23534 61376
rect 21364 60036 21416 60042
rect 21364 59978 21416 59984
rect 18604 3460 18656 3466
rect 18604 3402 18656 3408
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19444 480 19472 2994
rect 20640 480 20668 3402
rect 21376 3058 21404 59978
rect 23492 16574 23520 61367
rect 25502 57216 25558 57225
rect 25502 57151 25558 57160
rect 24860 29640 24912 29646
rect 24860 29582 24912 29588
rect 24872 16574 24900 29582
rect 23492 16546 24256 16574
rect 24872 16546 25360 16574
rect 21824 3664 21876 3670
rect 21824 3606 21876 3612
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 21836 480 21864 3606
rect 23020 3052 23072 3058
rect 23020 2994 23072 3000
rect 23032 480 23060 2994
rect 24228 480 24256 16546
rect 25332 480 25360 16546
rect 25516 3058 25544 57151
rect 25504 3052 25556 3058
rect 25504 2994 25556 3000
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 68167
rect 27620 62824 27672 62830
rect 27620 62766 27672 62772
rect 27632 16574 27660 62766
rect 30378 50280 30434 50289
rect 30378 50215 30434 50224
rect 30392 16574 30420 50215
rect 31760 35216 31812 35222
rect 31760 35158 31812 35164
rect 31772 16574 31800 35158
rect 27632 16546 27752 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 27724 480 27752 16546
rect 30104 14476 30156 14482
rect 30104 14418 30156 14424
rect 28908 6180 28960 6186
rect 28908 6122 28960 6128
rect 28920 480 28948 6122
rect 30116 480 30144 14418
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 33612 480 33640 3334
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 68546
rect 35164 65544 35216 65550
rect 35164 65486 35216 65492
rect 35176 3398 35204 65486
rect 35912 6914 35940 73782
rect 42800 71052 42852 71058
rect 42800 70994 42852 71000
rect 35992 69692 36044 69698
rect 35992 69634 36044 69640
rect 36004 16574 36032 69634
rect 40040 68400 40092 68406
rect 40040 68342 40092 68348
rect 39302 48920 39358 48929
rect 39302 48855 39358 48864
rect 36004 16546 36768 16574
rect 35912 6886 36032 6914
rect 35164 3392 35216 3398
rect 35164 3334 35216 3340
rect 36004 480 36032 6886
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 39316 3398 39344 48855
rect 40052 16574 40080 68342
rect 41418 54496 41474 54505
rect 41418 54431 41474 54440
rect 41432 16574 41460 54431
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 39580 3732 39632 3738
rect 39580 3674 39632 3680
rect 38384 3392 38436 3398
rect 38384 3334 38436 3340
rect 39304 3392 39356 3398
rect 39304 3334 39356 3340
rect 38396 480 38424 3334
rect 39592 480 39620 3674
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 70994
rect 44180 66904 44232 66910
rect 44180 66846 44232 66852
rect 44192 6914 44220 66846
rect 44270 47560 44326 47569
rect 44270 47495 44326 47504
rect 44284 16574 44312 47495
rect 45560 33788 45612 33794
rect 45560 33730 45612 33736
rect 45572 16574 45600 33730
rect 46952 16574 46980 77930
rect 66258 76664 66314 76673
rect 66258 76599 66314 76608
rect 52460 75200 52512 75206
rect 52460 75142 52512 75148
rect 48320 58676 48372 58682
rect 48320 58618 48372 58624
rect 48332 16574 48360 58618
rect 49698 46200 49754 46209
rect 49698 46135 49754 46144
rect 49712 16574 49740 46135
rect 44284 16546 45048 16574
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 44192 6886 44312 6914
rect 44284 480 44312 6886
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 52472 3398 52500 75142
rect 54482 73944 54538 73953
rect 54482 73879 54538 73888
rect 52552 65612 52604 65618
rect 52552 65554 52604 65560
rect 52460 3392 52512 3398
rect 52460 3334 52512 3340
rect 51356 3324 51408 3330
rect 51356 3266 51408 3272
rect 51368 480 51396 3266
rect 52564 480 52592 65554
rect 53380 3392 53432 3398
rect 53380 3334 53432 3340
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53392 354 53420 3334
rect 54496 3330 54524 73879
rect 60740 68672 60792 68678
rect 60740 68614 60792 68620
rect 59358 65648 59414 65657
rect 59358 65583 59414 65592
rect 57978 65512 58034 65521
rect 57978 65447 58034 65456
rect 57242 64288 57298 64297
rect 57242 64223 57298 64232
rect 56598 55992 56654 56001
rect 56598 55927 56654 55936
rect 56612 16574 56640 55927
rect 56612 16546 56824 16574
rect 54944 7608 54996 7614
rect 54944 7550 54996 7556
rect 54484 3324 54536 3330
rect 54484 3266 54536 3272
rect 54956 480 54984 7550
rect 56048 3392 56100 3398
rect 56048 3334 56100 3340
rect 56060 480 56088 3334
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 57256 3398 57284 64223
rect 57992 16574 58020 65447
rect 57992 16546 58480 16574
rect 57244 3392 57296 3398
rect 57244 3334 57296 3340
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 65583
rect 60752 6914 60780 68614
rect 60832 65680 60884 65686
rect 60832 65622 60884 65628
rect 60844 16574 60872 65622
rect 62120 60104 62172 60110
rect 62120 60046 62172 60052
rect 62132 16574 62160 60046
rect 63498 43480 63554 43489
rect 63498 43415 63554 43424
rect 63512 16574 63540 43415
rect 66272 16574 66300 76599
rect 67640 76560 67692 76566
rect 67640 76502 67692 76508
rect 60844 16546 61608 16574
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 66272 16546 66760 16574
rect 60752 6886 60872 6914
rect 60844 480 60872 6886
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 65524 3868 65576 3874
rect 65524 3810 65576 3816
rect 65536 480 65564 3810
rect 66732 480 66760 16546
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 76502
rect 88984 75948 89036 75954
rect 88984 75890 89036 75896
rect 71044 71120 71096 71126
rect 71044 71062 71096 71068
rect 70400 42084 70452 42090
rect 70400 42026 70452 42032
rect 70412 16574 70440 42026
rect 70412 16546 70992 16574
rect 69112 3800 69164 3806
rect 69112 3742 69164 3748
rect 69124 480 69152 3742
rect 70964 3482 70992 16546
rect 71056 3806 71084 71062
rect 85580 69828 85632 69834
rect 85580 69770 85632 69776
rect 77300 66972 77352 66978
rect 77300 66914 77352 66920
rect 75920 65748 75972 65754
rect 75920 65690 75972 65696
rect 72424 62892 72476 62898
rect 72424 62834 72476 62840
rect 71044 3800 71096 3806
rect 71044 3742 71096 3748
rect 70964 3454 71544 3482
rect 70308 2916 70360 2922
rect 70308 2858 70360 2864
rect 70320 480 70348 2858
rect 71516 480 71544 3454
rect 72436 2922 72464 62834
rect 75182 61568 75238 61577
rect 75182 61503 75238 61512
rect 74538 40624 74594 40633
rect 74538 40559 74594 40568
rect 74552 16574 74580 40559
rect 74552 16546 75040 16574
rect 73804 4140 73856 4146
rect 73804 4082 73856 4088
rect 72608 3868 72660 3874
rect 72608 3810 72660 3816
rect 72424 2916 72476 2922
rect 72424 2858 72476 2864
rect 72620 480 72648 3810
rect 73816 480 73844 4082
rect 75012 480 75040 16546
rect 75196 4146 75224 61503
rect 75184 4140 75236 4146
rect 75184 4082 75236 4088
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 65690
rect 77312 6914 77340 66914
rect 78680 65816 78732 65822
rect 78680 65758 78732 65764
rect 77392 39364 77444 39370
rect 77392 39306 77444 39312
rect 77404 16574 77432 39306
rect 78692 16574 78720 65758
rect 80058 57352 80114 57361
rect 80058 57287 80114 57296
rect 80072 16574 80100 57287
rect 84198 54632 84254 54641
rect 84198 54567 84254 54576
rect 81438 51776 81494 51785
rect 81438 51711 81494 51720
rect 81452 16574 81480 51711
rect 77404 16546 78168 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 77312 6886 77432 6914
rect 77404 480 77432 6886
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83280 3936 83332 3942
rect 83280 3878 83332 3884
rect 83292 480 83320 3878
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 54567
rect 85592 16574 85620 69770
rect 88340 64184 88392 64190
rect 88340 64126 88392 64132
rect 88352 16574 88380 64126
rect 85592 16546 86448 16574
rect 88352 16546 88932 16574
rect 85672 4004 85724 4010
rect 85672 3946 85724 3952
rect 85684 480 85712 3946
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 87512 10328 87564 10334
rect 87512 10270 87564 10276
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 10270
rect 88904 3482 88932 16546
rect 88996 4010 89024 75890
rect 89720 75472 89772 75478
rect 89720 75414 89772 75420
rect 89732 16574 89760 75414
rect 93124 65952 93176 65958
rect 93124 65894 93176 65900
rect 92478 53816 92534 53825
rect 92478 53751 92534 53760
rect 89732 16546 89944 16574
rect 88984 4004 89036 4010
rect 88984 3946 89036 3952
rect 88904 3454 89208 3482
rect 89180 480 89208 3454
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91560 3392 91612 3398
rect 91560 3334 91612 3340
rect 91572 480 91600 3334
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 53751
rect 93136 3398 93164 65894
rect 93858 58576 93914 58585
rect 93858 58511 93914 58520
rect 93872 16574 93900 58511
rect 95238 44840 95294 44849
rect 95238 44775 95294 44784
rect 95252 16574 95280 44775
rect 95896 33114 95924 153206
rect 96068 151088 96120 151094
rect 96068 151030 96120 151036
rect 95976 139596 96028 139602
rect 95976 139538 96028 139544
rect 95988 85542 96016 139538
rect 95976 85536 96028 85542
rect 95976 85478 96028 85484
rect 96080 79354 96108 151030
rect 96068 79348 96120 79354
rect 96068 79290 96120 79296
rect 96172 79234 96200 153954
rect 96080 79206 96200 79234
rect 96080 75750 96108 79206
rect 96160 79144 96212 79150
rect 96160 79086 96212 79092
rect 96172 77110 96200 79086
rect 96160 77104 96212 77110
rect 96160 77046 96212 77052
rect 96172 75954 96200 77046
rect 96160 75948 96212 75954
rect 96160 75890 96212 75896
rect 96068 75744 96120 75750
rect 96068 75686 96120 75692
rect 95976 73908 96028 73914
rect 95976 73850 96028 73856
rect 95884 33108 95936 33114
rect 95884 33050 95936 33056
rect 93872 16546 94728 16574
rect 95252 16546 95832 16574
rect 93124 3392 93176 3398
rect 93124 3334 93176 3340
rect 93952 3188 94004 3194
rect 93952 3130 94004 3136
rect 93964 480 93992 3130
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 95988 3194 96016 73850
rect 96264 41313 96292 154090
rect 96356 74526 96384 189722
rect 96448 76634 96476 193802
rect 97538 192536 97594 192545
rect 97448 192500 97500 192506
rect 97538 192471 97594 192480
rect 97448 192442 97500 192448
rect 97356 189848 97408 189854
rect 97356 189790 97408 189796
rect 97172 154080 97224 154086
rect 97172 154022 97224 154028
rect 96988 153944 97040 153950
rect 96988 153886 97040 153892
rect 96526 153776 96582 153785
rect 96526 153711 96582 153720
rect 96436 76628 96488 76634
rect 96436 76570 96488 76576
rect 96344 74520 96396 74526
rect 96344 74462 96396 74468
rect 96540 45554 96568 153711
rect 96620 72480 96672 72486
rect 96620 72422 96672 72428
rect 96448 45526 96568 45554
rect 96250 41304 96306 41313
rect 96250 41239 96306 41248
rect 96448 37233 96476 45526
rect 96526 41304 96582 41313
rect 96526 41239 96582 41248
rect 96540 40633 96568 41239
rect 96526 40624 96582 40633
rect 96526 40559 96582 40568
rect 96434 37224 96490 37233
rect 96434 37159 96490 37168
rect 96632 16574 96660 72422
rect 97000 67522 97028 153886
rect 97080 148436 97132 148442
rect 97080 148378 97132 148384
rect 97092 70378 97120 148378
rect 97080 70372 97132 70378
rect 97080 70314 97132 70320
rect 97184 68338 97212 154022
rect 97368 84194 97396 189790
rect 97276 84166 97396 84194
rect 97276 70281 97304 84166
rect 97356 75880 97408 75886
rect 97356 75822 97408 75828
rect 97368 75177 97396 75822
rect 97354 75168 97410 75177
rect 97354 75103 97410 75112
rect 97460 70922 97488 192442
rect 97448 70916 97500 70922
rect 97448 70858 97500 70864
rect 97262 70272 97318 70281
rect 97552 70242 97580 192471
rect 97644 73642 97672 199514
rect 97908 199504 97960 199510
rect 97908 199446 97960 199452
rect 97722 192672 97778 192681
rect 97722 192607 97778 192616
rect 97632 73636 97684 73642
rect 97632 73578 97684 73584
rect 97262 70207 97318 70216
rect 97540 70236 97592 70242
rect 97540 70178 97592 70184
rect 97172 68332 97224 68338
rect 97172 68274 97224 68280
rect 96988 67516 97040 67522
rect 96988 67458 97040 67464
rect 97736 66774 97764 192607
rect 97816 192568 97868 192574
rect 97816 192510 97868 192516
rect 97724 66768 97776 66774
rect 97724 66710 97776 66716
rect 97828 64870 97856 192510
rect 97816 64864 97868 64870
rect 97920 64841 97948 199446
rect 103150 199336 103206 199345
rect 103150 199271 103206 199280
rect 99286 199200 99342 199209
rect 99286 199135 99342 199144
rect 99196 191344 99248 191350
rect 99196 191286 99248 191292
rect 99104 191208 99156 191214
rect 99104 191150 99156 191156
rect 99012 191140 99064 191146
rect 99012 191082 99064 191088
rect 98920 187196 98972 187202
rect 98920 187138 98972 187144
rect 98736 187128 98788 187134
rect 98736 187070 98788 187076
rect 98644 151564 98696 151570
rect 98644 151506 98696 151512
rect 98552 151224 98604 151230
rect 98552 151166 98604 151172
rect 98460 148708 98512 148714
rect 98460 148650 98512 148656
rect 98472 71641 98500 148650
rect 98458 71632 98514 71641
rect 98458 71567 98514 71576
rect 98472 71233 98500 71567
rect 98458 71224 98514 71233
rect 98458 71159 98514 71168
rect 98564 70174 98592 151166
rect 98552 70168 98604 70174
rect 98552 70110 98604 70116
rect 97816 64806 97868 64812
rect 97906 64832 97962 64841
rect 97906 64767 97962 64776
rect 98656 60722 98684 151506
rect 98748 76945 98776 187070
rect 98828 186992 98880 186998
rect 98828 186934 98880 186940
rect 98734 76936 98790 76945
rect 98734 76871 98790 76880
rect 98748 76537 98776 76871
rect 98734 76528 98790 76537
rect 98734 76463 98790 76472
rect 98840 75818 98868 186934
rect 98828 75812 98880 75818
rect 98828 75754 98880 75760
rect 98932 74322 98960 187138
rect 99024 77178 99052 191082
rect 99012 77172 99064 77178
rect 99012 77114 99064 77120
rect 98920 74316 98972 74322
rect 98920 74258 98972 74264
rect 99116 71602 99144 191150
rect 99104 71596 99156 71602
rect 99104 71538 99156 71544
rect 99208 68542 99236 191286
rect 99300 69018 99328 199135
rect 100574 195256 100630 195265
rect 100574 195191 100630 195200
rect 100484 194132 100536 194138
rect 100484 194074 100536 194080
rect 100300 187468 100352 187474
rect 100300 187410 100352 187416
rect 100024 151428 100076 151434
rect 100024 151370 100076 151376
rect 99840 149728 99892 149734
rect 99840 149670 99892 149676
rect 99852 79762 99880 149670
rect 99932 148572 99984 148578
rect 99932 148514 99984 148520
rect 99840 79756 99892 79762
rect 99840 79698 99892 79704
rect 99944 78674 99972 148514
rect 99932 78668 99984 78674
rect 99932 78610 99984 78616
rect 99944 76378 99972 78610
rect 99852 76350 99972 76378
rect 99380 75744 99432 75750
rect 99380 75686 99432 75692
rect 99288 69012 99340 69018
rect 99288 68954 99340 68960
rect 99196 68536 99248 68542
rect 99196 68478 99248 68484
rect 98644 60716 98696 60722
rect 98644 60658 98696 60664
rect 98000 60648 98052 60654
rect 98000 60590 98052 60596
rect 98012 16574 98040 60590
rect 98656 60042 98684 60658
rect 98644 60036 98696 60042
rect 98644 59978 98696 59984
rect 99392 16574 99420 75686
rect 99852 68610 99880 76350
rect 99932 75948 99984 75954
rect 99932 75890 99984 75896
rect 99944 73001 99972 75890
rect 99930 72992 99986 73001
rect 99930 72927 99986 72936
rect 99840 68604 99892 68610
rect 99840 68546 99892 68552
rect 100036 67386 100064 151370
rect 100116 151360 100168 151366
rect 100116 151302 100168 151308
rect 100024 67380 100076 67386
rect 100024 67322 100076 67328
rect 100128 67318 100156 151302
rect 100206 151056 100262 151065
rect 100206 150991 100262 151000
rect 100220 70394 100248 150991
rect 100312 75410 100340 187410
rect 100392 187332 100444 187338
rect 100392 187274 100444 187280
rect 100300 75404 100352 75410
rect 100300 75346 100352 75352
rect 100220 70366 100340 70394
rect 100116 67312 100168 67318
rect 100116 67254 100168 67260
rect 100312 62121 100340 70366
rect 100404 67250 100432 187274
rect 100496 75954 100524 194074
rect 100484 75948 100536 75954
rect 100484 75890 100536 75896
rect 100484 75744 100536 75750
rect 100484 75686 100536 75692
rect 100496 75342 100524 75686
rect 100484 75336 100536 75342
rect 100484 75278 100536 75284
rect 100392 67244 100444 67250
rect 100392 67186 100444 67192
rect 100588 63510 100616 195191
rect 101680 192908 101732 192914
rect 101680 192850 101732 192856
rect 100666 191040 100722 191049
rect 100666 190975 100722 190984
rect 100576 63504 100628 63510
rect 100576 63446 100628 63452
rect 100588 62830 100616 63446
rect 100576 62824 100628 62830
rect 100576 62766 100628 62772
rect 100298 62112 100354 62121
rect 100298 62047 100354 62056
rect 100312 61441 100340 62047
rect 100298 61432 100354 61441
rect 100298 61367 100354 61376
rect 100680 50969 100708 190975
rect 101404 151700 101456 151706
rect 101404 151642 101456 151648
rect 101312 151156 101364 151162
rect 101312 151098 101364 151104
rect 101218 138680 101274 138689
rect 101218 138615 101274 138624
rect 101232 77246 101260 138615
rect 101324 78062 101352 151098
rect 101312 78056 101364 78062
rect 101312 77998 101364 78004
rect 101220 77240 101272 77246
rect 101220 77182 101272 77188
rect 101312 76084 101364 76090
rect 101312 76026 101364 76032
rect 101324 73658 101352 76026
rect 101416 75970 101444 151642
rect 101496 151292 101548 151298
rect 101496 151234 101548 151240
rect 101508 76090 101536 151234
rect 101586 148336 101642 148345
rect 101586 148271 101642 148280
rect 101496 76084 101548 76090
rect 101496 76026 101548 76032
rect 101416 75942 101536 75970
rect 101508 74118 101536 75942
rect 101496 74112 101548 74118
rect 101496 74054 101548 74060
rect 101508 73846 101536 74054
rect 101496 73840 101548 73846
rect 101496 73782 101548 73788
rect 101324 73630 101536 73658
rect 101508 71534 101536 73630
rect 101496 71528 101548 71534
rect 101496 71470 101548 71476
rect 101508 71058 101536 71470
rect 101496 71052 101548 71058
rect 101496 70994 101548 71000
rect 100760 59356 100812 59362
rect 100760 59298 100812 59304
rect 100772 58682 100800 59298
rect 100760 58676 100812 58682
rect 100760 58618 100812 58624
rect 99470 50960 99526 50969
rect 99470 50895 99526 50904
rect 100666 50960 100722 50969
rect 100666 50895 100722 50904
rect 99484 50289 99512 50895
rect 99470 50280 99526 50289
rect 99470 50215 99526 50224
rect 100758 49600 100814 49609
rect 100758 49535 100814 49544
rect 100772 48929 100800 49535
rect 100758 48920 100814 48929
rect 100758 48855 100814 48864
rect 101600 46889 101628 148271
rect 101692 69902 101720 192850
rect 101772 192840 101824 192846
rect 101772 192782 101824 192788
rect 101680 69896 101732 69902
rect 101680 69838 101732 69844
rect 101692 69698 101720 69838
rect 101680 69692 101732 69698
rect 101680 69634 101732 69640
rect 101784 66910 101812 192782
rect 103060 191276 103112 191282
rect 103060 191218 103112 191224
rect 101864 189984 101916 189990
rect 101864 189926 101916 189932
rect 101772 66904 101824 66910
rect 101772 66846 101824 66852
rect 101876 59362 101904 189926
rect 101956 187536 102008 187542
rect 101956 187478 102008 187484
rect 101864 59356 101916 59362
rect 101864 59298 101916 59304
rect 101968 55185 101996 187478
rect 102046 187096 102102 187105
rect 102046 187031 102102 187040
rect 101954 55176 102010 55185
rect 101954 55111 102010 55120
rect 101968 54505 101996 55111
rect 101954 54496 102010 54505
rect 101954 54431 102010 54440
rect 102060 49609 102088 187031
rect 102784 151632 102836 151638
rect 102784 151574 102836 151580
rect 102598 138816 102654 138825
rect 102598 138751 102654 138760
rect 102612 71670 102640 138751
rect 102690 112432 102746 112441
rect 102690 112367 102746 112376
rect 102600 71664 102652 71670
rect 102600 71606 102652 71612
rect 102046 49600 102102 49609
rect 102046 49535 102102 49544
rect 100758 46880 100814 46889
rect 100758 46815 100814 46824
rect 101586 46880 101642 46889
rect 101586 46815 101642 46824
rect 100772 46209 100800 46815
rect 100758 46200 100814 46209
rect 100758 46135 100814 46144
rect 102704 44169 102732 112367
rect 102796 80442 102824 151574
rect 102968 151496 103020 151502
rect 102968 151438 103020 151444
rect 102876 147144 102928 147150
rect 102876 147086 102928 147092
rect 102784 80436 102836 80442
rect 102784 80378 102836 80384
rect 102888 75206 102916 147086
rect 102876 75200 102928 75206
rect 102876 75142 102928 75148
rect 102782 69864 102838 69873
rect 102782 69799 102838 69808
rect 102796 69601 102824 69799
rect 102782 69592 102838 69601
rect 102782 69527 102784 69536
rect 102836 69527 102838 69536
rect 102784 69498 102836 69504
rect 102796 69467 102824 69498
rect 102784 69080 102836 69086
rect 102784 69022 102836 69028
rect 102138 44160 102194 44169
rect 102138 44095 102194 44104
rect 102690 44160 102746 44169
rect 102690 44095 102746 44104
rect 102152 43489 102180 44095
rect 102138 43480 102194 43489
rect 102138 43415 102194 43424
rect 102138 37224 102194 37233
rect 102138 37159 102194 37168
rect 102152 36553 102180 37159
rect 102138 36544 102194 36553
rect 102138 36479 102194 36488
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 95976 3188 96028 3194
rect 95976 3130 96028 3136
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 102152 3398 102180 36479
rect 102232 4072 102284 4078
rect 102232 4014 102284 4020
rect 102140 3392 102192 3398
rect 102140 3334 102192 3340
rect 101036 3324 101088 3330
rect 101036 3266 101088 3272
rect 101048 480 101076 3266
rect 102244 480 102272 4014
rect 102796 3330 102824 69022
rect 102980 68814 103008 151438
rect 103072 76809 103100 191218
rect 103164 77926 103192 199271
rect 103336 194064 103388 194070
rect 103336 194006 103388 194012
rect 103244 190188 103296 190194
rect 103244 190130 103296 190136
rect 103152 77920 103204 77926
rect 103152 77862 103204 77868
rect 103058 76800 103114 76809
rect 103058 76735 103114 76744
rect 103150 68912 103206 68921
rect 103150 68847 103206 68856
rect 102968 68808 103020 68814
rect 102968 68750 103020 68756
rect 103164 68474 103192 68847
rect 103152 68468 103204 68474
rect 103152 68410 103204 68416
rect 103164 68241 103192 68410
rect 103150 68232 103206 68241
rect 103150 68167 103206 68176
rect 103256 66094 103284 190130
rect 103348 68678 103376 194006
rect 104348 193928 104400 193934
rect 104348 193870 104400 193876
rect 103426 192944 103482 192953
rect 103426 192879 103482 192888
rect 103336 68672 103388 68678
rect 103336 68614 103388 68620
rect 103348 68406 103376 68614
rect 103336 68400 103388 68406
rect 103336 68342 103388 68348
rect 103440 67538 103468 192879
rect 104164 148980 104216 148986
rect 104164 148922 104216 148928
rect 104072 147076 104124 147082
rect 104072 147018 104124 147024
rect 103978 113792 104034 113801
rect 103978 113727 104034 113736
rect 103992 81161 104020 113727
rect 103978 81152 104034 81161
rect 103978 81087 104034 81096
rect 104084 78130 104112 147018
rect 104072 78124 104124 78130
rect 104072 78066 104124 78072
rect 104176 75750 104204 148922
rect 104256 140072 104308 140078
rect 104256 140014 104308 140020
rect 104164 75744 104216 75750
rect 104164 75686 104216 75692
rect 103348 67510 103468 67538
rect 103244 66088 103296 66094
rect 103244 66030 103296 66036
rect 103348 65550 103376 67510
rect 103428 66088 103480 66094
rect 103428 66030 103480 66036
rect 103440 65618 103468 66030
rect 104176 65754 104204 75686
rect 104164 65748 104216 65754
rect 104164 65690 104216 65696
rect 104268 65634 104296 140014
rect 104360 75478 104388 193870
rect 104440 187264 104492 187270
rect 104440 187206 104492 187212
rect 104348 75472 104400 75478
rect 104348 75414 104400 75420
rect 104452 67182 104480 187206
rect 104544 78266 104572 199582
rect 105728 198212 105780 198218
rect 105728 198154 105780 198160
rect 105636 198076 105688 198082
rect 105636 198018 105688 198024
rect 104716 196648 104768 196654
rect 104716 196590 104768 196596
rect 104622 195392 104678 195401
rect 104622 195327 104678 195336
rect 104532 78260 104584 78266
rect 104532 78202 104584 78208
rect 104636 72593 104664 195327
rect 104728 73137 104756 196590
rect 104808 191548 104860 191554
rect 104808 191490 104860 191496
rect 104714 73128 104770 73137
rect 104714 73063 104770 73072
rect 104622 72584 104678 72593
rect 104622 72519 104678 72528
rect 104440 67176 104492 67182
rect 104440 67118 104492 67124
rect 104452 66978 104480 67118
rect 104440 66972 104492 66978
rect 104440 66914 104492 66920
rect 104438 66192 104494 66201
rect 104438 66127 104440 66136
rect 104492 66127 104494 66136
rect 104440 66098 104492 66104
rect 104452 65657 104480 66098
rect 104728 65822 104756 73063
rect 104716 65816 104768 65822
rect 104716 65758 104768 65764
rect 103428 65612 103480 65618
rect 103428 65554 103480 65560
rect 104176 65606 104296 65634
rect 104438 65648 104494 65657
rect 103336 65544 103388 65550
rect 103336 65486 103388 65492
rect 104176 64802 104204 65606
rect 104438 65583 104494 65592
rect 104164 64796 104216 64802
rect 104164 64738 104216 64744
rect 103796 64728 103848 64734
rect 103796 64670 103848 64676
rect 103808 64297 103836 64670
rect 103980 64660 104032 64666
rect 103980 64602 104032 64608
rect 103794 64288 103850 64297
rect 103794 64223 103850 64232
rect 103992 64161 104020 64602
rect 104176 64190 104204 64738
rect 104164 64184 104216 64190
rect 103978 64152 104034 64161
rect 104164 64126 104216 64132
rect 103978 64087 104034 64096
rect 104820 63442 104848 191490
rect 105542 189680 105598 189689
rect 105542 189615 105598 189624
rect 105360 147280 105412 147286
rect 105360 147222 105412 147228
rect 105174 81424 105230 81433
rect 105174 81359 105230 81368
rect 105188 80850 105216 81359
rect 105176 80844 105228 80850
rect 105176 80786 105228 80792
rect 105372 76906 105400 147222
rect 105452 146940 105504 146946
rect 105452 146882 105504 146888
rect 105360 76900 105412 76906
rect 105360 76842 105412 76848
rect 105372 76566 105400 76842
rect 105360 76560 105412 76566
rect 105360 76502 105412 76508
rect 104898 71088 104954 71097
rect 104898 71023 104900 71032
rect 104952 71023 104954 71032
rect 104900 70994 104952 71000
rect 104348 63436 104400 63442
rect 104348 63378 104400 63384
rect 104808 63436 104860 63442
rect 104808 63378 104860 63384
rect 104360 62898 104388 63378
rect 104348 62892 104400 62898
rect 104348 62834 104400 62840
rect 103520 62756 103572 62762
rect 103520 62698 103572 62704
rect 103532 16574 103560 62698
rect 105464 53825 105492 146882
rect 105556 72282 105584 189615
rect 105648 89146 105676 198018
rect 105636 89140 105688 89146
rect 105636 89082 105688 89088
rect 105740 89026 105768 198154
rect 107384 197056 107436 197062
rect 107384 196998 107436 197004
rect 107292 196716 107344 196722
rect 107292 196658 107344 196664
rect 105820 195560 105872 195566
rect 105820 195502 105872 195508
rect 105648 88998 105768 89026
rect 105648 77994 105676 88998
rect 105728 88936 105780 88942
rect 105728 88878 105780 88884
rect 105636 77988 105688 77994
rect 105636 77930 105688 77936
rect 105648 77586 105676 77930
rect 105740 77654 105768 88878
rect 105728 77648 105780 77654
rect 105728 77590 105780 77596
rect 105636 77580 105688 77586
rect 105636 77522 105688 77528
rect 105544 72276 105596 72282
rect 105544 72218 105596 72224
rect 105556 69086 105584 72218
rect 105544 69080 105596 69086
rect 105544 69022 105596 69028
rect 105740 65686 105768 77590
rect 105832 69834 105860 195502
rect 106002 191312 106058 191321
rect 106002 191247 106058 191256
rect 105912 187400 105964 187406
rect 105912 187342 105964 187348
rect 105820 69828 105872 69834
rect 105820 69770 105872 69776
rect 105728 65680 105780 65686
rect 105728 65622 105780 65628
rect 105924 60654 105952 187342
rect 106016 61577 106044 191247
rect 106096 190256 106148 190262
rect 106096 190198 106148 190204
rect 106002 61568 106058 61577
rect 106002 61503 106058 61512
rect 105912 60648 105964 60654
rect 105912 60590 105964 60596
rect 106108 60586 106136 190198
rect 107198 190088 107254 190097
rect 107198 190023 107254 190032
rect 107014 189952 107070 189961
rect 107014 189887 107070 189896
rect 106186 187640 106242 187649
rect 106186 187575 106242 187584
rect 105820 60580 105872 60586
rect 105820 60522 105872 60528
rect 106096 60580 106148 60586
rect 106096 60522 106148 60528
rect 105832 60110 105860 60522
rect 105820 60104 105872 60110
rect 105820 60046 105872 60052
rect 106200 57905 106228 187575
rect 106924 187060 106976 187066
rect 106924 187002 106976 187008
rect 106740 148232 106792 148238
rect 106740 148174 106792 148180
rect 106752 77994 106780 148174
rect 106830 138952 106886 138961
rect 106830 138887 106886 138896
rect 106740 77988 106792 77994
rect 106740 77930 106792 77936
rect 106278 73944 106334 73953
rect 106278 73879 106334 73888
rect 106292 73846 106320 73879
rect 106280 73840 106332 73846
rect 106280 73782 106332 73788
rect 106280 68332 106332 68338
rect 106280 68274 106332 68280
rect 106186 57896 106242 57905
rect 106186 57831 106242 57840
rect 105450 53816 105506 53825
rect 105450 53751 105506 53760
rect 106292 16574 106320 68274
rect 106844 62082 106872 138887
rect 106936 79558 106964 187002
rect 106924 79552 106976 79558
rect 106924 79494 106976 79500
rect 107028 78198 107056 189887
rect 107106 189816 107162 189825
rect 107106 189751 107162 189760
rect 107016 78192 107068 78198
rect 107016 78134 107068 78140
rect 107016 75268 107068 75274
rect 107016 75210 107068 75216
rect 106924 67040 106976 67046
rect 106924 66982 106976 66988
rect 106832 62076 106884 62082
rect 106832 62018 106884 62024
rect 103532 16546 104112 16574
rect 106292 16546 106504 16574
rect 103336 3392 103388 3398
rect 103336 3334 103388 3340
rect 102784 3324 102836 3330
rect 102784 3266 102836 3272
rect 103348 480 103376 3334
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105728 3392 105780 3398
rect 105728 3334 105780 3340
rect 105740 480 105768 3334
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 106936 3398 106964 66982
rect 107028 65958 107056 75210
rect 107120 73914 107148 189751
rect 107108 73908 107160 73914
rect 107108 73850 107160 73856
rect 107212 69494 107240 190023
rect 107304 72486 107332 196658
rect 107292 72480 107344 72486
rect 107292 72422 107344 72428
rect 107396 71126 107424 196998
rect 107476 191480 107528 191486
rect 107476 191422 107528 191428
rect 107488 75274 107516 191422
rect 107476 75268 107528 75274
rect 107476 75210 107528 75216
rect 107384 71120 107436 71126
rect 107384 71062 107436 71068
rect 107200 69488 107252 69494
rect 107200 69430 107252 69436
rect 107580 66978 107608 200398
rect 108396 198008 108448 198014
rect 108396 197950 108448 197956
rect 108304 194200 108356 194206
rect 108304 194142 108356 194148
rect 108212 192704 108264 192710
rect 108212 192646 108264 192652
rect 108120 189916 108172 189922
rect 108120 189858 108172 189864
rect 108028 79484 108080 79490
rect 108028 79426 108080 79432
rect 107752 75404 107804 75410
rect 107752 75346 107804 75352
rect 107764 75206 107792 75346
rect 107752 75200 107804 75206
rect 107752 75142 107804 75148
rect 108040 71330 108068 79426
rect 108132 79257 108160 189858
rect 108224 79354 108252 192646
rect 108212 79348 108264 79354
rect 108212 79290 108264 79296
rect 108118 79248 108174 79257
rect 108118 79183 108174 79192
rect 108316 78334 108344 194142
rect 108408 79422 108436 197950
rect 108488 195832 108540 195838
rect 108488 195774 108540 195780
rect 108396 79416 108448 79422
rect 108396 79358 108448 79364
rect 108304 78328 108356 78334
rect 108304 78270 108356 78276
rect 107660 71324 107712 71330
rect 107660 71266 107712 71272
rect 108028 71324 108080 71330
rect 108028 71266 108080 71272
rect 107568 66972 107620 66978
rect 107568 66914 107620 66920
rect 107016 65952 107068 65958
rect 107016 65894 107068 65900
rect 107672 16574 107700 71266
rect 108316 62762 108344 78270
rect 108500 75070 108528 195774
rect 108672 194336 108724 194342
rect 108672 194278 108724 194284
rect 108580 192772 108632 192778
rect 108580 192714 108632 192720
rect 108488 75064 108540 75070
rect 108488 75006 108540 75012
rect 108592 70106 108620 192714
rect 108684 79490 108712 194278
rect 108764 193996 108816 194002
rect 108764 193938 108816 193944
rect 108672 79484 108724 79490
rect 108672 79426 108724 79432
rect 108670 79248 108726 79257
rect 108670 79183 108726 79192
rect 108684 71738 108712 79183
rect 108672 71732 108724 71738
rect 108672 71674 108724 71680
rect 108580 70100 108632 70106
rect 108580 70042 108632 70048
rect 108776 68746 108804 193938
rect 108856 191616 108908 191622
rect 108856 191558 108908 191564
rect 108764 68740 108816 68746
rect 108764 68682 108816 68688
rect 108868 62830 108896 191558
rect 108960 70038 108988 200534
rect 109684 194268 109736 194274
rect 109684 194210 109736 194216
rect 109592 147348 109644 147354
rect 109592 147290 109644 147296
rect 109408 147008 109460 147014
rect 109408 146950 109460 146956
rect 108948 70032 109000 70038
rect 108948 69974 109000 69980
rect 109420 67046 109448 146950
rect 109498 123448 109554 123457
rect 109498 123383 109554 123392
rect 109512 80918 109540 123383
rect 109500 80912 109552 80918
rect 109500 80854 109552 80860
rect 109604 77858 109632 147290
rect 109696 79626 109724 194210
rect 109788 144498 109816 262618
rect 110328 198144 110380 198150
rect 110328 198086 110380 198092
rect 109958 196616 110014 196625
rect 109958 196551 110014 196560
rect 109868 195628 109920 195634
rect 109868 195570 109920 195576
rect 109776 144492 109828 144498
rect 109776 144434 109828 144440
rect 109684 79620 109736 79626
rect 109684 79562 109736 79568
rect 109592 77852 109644 77858
rect 109592 77794 109644 77800
rect 109880 72758 109908 195570
rect 109868 72752 109920 72758
rect 109868 72694 109920 72700
rect 109972 72350 110000 196551
rect 110236 195696 110288 195702
rect 110236 195638 110288 195644
rect 110144 190120 110196 190126
rect 110144 190062 110196 190068
rect 110052 190052 110104 190058
rect 110052 189994 110104 190000
rect 109960 72344 110012 72350
rect 109960 72286 110012 72292
rect 109408 67040 109460 67046
rect 109408 66982 109460 66988
rect 110064 66230 110092 189994
rect 110052 66224 110104 66230
rect 110156 66201 110184 190062
rect 110248 69902 110276 195638
rect 110236 69896 110288 69902
rect 110236 69838 110288 69844
rect 110052 66166 110104 66172
rect 110142 66192 110198 66201
rect 110142 66127 110198 66136
rect 110340 65958 110368 198086
rect 111248 195356 111300 195362
rect 111248 195298 111300 195304
rect 111156 152516 111208 152522
rect 111156 152458 111208 152464
rect 110788 148912 110840 148918
rect 110788 148854 110840 148860
rect 110696 147212 110748 147218
rect 110696 147154 110748 147160
rect 110328 65952 110380 65958
rect 110708 65929 110736 147154
rect 110800 68406 110828 148854
rect 111064 148776 111116 148782
rect 111064 148718 111116 148724
rect 110972 146124 111024 146130
rect 110972 146066 111024 146072
rect 110880 144764 110932 144770
rect 110880 144706 110932 144712
rect 110892 72418 110920 144706
rect 110880 72412 110932 72418
rect 110880 72354 110932 72360
rect 110984 69970 111012 146066
rect 111076 71262 111104 148718
rect 111168 75177 111196 152458
rect 111260 78946 111288 195298
rect 111340 195288 111392 195294
rect 111340 195230 111392 195236
rect 111352 79286 111380 195230
rect 111444 145994 111472 262783
rect 111432 145988 111484 145994
rect 111432 145930 111484 145936
rect 111536 144634 111564 263570
rect 113824 263016 113876 263022
rect 113824 262958 113876 262964
rect 112352 262948 112404 262954
rect 112352 262890 112404 262896
rect 111708 196988 111760 196994
rect 111708 196930 111760 196936
rect 111616 196784 111668 196790
rect 111616 196726 111668 196732
rect 111524 144628 111576 144634
rect 111524 144570 111576 144576
rect 111340 79280 111392 79286
rect 111340 79222 111392 79228
rect 111248 78940 111300 78946
rect 111248 78882 111300 78888
rect 111246 77208 111302 77217
rect 111246 77143 111302 77152
rect 111260 76566 111288 77143
rect 111628 76974 111656 196726
rect 111616 76968 111668 76974
rect 111616 76910 111668 76916
rect 111248 76560 111300 76566
rect 111248 76502 111300 76508
rect 111154 75168 111210 75177
rect 111154 75103 111210 75112
rect 111064 71256 111116 71262
rect 111064 71198 111116 71204
rect 110972 69964 111024 69970
rect 110972 69906 111024 69912
rect 110788 68400 110840 68406
rect 110788 68342 110840 68348
rect 110328 65894 110380 65900
rect 110694 65920 110750 65929
rect 110694 65855 110750 65864
rect 108856 62824 108908 62830
rect 108856 62766 108908 62772
rect 108304 62756 108356 62762
rect 108304 62698 108356 62704
rect 109592 55208 109644 55214
rect 109592 55150 109644 55156
rect 109604 54641 109632 55150
rect 109590 54632 109646 54641
rect 109590 54567 109646 54576
rect 110420 50380 110472 50386
rect 110420 50322 110472 50328
rect 110432 16574 110460 50322
rect 107672 16546 108160 16574
rect 110432 16546 110552 16574
rect 106924 3392 106976 3398
rect 106924 3334 106976 3340
rect 108132 480 108160 16546
rect 109316 3392 109368 3398
rect 109316 3334 109368 3340
rect 109328 480 109356 3334
rect 110524 480 110552 16546
rect 111260 3398 111288 76502
rect 111720 69630 111748 196930
rect 112260 192636 112312 192642
rect 112260 192578 112312 192584
rect 112272 80753 112300 192578
rect 112364 148374 112392 262890
rect 112628 262812 112680 262818
rect 112628 262754 112680 262760
rect 112536 259684 112588 259690
rect 112536 259626 112588 259632
rect 112444 195492 112496 195498
rect 112444 195434 112496 195440
rect 112352 148368 112404 148374
rect 112352 148310 112404 148316
rect 112350 139360 112406 139369
rect 112350 139295 112406 139304
rect 112258 80744 112314 80753
rect 112364 80714 112392 139295
rect 112456 80782 112484 195434
rect 112548 144362 112576 259626
rect 112640 146198 112668 262754
rect 112812 259616 112864 259622
rect 112812 259558 112864 259564
rect 112720 192976 112772 192982
rect 112720 192918 112772 192924
rect 112628 146192 112680 146198
rect 112628 146134 112680 146140
rect 112536 144356 112588 144362
rect 112536 144298 112588 144304
rect 112628 141772 112680 141778
rect 112628 141714 112680 141720
rect 112534 138544 112590 138553
rect 112534 138479 112590 138488
rect 112444 80776 112496 80782
rect 112444 80718 112496 80724
rect 112258 80679 112314 80688
rect 112352 80708 112404 80714
rect 112352 80650 112404 80656
rect 112548 79082 112576 138479
rect 112536 79076 112588 79082
rect 112536 79018 112588 79024
rect 112640 76430 112668 141714
rect 112628 76424 112680 76430
rect 112628 76366 112680 76372
rect 112732 75585 112760 192918
rect 112824 142118 112852 259558
rect 113732 259548 113784 259554
rect 113732 259490 113784 259496
rect 112904 259480 112956 259486
rect 112904 259422 112956 259428
rect 112812 142112 112864 142118
rect 112812 142054 112864 142060
rect 112916 142050 112944 259422
rect 112996 199164 113048 199170
rect 112996 199106 113048 199112
rect 112904 142044 112956 142050
rect 112904 141986 112956 141992
rect 112812 141432 112864 141438
rect 112812 141374 112864 141380
rect 112718 75576 112774 75585
rect 112718 75511 112774 75520
rect 112442 72720 112498 72729
rect 112442 72655 112498 72664
rect 112456 72486 112484 72655
rect 111800 72480 111852 72486
rect 111800 72422 111852 72428
rect 112444 72480 112496 72486
rect 112444 72422 112496 72428
rect 111708 69624 111760 69630
rect 111708 69566 111760 69572
rect 111812 16574 111840 72422
rect 112824 71777 112852 141374
rect 112904 140548 112956 140554
rect 112904 140490 112956 140496
rect 112810 71768 112866 71777
rect 112810 71703 112866 71712
rect 112916 68610 112944 140490
rect 113008 75478 113036 199106
rect 113088 199028 113140 199034
rect 113088 198970 113140 198976
rect 113100 75682 113128 198970
rect 113546 147520 113602 147529
rect 113546 147455 113602 147464
rect 113178 138952 113234 138961
rect 113178 138887 113234 138896
rect 113192 138417 113220 138887
rect 113178 138408 113234 138417
rect 113178 138343 113234 138352
rect 113272 76492 113324 76498
rect 113272 76434 113324 76440
rect 113088 75676 113140 75682
rect 113088 75618 113140 75624
rect 112996 75472 113048 75478
rect 112996 75414 113048 75420
rect 113284 74633 113312 76434
rect 113270 74624 113326 74633
rect 113270 74559 113326 74568
rect 112904 68604 112956 68610
rect 112904 68546 112956 68552
rect 113180 65816 113232 65822
rect 113180 65758 113232 65764
rect 111812 16546 112392 16574
rect 111616 4004 111668 4010
rect 111616 3946 111668 3952
rect 111248 3392 111300 3398
rect 111248 3334 111300 3340
rect 111628 480 111656 3946
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 113192 3482 113220 65758
rect 113284 4078 113312 74559
rect 113560 70854 113588 147455
rect 113744 144090 113772 259490
rect 113836 146266 113864 262958
rect 114100 262880 114152 262886
rect 114100 262822 114152 262828
rect 113916 262744 113968 262750
rect 113916 262686 113968 262692
rect 113824 146260 113876 146266
rect 113824 146202 113876 146208
rect 113824 145648 113876 145654
rect 113824 145590 113876 145596
rect 113732 144084 113784 144090
rect 113732 144026 113784 144032
rect 113732 141500 113784 141506
rect 113732 141442 113784 141448
rect 113640 139460 113692 139466
rect 113640 139402 113692 139408
rect 113652 79490 113680 139402
rect 113744 79830 113772 141442
rect 113836 80889 113864 145590
rect 113928 143138 113956 262686
rect 114008 196852 114060 196858
rect 114008 196794 114060 196800
rect 113916 143132 113968 143138
rect 113916 143074 113968 143080
rect 113822 80880 113878 80889
rect 113822 80815 113878 80824
rect 113732 79824 113784 79830
rect 113732 79766 113784 79772
rect 113640 79484 113692 79490
rect 113640 79426 113692 79432
rect 114020 76770 114048 196794
rect 114112 141914 114140 262822
rect 114204 144838 114232 265134
rect 115480 263764 115532 263770
rect 115480 263706 115532 263712
rect 115388 262472 115440 262478
rect 115388 262414 115440 262420
rect 115296 261384 115348 261390
rect 115296 261326 115348 261332
rect 115204 259820 115256 259826
rect 115204 259762 115256 259768
rect 114468 199300 114520 199306
rect 114468 199242 114520 199248
rect 114284 199096 114336 199102
rect 114284 199038 114336 199044
rect 114192 144832 114244 144838
rect 114192 144774 114244 144780
rect 114192 143268 114244 143274
rect 114192 143210 114244 143216
rect 114100 141908 114152 141914
rect 114100 141850 114152 141856
rect 114100 140344 114152 140350
rect 114100 140286 114152 140292
rect 114008 76764 114060 76770
rect 114008 76706 114060 76712
rect 113548 70848 113600 70854
rect 113548 70790 113600 70796
rect 114112 68950 114140 140286
rect 114204 72214 114232 143210
rect 114296 77042 114324 199038
rect 114376 195424 114428 195430
rect 114376 195366 114428 195372
rect 114284 77036 114336 77042
rect 114284 76978 114336 76984
rect 114388 72962 114416 195366
rect 114480 75721 114508 199242
rect 114928 151768 114980 151774
rect 114928 151710 114980 151716
rect 114836 148504 114888 148510
rect 114836 148446 114888 148452
rect 114466 75712 114522 75721
rect 114466 75647 114522 75656
rect 114848 74458 114876 148446
rect 114940 81054 114968 151710
rect 115018 144528 115074 144537
rect 115018 144463 115074 144472
rect 115032 110673 115060 144463
rect 115216 142934 115244 259762
rect 115308 144702 115336 261326
rect 115296 144696 115348 144702
rect 115296 144638 115348 144644
rect 115400 143546 115428 262414
rect 115492 144906 115520 263706
rect 115572 263696 115624 263702
rect 115572 263638 115624 263644
rect 115480 144900 115532 144906
rect 115480 144842 115532 144848
rect 115388 143540 115440 143546
rect 115388 143482 115440 143488
rect 115204 142928 115256 142934
rect 115204 142870 115256 142876
rect 115480 141976 115532 141982
rect 115480 141918 115532 141924
rect 115112 141636 115164 141642
rect 115112 141578 115164 141584
rect 115018 110664 115074 110673
rect 115018 110599 115074 110608
rect 115020 110492 115072 110498
rect 115020 110434 115072 110440
rect 114928 81048 114980 81054
rect 114928 80990 114980 80996
rect 114836 74452 114888 74458
rect 114836 74394 114888 74400
rect 114376 72956 114428 72962
rect 114376 72898 114428 72904
rect 114192 72208 114244 72214
rect 114192 72150 114244 72156
rect 114560 71732 114612 71738
rect 114560 71674 114612 71680
rect 114100 68944 114152 68950
rect 114100 68886 114152 68892
rect 114572 16574 114600 71674
rect 115032 70242 115060 110434
rect 115124 79014 115152 141578
rect 115296 140208 115348 140214
rect 115296 140150 115348 140156
rect 115202 139224 115258 139233
rect 115202 139159 115258 139168
rect 115112 79008 115164 79014
rect 115112 78950 115164 78956
rect 115216 75449 115244 139159
rect 115202 75440 115258 75449
rect 115202 75375 115258 75384
rect 115308 71466 115336 140150
rect 115296 71460 115348 71466
rect 115296 71402 115348 71408
rect 115020 70236 115072 70242
rect 115020 70178 115072 70184
rect 115492 68882 115520 141918
rect 115584 141846 115612 263638
rect 118148 263084 118200 263090
rect 118148 263026 118200 263032
rect 116860 262404 116912 262410
rect 116860 262346 116912 262352
rect 116492 261248 116544 261254
rect 116492 261190 116544 261196
rect 116400 260092 116452 260098
rect 116400 260034 116452 260040
rect 115664 199368 115716 199374
rect 115664 199310 115716 199316
rect 115572 141840 115624 141846
rect 115572 141782 115624 141788
rect 115676 76838 115704 199310
rect 115848 199232 115900 199238
rect 115848 199174 115900 199180
rect 115756 198960 115808 198966
rect 115756 198902 115808 198908
rect 115664 76832 115716 76838
rect 115664 76774 115716 76780
rect 115768 73098 115796 198902
rect 115756 73092 115808 73098
rect 115756 73034 115808 73040
rect 115860 72826 115888 199174
rect 116412 145926 116440 260034
rect 116400 145920 116452 145926
rect 116400 145862 116452 145868
rect 116216 145852 116268 145858
rect 116216 145794 116268 145800
rect 116228 78985 116256 145794
rect 116308 145716 116360 145722
rect 116308 145658 116360 145664
rect 116320 79529 116348 145658
rect 116504 145518 116532 261190
rect 116676 260024 116728 260030
rect 116676 259966 116728 259972
rect 116584 259752 116636 259758
rect 116584 259694 116636 259700
rect 116492 145512 116544 145518
rect 116492 145454 116544 145460
rect 116596 142866 116624 259694
rect 116688 143002 116716 259966
rect 116768 191412 116820 191418
rect 116768 191354 116820 191360
rect 116676 142996 116728 143002
rect 116676 142938 116728 142944
rect 116584 142860 116636 142866
rect 116584 142802 116636 142808
rect 116400 141704 116452 141710
rect 116400 141646 116452 141652
rect 116306 79520 116362 79529
rect 116306 79455 116362 79464
rect 116412 79218 116440 141646
rect 116676 140412 116728 140418
rect 116676 140354 116728 140360
rect 116400 79212 116452 79218
rect 116400 79154 116452 79160
rect 116214 78976 116270 78985
rect 116214 78911 116270 78920
rect 116688 74225 116716 140354
rect 116674 74216 116730 74225
rect 116674 74151 116730 74160
rect 116780 74050 116808 191354
rect 116872 143342 116900 262346
rect 118056 261112 118108 261118
rect 118056 261054 118108 261060
rect 117872 260772 117924 260778
rect 117872 260714 117924 260720
rect 117228 200252 117280 200258
rect 117228 200194 117280 200200
rect 116952 199436 117004 199442
rect 116952 199378 117004 199384
rect 116860 143336 116912 143342
rect 116860 143278 116912 143284
rect 116860 141568 116912 141574
rect 116860 141510 116912 141516
rect 116768 74044 116820 74050
rect 116768 73986 116820 73992
rect 115848 72820 115900 72826
rect 115848 72762 115900 72768
rect 116872 71505 116900 141510
rect 116964 76702 116992 199378
rect 117136 198892 117188 198898
rect 117136 198834 117188 198840
rect 117044 196512 117096 196518
rect 117044 196454 117096 196460
rect 116952 76696 117004 76702
rect 116952 76638 117004 76644
rect 117056 72622 117084 196454
rect 117148 75206 117176 198834
rect 117136 75200 117188 75206
rect 117136 75142 117188 75148
rect 117240 72894 117268 200194
rect 117780 194540 117832 194546
rect 117780 194482 117832 194488
rect 117792 145790 117820 194482
rect 117884 150521 117912 260714
rect 117964 259888 118016 259894
rect 117964 259830 118016 259836
rect 117870 150512 117926 150521
rect 117870 150447 117926 150456
rect 117780 145784 117832 145790
rect 117780 145726 117832 145732
rect 117688 144152 117740 144158
rect 117688 144094 117740 144100
rect 117700 74089 117728 144094
rect 117884 142089 117912 150447
rect 117976 143070 118004 259830
rect 118068 143206 118096 261054
rect 118160 143410 118188 263026
rect 118240 195764 118292 195770
rect 118240 195706 118292 195712
rect 118148 143404 118200 143410
rect 118148 143346 118200 143352
rect 118056 143200 118108 143206
rect 118056 143142 118108 143148
rect 117964 143064 118016 143070
rect 117964 143006 118016 143012
rect 117870 142080 117926 142089
rect 117870 142015 117926 142024
rect 117964 140684 118016 140690
rect 117964 140626 118016 140632
rect 117872 140480 117924 140486
rect 117872 140422 117924 140428
rect 117780 140140 117832 140146
rect 117780 140082 117832 140088
rect 117792 81025 117820 140082
rect 117778 81016 117834 81025
rect 117778 80951 117834 80960
rect 117884 79121 117912 140422
rect 117870 79112 117926 79121
rect 117870 79047 117926 79056
rect 117976 74186 118004 140626
rect 118056 140616 118108 140622
rect 118056 140558 118108 140564
rect 117964 74180 118016 74186
rect 117964 74122 118016 74128
rect 117686 74080 117742 74089
rect 117686 74015 117742 74024
rect 118068 73778 118096 140558
rect 118056 73772 118108 73778
rect 118056 73714 118108 73720
rect 117228 72888 117280 72894
rect 117228 72830 117280 72836
rect 118252 72729 118280 195706
rect 118344 141545 118372 265202
rect 119988 265124 120040 265130
rect 119988 265066 120040 265072
rect 119896 265056 119948 265062
rect 119896 264998 119948 265004
rect 119710 262712 119766 262721
rect 119710 262647 119766 262656
rect 119528 261044 119580 261050
rect 119528 260986 119580 260992
rect 119252 260908 119304 260914
rect 119252 260850 119304 260856
rect 118608 200388 118660 200394
rect 118608 200330 118660 200336
rect 118516 200320 118568 200326
rect 118516 200262 118568 200268
rect 118424 198824 118476 198830
rect 118424 198766 118476 198772
rect 118330 141536 118386 141545
rect 118330 141471 118386 141480
rect 118332 141364 118384 141370
rect 118332 141306 118384 141312
rect 118238 72720 118294 72729
rect 118238 72655 118294 72664
rect 117044 72616 117096 72622
rect 117044 72558 117096 72564
rect 116858 71496 116914 71505
rect 116858 71431 116914 71440
rect 115480 68876 115532 68882
rect 115480 68818 115532 68824
rect 118344 68649 118372 141306
rect 118436 75313 118464 198766
rect 118422 75304 118478 75313
rect 118422 75239 118478 75248
rect 118528 73574 118556 200262
rect 118516 73568 118568 73574
rect 118516 73510 118568 73516
rect 118620 72554 118648 200330
rect 118700 198348 118752 198354
rect 118700 198290 118752 198296
rect 118712 80646 118740 198290
rect 119264 197198 119292 260850
rect 119436 260840 119488 260846
rect 119436 260782 119488 260788
rect 119344 259956 119396 259962
rect 119344 259898 119396 259904
rect 119252 197192 119304 197198
rect 119252 197134 119304 197140
rect 119356 154222 119384 259898
rect 119448 200122 119476 260782
rect 119436 200116 119488 200122
rect 119436 200058 119488 200064
rect 119540 196586 119568 260986
rect 119620 260976 119672 260982
rect 119620 260918 119672 260924
rect 119528 196580 119580 196586
rect 119528 196522 119580 196528
rect 119632 196314 119660 260918
rect 119620 196308 119672 196314
rect 119620 196250 119672 196256
rect 119528 193180 119580 193186
rect 119528 193122 119580 193128
rect 119436 193112 119488 193118
rect 119436 193054 119488 193060
rect 119344 154216 119396 154222
rect 119344 154158 119396 154164
rect 118976 151020 119028 151026
rect 118976 150962 119028 150968
rect 118884 149048 118936 149054
rect 118884 148990 118936 148996
rect 118792 148640 118844 148646
rect 118792 148582 118844 148588
rect 118700 80640 118752 80646
rect 118700 80582 118752 80588
rect 118608 72548 118660 72554
rect 118608 72490 118660 72496
rect 118804 69834 118832 148582
rect 118896 71194 118924 148990
rect 118884 71188 118936 71194
rect 118884 71130 118936 71136
rect 118792 69828 118844 69834
rect 118792 69770 118844 69776
rect 118330 68640 118386 68649
rect 118330 68575 118386 68584
rect 118988 68270 119016 150962
rect 119344 144288 119396 144294
rect 119344 144230 119396 144236
rect 119068 140888 119120 140894
rect 119068 140830 119120 140836
rect 119080 137970 119108 140830
rect 119252 140004 119304 140010
rect 119252 139946 119304 139952
rect 119068 137964 119120 137970
rect 119068 137906 119120 137912
rect 119158 137864 119214 137873
rect 119158 137799 119214 137808
rect 119172 80209 119200 137799
rect 119158 80200 119214 80209
rect 119158 80135 119214 80144
rect 119264 74254 119292 139946
rect 119356 75546 119384 144230
rect 119448 78538 119476 193054
rect 119436 78532 119488 78538
rect 119436 78474 119488 78480
rect 119540 78402 119568 193122
rect 119724 144430 119752 262647
rect 119804 198280 119856 198286
rect 119804 198222 119856 198228
rect 119712 144424 119764 144430
rect 119712 144366 119764 144372
rect 119816 79150 119844 198222
rect 119908 146062 119936 264998
rect 119896 146056 119948 146062
rect 119896 145998 119948 146004
rect 120000 144566 120028 265066
rect 120724 264988 120776 264994
rect 120724 264930 120776 264936
rect 120632 200660 120684 200666
rect 120632 200602 120684 200608
rect 120644 200462 120672 200602
rect 120632 200456 120684 200462
rect 120632 200398 120684 200404
rect 120540 197940 120592 197946
rect 120540 197882 120592 197888
rect 120356 196376 120408 196382
rect 120356 196318 120408 196324
rect 119988 144560 120040 144566
rect 119988 144502 120040 144508
rect 120080 80844 120132 80850
rect 120080 80786 120132 80792
rect 120092 80617 120120 80786
rect 120078 80608 120134 80617
rect 120078 80543 120134 80552
rect 119804 79144 119856 79150
rect 119804 79086 119856 79092
rect 119802 78432 119858 78441
rect 119528 78396 119580 78402
rect 119802 78367 119858 78376
rect 119528 78338 119580 78344
rect 119344 75540 119396 75546
rect 119344 75482 119396 75488
rect 119252 74248 119304 74254
rect 119252 74190 119304 74196
rect 118976 68264 119028 68270
rect 118976 68206 119028 68212
rect 117226 65512 117282 65521
rect 117226 65447 117282 65456
rect 115940 62824 115992 62830
rect 115940 62766 115992 62772
rect 116952 62824 117004 62830
rect 116952 62766 117004 62772
rect 115952 16574 115980 62766
rect 116964 61849 116992 62766
rect 117240 62082 117268 65447
rect 118988 64874 119016 68206
rect 119816 67454 119844 78367
rect 120368 70990 120396 196318
rect 120552 79694 120580 197882
rect 120736 194585 120764 264930
rect 120814 262440 120870 262449
rect 120814 262375 120870 262384
rect 120722 194576 120778 194585
rect 120828 194546 120856 262375
rect 120722 194511 120778 194520
rect 120816 194540 120868 194546
rect 120816 194482 120868 194488
rect 120816 190324 120868 190330
rect 120816 190266 120868 190272
rect 120632 142384 120684 142390
rect 120632 142326 120684 142332
rect 120644 138718 120672 142326
rect 120724 140276 120776 140282
rect 120724 140218 120776 140224
rect 120632 138712 120684 138718
rect 120632 138654 120684 138660
rect 120736 110498 120764 140218
rect 120828 138145 120856 190266
rect 120920 153882 120948 267706
rect 125968 263084 126020 263090
rect 125968 263026 126020 263032
rect 131120 263084 131172 263090
rect 131120 263026 131172 263032
rect 131764 263084 131816 263090
rect 131764 263026 131816 263032
rect 123208 262472 123260 262478
rect 123208 262414 123260 262420
rect 121368 262336 121420 262342
rect 121368 262278 121420 262284
rect 121276 261180 121328 261186
rect 121276 261122 121328 261128
rect 121184 198552 121236 198558
rect 121184 198494 121236 198500
rect 121092 198416 121144 198422
rect 121092 198358 121144 198364
rect 121000 197124 121052 197130
rect 121000 197066 121052 197072
rect 120908 153876 120960 153882
rect 120908 153818 120960 153824
rect 120908 148300 120960 148306
rect 120908 148242 120960 148248
rect 120814 138136 120870 138145
rect 120814 138071 120870 138080
rect 120724 110492 120776 110498
rect 120724 110434 120776 110440
rect 120724 81048 120776 81054
rect 120724 80990 120776 80996
rect 120630 80472 120686 80481
rect 120630 80407 120686 80416
rect 120540 79688 120592 79694
rect 120540 79630 120592 79636
rect 120644 72865 120672 80407
rect 120630 72856 120686 72865
rect 120630 72791 120686 72800
rect 120356 70984 120408 70990
rect 120356 70926 120408 70932
rect 120080 69488 120132 69494
rect 120080 69430 120132 69436
rect 119804 67448 119856 67454
rect 119804 67390 119856 67396
rect 120092 66910 120120 69430
rect 120736 69426 120764 80990
rect 120816 80912 120868 80918
rect 120816 80854 120868 80860
rect 120172 69420 120224 69426
rect 120172 69362 120224 69368
rect 120724 69420 120776 69426
rect 120724 69362 120776 69368
rect 120080 66904 120132 66910
rect 120080 66846 120132 66852
rect 120184 64874 120212 69362
rect 120724 66904 120776 66910
rect 120724 66846 120776 66852
rect 120264 66836 120316 66842
rect 120264 66778 120316 66784
rect 120276 65822 120304 66778
rect 120264 65816 120316 65822
rect 120264 65758 120316 65764
rect 118988 64846 119384 64874
rect 117228 62076 117280 62082
rect 117228 62018 117280 62024
rect 116950 61840 117006 61849
rect 116950 61775 117006 61784
rect 117240 60738 117268 62018
rect 117240 60710 117360 60738
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 113272 4072 113324 4078
rect 113272 4014 113324 4020
rect 113192 3454 114048 3482
rect 114020 480 114048 3454
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 60710
rect 119356 50386 119384 64846
rect 120092 64846 120212 64874
rect 119344 50380 119396 50386
rect 119344 50322 119396 50328
rect 120092 16574 120120 64846
rect 120092 16546 120672 16574
rect 119896 4072 119948 4078
rect 119896 4014 119948 4020
rect 118792 3052 118844 3058
rect 118792 2994 118844 3000
rect 118804 480 118832 2994
rect 119908 480 119936 4014
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 120736 3058 120764 66846
rect 120828 66842 120856 80854
rect 120920 71233 120948 148242
rect 121012 80850 121040 197066
rect 121000 80844 121052 80850
rect 121000 80786 121052 80792
rect 121104 80578 121132 198358
rect 121092 80572 121144 80578
rect 121092 80514 121144 80520
rect 121196 80510 121224 198494
rect 121288 197334 121316 261122
rect 121276 197328 121328 197334
rect 121276 197270 121328 197276
rect 121380 197266 121408 262278
rect 122840 260772 122892 260778
rect 122840 260714 122892 260720
rect 122852 259978 122880 260714
rect 123220 259978 123248 262414
rect 125600 261044 125652 261050
rect 125600 260986 125652 260992
rect 124312 260840 124364 260846
rect 124312 260782 124364 260788
rect 124324 259978 124352 260782
rect 125612 259978 125640 260986
rect 125980 259978 126008 263026
rect 130108 263016 130160 263022
rect 130108 262958 130160 262964
rect 128360 262948 128412 262954
rect 128360 262890 128412 262896
rect 127624 262404 127676 262410
rect 127624 262346 127676 262352
rect 127072 260976 127124 260982
rect 127072 260918 127124 260924
rect 127084 259978 127112 260918
rect 127636 259978 127664 262346
rect 128372 259978 128400 262890
rect 128728 262336 128780 262342
rect 128728 262278 128780 262284
rect 128740 259978 128768 262278
rect 130120 259978 130148 262958
rect 131132 262818 131160 263026
rect 131120 262812 131172 262818
rect 131120 262754 131172 262760
rect 131120 261112 131172 261118
rect 131120 261054 131172 261060
rect 130384 260908 130436 260914
rect 130384 260850 130436 260856
rect 130396 259978 130424 260850
rect 131132 259978 131160 261054
rect 131776 259978 131804 263026
rect 132040 262404 132092 262410
rect 132040 262346 132092 262352
rect 132052 261186 132080 262346
rect 132040 261180 132092 261186
rect 132040 261122 132092 261128
rect 132052 259978 132080 261122
rect 122852 259950 123004 259978
rect 123220 259950 123556 259978
rect 124324 259950 124660 259978
rect 125612 259950 125764 259978
rect 125980 259950 126316 259978
rect 127084 259950 127420 259978
rect 127636 259950 127972 259978
rect 128372 259950 128524 259978
rect 128740 259950 129076 259978
rect 130120 259950 130180 259978
rect 130396 259950 130732 259978
rect 131132 259950 131436 259978
rect 131776 259950 131836 259978
rect 132052 259950 132388 259978
rect 132512 259962 132540 271866
rect 134432 263764 134484 263770
rect 134432 263706 134484 263712
rect 133052 262744 133104 262750
rect 133052 262686 133104 262692
rect 133064 261322 133092 262686
rect 133052 261316 133104 261322
rect 133052 261258 133104 261264
rect 133064 259978 133092 261258
rect 134340 261248 134392 261254
rect 134340 261190 134392 261196
rect 134352 260370 134380 261190
rect 134340 260364 134392 260370
rect 134340 260306 134392 260312
rect 134352 259978 134380 260306
rect 132500 259956 132552 259962
rect 124864 259616 124916 259622
rect 123758 259584 123814 259593
rect 123814 259542 124108 259570
rect 131408 259593 131436 259950
rect 132940 259950 133092 259978
rect 133156 259962 133492 259978
rect 133144 259956 133492 259962
rect 132500 259898 132552 259904
rect 133196 259950 133492 259956
rect 134044 259950 134380 259978
rect 134444 259978 134472 263706
rect 134536 262886 134564 324294
rect 134616 298172 134668 298178
rect 134616 298114 134668 298120
rect 134628 263770 134656 298114
rect 134616 263764 134668 263770
rect 134616 263706 134668 263712
rect 134524 262880 134576 262886
rect 134524 262822 134576 262828
rect 134800 262880 134852 262886
rect 134800 262822 134852 262828
rect 134812 259978 134840 262822
rect 135272 260273 135300 351902
rect 135904 311908 135956 311914
rect 135904 311850 135956 311856
rect 135916 265198 135944 311850
rect 137284 276684 137336 276690
rect 137284 276626 137336 276632
rect 135904 265192 135956 265198
rect 135904 265134 135956 265140
rect 135258 260264 135314 260273
rect 135258 260199 135314 260208
rect 135916 259978 135944 265134
rect 137296 263702 137324 276626
rect 137376 271244 137428 271250
rect 137376 271186 137428 271192
rect 137284 263696 137336 263702
rect 137284 263638 137336 263644
rect 137388 263634 137416 271186
rect 137560 263696 137612 263702
rect 137560 263638 137612 263644
rect 137376 263628 137428 263634
rect 137376 263570 137428 263576
rect 136224 260264 136280 260273
rect 136224 260199 136280 260208
rect 134444 259950 134596 259978
rect 134812 259950 135148 259978
rect 135700 259950 135944 259978
rect 136238 259964 136266 260199
rect 137388 260148 137416 263570
rect 137468 263492 137520 263498
rect 137468 263434 137520 263440
rect 137480 261390 137508 263434
rect 137468 261384 137520 261390
rect 137468 261326 137520 261332
rect 137204 260120 137416 260148
rect 137204 259978 137232 260120
rect 137480 259978 137508 261326
rect 136804 259950 137232 259978
rect 137356 259950 137508 259978
rect 137572 259978 137600 263638
rect 138676 262682 138704 430578
rect 138756 418192 138808 418198
rect 138756 418134 138808 418140
rect 138768 265266 138796 418134
rect 139412 267734 139440 484366
rect 140044 470620 140096 470626
rect 140044 470562 140096 470568
rect 140056 267734 140084 470562
rect 141424 278044 141476 278050
rect 141424 277986 141476 277992
rect 139412 267706 139716 267734
rect 140056 267706 140268 267734
rect 138756 265260 138808 265266
rect 138756 265202 138808 265208
rect 138664 262676 138716 262682
rect 138664 262618 138716 262624
rect 138676 259978 138704 262618
rect 137572 259950 137908 259978
rect 138460 259950 138704 259978
rect 138768 259978 138796 265202
rect 139492 264240 139544 264246
rect 139492 264182 139544 264188
rect 139400 260024 139452 260030
rect 138768 259950 139012 259978
rect 139504 259978 139532 264182
rect 139452 259972 139532 259978
rect 139400 259966 139532 259972
rect 139412 259950 139532 259966
rect 133144 259898 133196 259904
rect 139504 259842 139532 259950
rect 139688 259978 139716 267706
rect 140240 262585 140268 267706
rect 141332 265736 141384 265742
rect 141332 265678 141384 265684
rect 140226 262576 140282 262585
rect 140226 262511 140282 262520
rect 140240 259978 140268 262511
rect 139688 259950 140116 259978
rect 140240 259950 140668 259978
rect 139504 259814 139564 259842
rect 139688 259826 139716 259950
rect 140872 259888 140924 259894
rect 141344 259842 141372 265678
rect 141436 263809 141464 277986
rect 141422 263800 141478 263809
rect 141422 263735 141478 263744
rect 141436 259978 141464 263735
rect 141436 259950 141772 259978
rect 140924 259836 141372 259842
rect 140872 259830 141372 259836
rect 139676 259820 139728 259826
rect 140884 259814 141372 259830
rect 139676 259762 139728 259768
rect 142172 259690 142200 590650
rect 142436 563100 142488 563106
rect 142436 563042 142488 563048
rect 142250 262848 142306 262857
rect 142250 262783 142306 262792
rect 142264 259978 142292 262783
rect 142448 259978 142476 563042
rect 142804 524476 142856 524482
rect 142804 524418 142856 524424
rect 142816 262857 142844 524418
rect 142802 262848 142858 262857
rect 142802 262783 142858 262792
rect 143552 260273 143580 616830
rect 144184 576904 144236 576910
rect 144184 576846 144236 576852
rect 144196 265169 144224 576846
rect 145564 286340 145616 286346
rect 145564 286282 145616 286288
rect 144920 279472 144972 279478
rect 144920 279414 144972 279420
rect 143630 265160 143686 265169
rect 143630 265095 143686 265104
rect 144182 265160 144238 265169
rect 144182 265095 144238 265104
rect 143538 260264 143594 260273
rect 143538 260199 143594 260208
rect 143644 259978 143672 265095
rect 144504 260264 144560 260273
rect 144504 260199 144560 260208
rect 142264 259950 142324 259978
rect 142448 259950 142876 259978
rect 143644 259950 143980 259978
rect 144518 259964 144546 260199
rect 144932 260001 144960 279414
rect 145576 265033 145604 286282
rect 146208 268388 146260 268394
rect 146208 268330 146260 268336
rect 145562 265024 145618 265033
rect 145562 264959 145618 264968
rect 144918 259992 144974 260001
rect 142448 259758 142476 259950
rect 145576 259978 145604 264959
rect 146220 263673 146248 268330
rect 146206 263664 146262 263673
rect 146206 263599 146262 263608
rect 146220 260250 146248 263599
rect 146174 260222 146248 260250
rect 144974 259950 145084 259978
rect 145576 259950 145636 259978
rect 146174 259964 146202 260222
rect 146312 259978 146340 696934
rect 146944 683188 146996 683194
rect 146944 683130 146996 683136
rect 146956 265130 146984 683130
rect 147956 280832 148008 280838
rect 147956 280774 148008 280780
rect 147772 269816 147824 269822
rect 147772 269758 147824 269764
rect 146944 265124 146996 265130
rect 146944 265066 146996 265072
rect 146956 259978 146984 265066
rect 147784 260137 147812 269758
rect 147770 260128 147826 260137
rect 147968 260098 147996 280774
rect 148336 267734 148364 700266
rect 149704 660340 149756 660346
rect 149704 660282 149756 660288
rect 149060 271176 149112 271182
rect 149060 271118 149112 271124
rect 148336 267706 148548 267734
rect 148520 265062 148548 267706
rect 148508 265056 148560 265062
rect 148508 264998 148560 265004
rect 147770 260063 147826 260072
rect 147956 260092 148008 260098
rect 147784 259978 147812 260063
rect 147956 260034 148008 260040
rect 147968 259978 147996 260034
rect 148520 259978 148548 264998
rect 149072 259978 149100 271118
rect 149716 262721 149744 660282
rect 152464 371272 152516 371278
rect 152464 371214 152516 371220
rect 151084 287700 151136 287706
rect 151084 287642 151136 287648
rect 150438 281616 150494 281625
rect 150438 281551 150494 281560
rect 150452 267734 150480 281551
rect 150452 267706 151032 267734
rect 150716 264988 150768 264994
rect 150716 264930 150768 264936
rect 149702 262712 149758 262721
rect 149702 262647 149758 262656
rect 149716 259978 149744 262647
rect 150728 259978 150756 264930
rect 150900 263628 150952 263634
rect 150900 263570 150952 263576
rect 151004 263594 151032 267706
rect 151096 264994 151124 287642
rect 151820 282940 151872 282946
rect 151820 282882 151872 282888
rect 151832 267734 151860 282882
rect 151832 267706 152412 267734
rect 151084 264988 151136 264994
rect 151084 264930 151136 264936
rect 146312 259950 146740 259978
rect 146956 259950 147292 259978
rect 147784 259950 147844 259978
rect 147968 259950 148396 259978
rect 148520 259950 148948 259978
rect 149072 259950 149500 259978
rect 149716 259950 150052 259978
rect 150604 259950 150756 259978
rect 150912 259978 150940 263570
rect 151004 263566 151308 263594
rect 151280 259978 151308 263566
rect 152186 262848 152242 262857
rect 152186 262783 152242 262792
rect 152200 262449 152228 262783
rect 152186 262440 152242 262449
rect 152186 262375 152242 262384
rect 150912 259950 151156 259978
rect 151280 259950 151708 259978
rect 144918 259927 144974 259936
rect 144932 259867 144960 259927
rect 142436 259752 142488 259758
rect 146496 259729 146524 259950
rect 149256 259865 149284 259950
rect 149242 259856 149298 259865
rect 152200 259842 152228 262375
rect 152384 259978 152412 267706
rect 152476 265810 152504 371214
rect 152464 265804 152516 265810
rect 152464 265746 152516 265752
rect 153212 263702 153240 702406
rect 157340 700732 157392 700738
rect 157340 700674 157392 700680
rect 155960 700664 156012 700670
rect 155960 700606 156012 700612
rect 153290 289912 153346 289921
rect 153290 289847 153346 289856
rect 153200 263696 153252 263702
rect 153304 263673 153332 289847
rect 154580 284368 154632 284374
rect 154580 284310 154632 284316
rect 153384 274712 153436 274718
rect 153384 274654 153436 274660
rect 153200 263638 153252 263644
rect 153290 263664 153346 263673
rect 153290 263599 153346 263608
rect 153290 263528 153346 263537
rect 153200 263492 153252 263498
rect 153396 263498 153424 274654
rect 154396 266484 154448 266490
rect 154396 266426 154448 266432
rect 153290 263463 153346 263472
rect 153384 263492 153436 263498
rect 153200 263434 153252 263440
rect 153212 259978 153240 263434
rect 153304 260148 153332 263463
rect 153384 263434 153436 263440
rect 153304 260120 153516 260148
rect 153488 259978 153516 260120
rect 154408 259978 154436 266426
rect 154592 259978 154620 284310
rect 155868 262880 155920 262886
rect 155868 262822 155920 262828
rect 155880 259978 155908 262822
rect 155972 260273 156000 700606
rect 157248 700596 157300 700602
rect 157248 700538 157300 700544
rect 156052 273284 156104 273290
rect 156052 273226 156104 273232
rect 155958 260264 156014 260273
rect 155958 260199 156014 260208
rect 152384 259950 152812 259978
rect 153212 259950 153364 259978
rect 153488 259950 153916 259978
rect 154408 259950 154468 259978
rect 154592 259950 155020 259978
rect 155572 259950 155908 259978
rect 156064 259978 156092 273226
rect 157260 265062 157288 700538
rect 157248 265056 157300 265062
rect 157248 264998 157300 265004
rect 156648 260264 156704 260273
rect 157260 260250 157288 264998
rect 156648 260199 156704 260208
rect 157214 260222 157288 260250
rect 156064 259950 156124 259978
rect 152200 259814 152260 259842
rect 149242 259791 149298 259800
rect 146482 259720 146538 259729
rect 142436 259694 142488 259700
rect 143092 259690 143428 259706
rect 142160 259684 142212 259690
rect 142160 259626 142212 259632
rect 143080 259684 143428 259690
rect 143132 259678 143428 259684
rect 156662 259706 156690 260199
rect 157214 259964 157242 260222
rect 157352 260166 157380 700674
rect 160744 700528 160796 700534
rect 160744 700470 160796 700476
rect 157432 447840 157484 447846
rect 157432 447782 157484 447788
rect 157340 260160 157392 260166
rect 157340 260102 157392 260108
rect 157444 259978 157472 447782
rect 160100 275324 160152 275330
rect 160100 275266 160152 275272
rect 159364 273964 159416 273970
rect 159364 273906 159416 273912
rect 158720 265668 158772 265674
rect 158720 265610 158772 265616
rect 158732 263770 158760 265610
rect 158720 263764 158772 263770
rect 158720 263706 158772 263712
rect 159272 263764 159324 263770
rect 159272 263706 159324 263712
rect 158812 263696 158864 263702
rect 158812 263638 158864 263644
rect 158306 260160 158358 260166
rect 158306 260102 158358 260108
rect 158318 259978 158346 260102
rect 158824 259978 158852 263638
rect 159284 259978 159312 263706
rect 159376 262818 159404 273906
rect 159364 262812 159416 262818
rect 159364 262754 159416 262760
rect 159916 262812 159968 262818
rect 159916 262754 159968 262760
rect 159928 259978 159956 262754
rect 160112 260001 160140 275266
rect 160756 267734 160784 700470
rect 162216 700460 162268 700466
rect 162216 700402 162268 700408
rect 162124 700392 162176 700398
rect 162124 700334 162176 700340
rect 161480 683256 161532 683262
rect 161480 683198 161532 683204
rect 160756 267706 160876 267734
rect 160848 265198 160876 267706
rect 160836 265192 160888 265198
rect 160836 265134 160888 265140
rect 160098 259992 160154 260001
rect 157444 259950 158116 259978
rect 158318 259964 158668 259978
rect 158332 259950 158668 259964
rect 158824 259950 158884 259978
rect 159284 259950 159436 259978
rect 159928 259950 159988 259978
rect 158088 259758 158116 259950
rect 158076 259752 158128 259758
rect 156786 259720 156842 259729
rect 156662 259692 156786 259706
rect 156676 259678 156786 259692
rect 146482 259655 146538 259664
rect 158076 259694 158128 259700
rect 158640 259690 158668 259950
rect 160848 259978 160876 265134
rect 161492 260817 161520 683198
rect 162136 267734 162164 700334
rect 162044 267706 162164 267734
rect 162044 262585 162072 267706
rect 162228 262682 162256 700402
rect 163504 670744 163556 670750
rect 163504 670686 163556 670692
rect 163516 265130 163544 670686
rect 163596 656940 163648 656946
rect 163596 656882 163648 656888
rect 163504 265124 163556 265130
rect 163504 265066 163556 265072
rect 163410 263120 163466 263129
rect 163410 263055 163466 263064
rect 162216 262676 162268 262682
rect 162216 262618 162268 262624
rect 162030 262576 162086 262585
rect 162030 262511 162086 262520
rect 161478 260808 161534 260817
rect 161478 260743 161534 260752
rect 160540 259950 160876 259978
rect 160926 259992 160982 260001
rect 160098 259927 160154 259936
rect 162044 259978 162072 262511
rect 162228 260250 162256 262618
rect 163424 262449 163452 263055
rect 163410 262440 163466 262449
rect 163410 262375 163466 262384
rect 162674 260808 162730 260817
rect 162674 260743 162730 260752
rect 160982 259950 161092 259978
rect 161644 259950 162072 259978
rect 162182 260222 162256 260250
rect 162182 259964 162210 260222
rect 160926 259927 160982 259936
rect 162582 259856 162638 259865
rect 162688 259842 162716 260743
rect 163424 259978 163452 262375
rect 163300 259950 163452 259978
rect 163516 259978 163544 265066
rect 163608 263129 163636 656882
rect 164240 632120 164292 632126
rect 164240 632062 164292 632068
rect 163594 263120 163650 263129
rect 163594 263055 163650 263064
rect 164252 259978 164280 632062
rect 164884 618316 164936 618322
rect 164884 618258 164936 618264
rect 164896 265470 164924 618258
rect 164976 605872 165028 605878
rect 164976 605814 165028 605820
rect 164884 265464 164936 265470
rect 164884 265406 164936 265412
rect 164988 262954 165016 605814
rect 165620 579692 165672 579698
rect 165620 579634 165672 579640
rect 165436 265464 165488 265470
rect 165436 265406 165488 265412
rect 165448 264994 165476 265406
rect 165436 264988 165488 264994
rect 165436 264930 165488 264936
rect 164976 262948 165028 262954
rect 164976 262890 165028 262896
rect 164988 260250 165016 262890
rect 164942 260222 165016 260250
rect 164376 260128 164432 260137
rect 164376 260063 164432 260072
rect 164390 259978 164418 260063
rect 163516 259950 163852 259978
rect 164252 259964 164418 259978
rect 164942 259964 164970 260222
rect 165448 259978 165476 264930
rect 165632 259978 165660 579634
rect 167644 565888 167696 565894
rect 167644 565830 167696 565836
rect 165712 553444 165764 553450
rect 165712 553386 165764 553392
rect 165724 260166 165752 553386
rect 167000 527196 167052 527202
rect 167000 527138 167052 527144
rect 166632 260296 166684 260302
rect 166598 260244 166632 260250
rect 166598 260238 166684 260244
rect 166598 260222 166672 260238
rect 166598 260166 166626 260222
rect 165712 260160 165764 260166
rect 165712 260102 165764 260108
rect 166586 260160 166638 260166
rect 166586 260102 166638 260108
rect 164252 259950 164404 259964
rect 165448 259950 165508 259978
rect 165632 259962 166396 259978
rect 166598 259964 166626 260102
rect 167012 260098 167040 527138
rect 167276 501016 167328 501022
rect 167276 500958 167328 500964
rect 167288 260846 167316 500958
rect 167656 267734 167684 565830
rect 169772 447846 169800 702406
rect 202800 700670 202828 703520
rect 202788 700664 202840 700670
rect 202788 700606 202840 700612
rect 218992 700602 219020 703520
rect 218980 700596 219032 700602
rect 218980 700538 219032 700544
rect 185584 670744 185636 670750
rect 185584 670686 185636 670692
rect 182824 643136 182876 643142
rect 182824 643078 182876 643084
rect 181444 510672 181496 510678
rect 181444 510614 181496 510620
rect 170404 462392 170456 462398
rect 170404 462334 170456 462340
rect 169760 447840 169812 447846
rect 169760 447782 169812 447788
rect 169760 422340 169812 422346
rect 169760 422282 169812 422288
rect 169024 289128 169076 289134
rect 169024 289070 169076 289076
rect 167564 267706 167684 267734
rect 168380 267776 168432 267782
rect 168432 267724 168972 267734
rect 168380 267718 168972 267724
rect 168392 267706 168972 267718
rect 167564 265033 167592 267706
rect 168748 265260 168800 265266
rect 168748 265202 168800 265208
rect 167550 265024 167606 265033
rect 167550 264959 167606 264968
rect 167276 260840 167328 260846
rect 167276 260782 167328 260788
rect 167000 260092 167052 260098
rect 167000 260034 167052 260040
rect 167564 259978 167592 264959
rect 168196 260840 168248 260846
rect 168196 260782 168248 260788
rect 167690 260092 167742 260098
rect 167690 260034 167742 260040
rect 165632 259956 166408 259962
rect 165632 259950 166356 259956
rect 167164 259950 167592 259978
rect 167702 259964 167730 260034
rect 166356 259898 166408 259904
rect 168208 259842 168236 260782
rect 168760 259978 168788 265202
rect 168944 259978 168972 267706
rect 169036 265266 169064 289070
rect 169024 265260 169076 265266
rect 169024 265202 169076 265208
rect 169772 260166 169800 422282
rect 170220 265464 170272 265470
rect 170220 265406 170272 265412
rect 169760 260160 169812 260166
rect 169760 260102 169812 260108
rect 170232 259978 170260 265406
rect 170416 265334 170444 462334
rect 180064 456816 180116 456822
rect 180064 456758 180116 456764
rect 170496 448588 170548 448594
rect 170496 448530 170548 448536
rect 170508 265470 170536 448530
rect 171784 409896 171836 409902
rect 171784 409838 171836 409844
rect 170496 265464 170548 265470
rect 170496 265406 170548 265412
rect 171796 265402 171824 409838
rect 171876 397520 171928 397526
rect 171876 397462 171928 397468
rect 171784 265396 171836 265402
rect 171784 265338 171836 265344
rect 170404 265328 170456 265334
rect 170404 265270 170456 265276
rect 170680 265328 170732 265334
rect 170680 265270 170732 265276
rect 170692 259978 170720 265270
rect 171692 263288 171744 263294
rect 171692 263230 171744 263236
rect 171704 262750 171732 263230
rect 171692 262744 171744 262750
rect 171692 262686 171744 262692
rect 171002 260160 171054 260166
rect 171002 260102 171054 260108
rect 168760 259950 168820 259978
rect 168944 259950 169372 259978
rect 169924 259950 170260 259978
rect 170476 259950 170720 259978
rect 171014 259964 171042 260102
rect 171704 259978 171732 262686
rect 171580 259950 171732 259978
rect 171796 259978 171824 265338
rect 171888 263294 171916 397462
rect 178684 378208 178736 378214
rect 178684 378150 178736 378156
rect 173900 318844 173952 318850
rect 173900 318786 173952 318792
rect 173164 291848 173216 291854
rect 173164 291790 173216 291796
rect 172704 269884 172756 269890
rect 172704 269826 172756 269832
rect 172716 267734 172744 269826
rect 173176 267734 173204 291790
rect 172716 267706 172836 267734
rect 173176 267706 173480 267734
rect 172808 265606 172836 267706
rect 173348 265804 173400 265810
rect 173348 265746 173400 265752
rect 172796 265600 172848 265606
rect 172796 265542 172848 265548
rect 172612 263900 172664 263906
rect 172612 263842 172664 263848
rect 171876 263288 171928 263294
rect 171876 263230 171928 263236
rect 171796 259950 172132 259978
rect 172624 259842 172652 263842
rect 172808 259978 172836 265542
rect 173360 263906 173388 265746
rect 173452 265538 173480 267706
rect 173440 265532 173492 265538
rect 173440 265474 173492 265480
rect 173348 263900 173400 263906
rect 173348 263842 173400 263848
rect 173452 259978 173480 265474
rect 173912 260438 173940 318786
rect 175924 305040 175976 305046
rect 175924 304982 175976 304988
rect 174544 292596 174596 292602
rect 174544 292538 174596 292544
rect 174556 265674 174584 292538
rect 175936 267734 175964 304982
rect 178696 271250 178724 378150
rect 178684 271244 178736 271250
rect 178684 271186 178736 271192
rect 175752 267706 175964 267734
rect 174544 265668 174596 265674
rect 174544 265610 174596 265616
rect 173900 260432 173952 260438
rect 173900 260374 173952 260380
rect 173912 259978 173940 260374
rect 174556 259978 174584 265610
rect 175752 263838 175780 267706
rect 175924 266416 175976 266422
rect 175924 266358 175976 266364
rect 175740 263832 175792 263838
rect 175740 263774 175792 263780
rect 175752 259978 175780 263774
rect 172808 259950 173236 259978
rect 173452 259950 173788 259978
rect 173912 259950 174340 259978
rect 174556 259950 174892 259978
rect 175444 259950 175780 259978
rect 175936 259978 175964 266358
rect 180076 264246 180104 456758
rect 181456 265742 181484 510614
rect 182836 279478 182864 643078
rect 184204 404388 184256 404394
rect 184204 404330 184256 404336
rect 182824 279472 182876 279478
rect 182824 279414 182876 279420
rect 184216 276690 184244 404330
rect 184204 276684 184256 276690
rect 184204 276626 184256 276632
rect 185596 268394 185624 670686
rect 198004 630692 198056 630698
rect 198004 630634 198056 630640
rect 188344 536852 188396 536858
rect 188344 536794 188396 536800
rect 188356 278050 188384 536794
rect 198016 286346 198044 630634
rect 198004 286340 198056 286346
rect 198004 286282 198056 286288
rect 189080 284980 189132 284986
rect 189080 284922 189132 284928
rect 189092 284374 189120 284922
rect 189080 284368 189132 284374
rect 189080 284310 189132 284316
rect 188344 278044 188396 278050
rect 188344 277986 188396 277992
rect 187700 275324 187752 275330
rect 187700 275266 187752 275272
rect 187712 274718 187740 275266
rect 187700 274712 187752 274718
rect 187700 274654 187752 274660
rect 185584 268388 185636 268394
rect 185584 268330 185636 268336
rect 181444 265736 181496 265742
rect 181444 265678 181496 265684
rect 180064 264240 180116 264246
rect 180064 264182 180116 264188
rect 177764 263220 177816 263226
rect 177764 263162 177816 263168
rect 176752 262608 176804 262614
rect 176752 262550 176804 262556
rect 176764 261390 176792 262550
rect 177776 261458 177804 263162
rect 178040 263152 178092 263158
rect 178040 263094 178092 263100
rect 178052 262478 178080 263094
rect 182916 262608 182968 262614
rect 182916 262550 182968 262556
rect 178408 262540 178460 262546
rect 178408 262482 178460 262488
rect 178040 262472 178092 262478
rect 178040 262414 178092 262420
rect 177764 261452 177816 261458
rect 177764 261394 177816 261400
rect 176752 261384 176804 261390
rect 176752 261326 176804 261332
rect 176200 260228 176252 260234
rect 176200 260170 176252 260176
rect 175936 259950 176148 259978
rect 176120 259894 176148 259950
rect 176108 259888 176160 259894
rect 162638 259814 162748 259842
rect 168116 259826 168268 259842
rect 168104 259820 168268 259826
rect 162582 259791 162638 259800
rect 168156 259814 168268 259820
rect 172624 259814 172684 259842
rect 176108 259830 176160 259836
rect 176212 259842 176240 260170
rect 176764 259978 176792 261326
rect 176764 259950 177100 259978
rect 177776 259842 177804 261394
rect 178052 259978 178080 262414
rect 178420 261050 178448 262482
rect 181260 262268 181312 262274
rect 181260 262210 181312 262216
rect 180156 261248 180208 261254
rect 180156 261190 180208 261196
rect 178408 261044 178460 261050
rect 178408 260986 178460 260992
rect 178420 259978 178448 260986
rect 180168 259978 180196 261190
rect 180524 261180 180576 261186
rect 180524 261122 180576 261128
rect 180536 259978 180564 261122
rect 181272 259978 181300 262210
rect 181996 261112 182048 261118
rect 181996 261054 182048 261060
rect 181812 260976 181864 260982
rect 181812 260918 181864 260924
rect 181824 259978 181852 260918
rect 181904 260432 181956 260438
rect 181904 260374 181956 260380
rect 181916 260098 181944 260374
rect 181904 260092 181956 260098
rect 181904 260034 181956 260040
rect 178052 259950 178204 259978
rect 178420 259950 178756 259978
rect 179860 259950 180196 259978
rect 180412 259950 180564 259978
rect 180964 259950 181300 259978
rect 181516 259950 181852 259978
rect 182008 259978 182036 261054
rect 182928 259978 182956 262550
rect 183468 262336 183520 262342
rect 183468 262278 183520 262284
rect 183480 259978 183508 262278
rect 184756 260908 184808 260914
rect 184756 260850 184808 260856
rect 184112 260228 184164 260234
rect 184112 260170 184164 260176
rect 182008 259950 182068 259978
rect 182620 259950 182956 259978
rect 183172 259950 183508 259978
rect 176212 259814 176548 259842
rect 177652 259814 177804 259842
rect 168104 259762 168156 259768
rect 156786 259655 156842 259664
rect 158628 259684 158680 259690
rect 143080 259626 143132 259632
rect 158628 259626 158680 259632
rect 131394 259584 131450 259593
rect 124916 259564 125212 259570
rect 124864 259558 125212 259564
rect 124876 259542 125212 259558
rect 126532 259542 126868 259570
rect 129292 259554 129628 259570
rect 129280 259548 129628 259554
rect 123758 259519 123814 259528
rect 126532 259486 126560 259542
rect 129332 259542 129628 259548
rect 131394 259519 131450 259528
rect 129280 259490 129332 259496
rect 176396 259486 176424 259814
rect 184124 259690 184152 260170
rect 184768 259978 184796 260850
rect 185674 260264 185730 260273
rect 185674 260199 185730 260208
rect 184768 259950 184828 259978
rect 185688 259729 185716 260199
rect 185674 259720 185730 259729
rect 184276 259690 184612 259706
rect 184112 259684 184164 259690
rect 184276 259684 184624 259690
rect 184276 259678 184572 259684
rect 184112 259626 184164 259632
rect 185674 259655 185730 259664
rect 184572 259626 184624 259632
rect 179420 259616 179472 259622
rect 179308 259564 179420 259570
rect 179308 259558 179472 259564
rect 179308 259542 179460 259558
rect 183724 259554 184060 259570
rect 183724 259548 184072 259554
rect 183724 259542 184020 259548
rect 185380 259542 185716 259570
rect 184020 259490 184072 259496
rect 126520 259480 126572 259486
rect 126520 259422 126572 259428
rect 176384 259480 176436 259486
rect 185688 259457 185716 259542
rect 176384 259422 176436 259428
rect 185674 259448 185730 259457
rect 185674 259383 185730 259392
rect 187148 200864 187200 200870
rect 187148 200806 187200 200812
rect 123944 200728 123996 200734
rect 123944 200670 123996 200676
rect 131856 200728 131908 200734
rect 132040 200728 132092 200734
rect 131856 200670 131908 200676
rect 131946 200696 132002 200705
rect 123956 200530 123984 200670
rect 128726 200560 128782 200569
rect 123944 200524 123996 200530
rect 128726 200495 128782 200504
rect 129004 200524 129056 200530
rect 123944 200466 123996 200472
rect 127622 200152 127678 200161
rect 125048 200116 125100 200122
rect 127622 200087 127678 200096
rect 125048 200058 125100 200064
rect 123576 199436 123628 199442
rect 123576 199378 123628 199384
rect 122102 199064 122158 199073
rect 122102 198999 122158 199008
rect 121368 197260 121420 197266
rect 121368 197202 121420 197208
rect 122116 138825 122144 198999
rect 123588 198898 123616 199378
rect 123576 198892 123628 198898
rect 123576 198834 123628 198840
rect 123576 198484 123628 198490
rect 123576 198426 123628 198432
rect 123484 196920 123536 196926
rect 123484 196862 123536 196868
rect 123496 196518 123524 196862
rect 123484 196512 123536 196518
rect 123484 196454 123536 196460
rect 123588 195974 123616 198426
rect 124864 197328 124916 197334
rect 124864 197270 124916 197276
rect 123496 195946 123616 195974
rect 122288 195900 122340 195906
rect 122288 195842 122340 195848
rect 122194 195664 122250 195673
rect 122194 195599 122250 195608
rect 122208 139466 122236 195599
rect 122196 139460 122248 139466
rect 122196 139402 122248 139408
rect 122102 138816 122158 138825
rect 122102 138751 122158 138760
rect 122300 138553 122328 195842
rect 122378 195800 122434 195809
rect 122378 195735 122434 195744
rect 122392 139777 122420 195735
rect 122472 148844 122524 148850
rect 122472 148786 122524 148792
rect 122484 140865 122512 148786
rect 123496 142154 123524 195946
rect 123944 193044 123996 193050
rect 123944 192986 123996 192992
rect 123574 148880 123630 148889
rect 123574 148815 123630 148824
rect 123404 142126 123524 142154
rect 122470 140856 122526 140865
rect 122470 140791 122526 140800
rect 123404 140554 123432 142126
rect 123392 140548 123444 140554
rect 123392 140490 123444 140496
rect 122378 139768 122434 139777
rect 122378 139703 122434 139712
rect 122746 138816 122802 138825
rect 122746 138751 122802 138760
rect 122286 138544 122342 138553
rect 122286 138479 122342 138488
rect 122760 138009 122788 138751
rect 123588 138417 123616 148815
rect 123666 142080 123722 142089
rect 123666 142015 123722 142024
rect 123680 139890 123708 142015
rect 123680 139862 123832 139890
rect 123956 138825 123984 192986
rect 124036 150952 124088 150958
rect 124036 150894 124088 150900
rect 123942 138816 123998 138825
rect 123942 138751 123998 138760
rect 123574 138408 123630 138417
rect 123574 138343 123630 138352
rect 124048 138145 124076 150894
rect 124220 143540 124272 143546
rect 124220 143482 124272 143488
rect 124232 140865 124260 143482
rect 124876 143478 124904 197270
rect 124956 197192 125008 197198
rect 124956 197134 125008 197140
rect 124968 144226 124996 197134
rect 125060 150482 125088 200058
rect 126612 200048 126664 200054
rect 126612 199990 126664 199996
rect 126336 197192 126388 197198
rect 126336 197134 126388 197140
rect 126244 195968 126296 195974
rect 126244 195910 126296 195916
rect 125048 150476 125100 150482
rect 125048 150418 125100 150424
rect 124956 144220 125008 144226
rect 124956 144162 125008 144168
rect 124864 143472 124916 143478
rect 124864 143414 124916 143420
rect 124862 142624 124918 142633
rect 124862 142559 124918 142568
rect 124876 142225 124904 142559
rect 124862 142216 124918 142225
rect 124862 142151 124918 142160
rect 124218 140856 124274 140865
rect 124218 140791 124274 140800
rect 124678 140856 124734 140865
rect 124678 140791 124734 140800
rect 124692 139890 124720 140791
rect 124384 139862 124720 139890
rect 124876 139890 124904 142151
rect 125060 139890 125088 150418
rect 125692 149116 125744 149122
rect 125692 149058 125744 149064
rect 125508 142112 125560 142118
rect 125560 142060 125640 142066
rect 125508 142054 125640 142060
rect 125520 142038 125640 142054
rect 124876 139862 124936 139890
rect 125060 139862 125488 139890
rect 125612 139482 125640 142038
rect 125704 139942 125732 149058
rect 125692 139936 125744 139942
rect 125692 139878 125744 139884
rect 125612 139466 126192 139482
rect 125612 139460 126204 139466
rect 125612 139454 126152 139460
rect 126152 139402 126204 139408
rect 126256 139369 126284 195910
rect 126348 140593 126376 197134
rect 126520 196580 126572 196586
rect 126520 196522 126572 196528
rect 126426 195528 126482 195537
rect 126426 195463 126482 195472
rect 126334 140584 126390 140593
rect 126334 140519 126390 140528
rect 126440 140010 126468 195463
rect 126532 149122 126560 196522
rect 126624 194177 126652 199990
rect 127164 199844 127216 199850
rect 127164 199786 127216 199792
rect 126980 199776 127032 199782
rect 126980 199718 127032 199724
rect 126610 194168 126666 194177
rect 126992 194138 127020 199718
rect 127176 198257 127204 199786
rect 127162 198248 127218 198257
rect 127162 198183 127218 198192
rect 126610 194103 126666 194112
rect 126980 194132 127032 194138
rect 126980 194074 127032 194080
rect 126520 149116 126572 149122
rect 126520 149058 126572 149064
rect 127440 143404 127492 143410
rect 127440 143346 127492 143352
rect 127452 141137 127480 143346
rect 127532 142044 127584 142050
rect 127532 141986 127584 141992
rect 127438 141128 127494 141137
rect 127438 141063 127494 141072
rect 126428 140004 126480 140010
rect 126428 139946 126480 139952
rect 126336 139936 126388 139942
rect 127452 139890 127480 141063
rect 127544 141001 127572 141986
rect 127530 140992 127586 141001
rect 127530 140927 127586 140936
rect 126388 139884 126592 139890
rect 126336 139878 126592 139884
rect 126348 139862 126592 139878
rect 127144 139862 127480 139890
rect 127544 139890 127572 140927
rect 127636 140321 127664 200087
rect 128740 199889 128768 200495
rect 129004 200466 129056 200472
rect 128726 199880 128782 199889
rect 128726 199815 128782 199824
rect 127900 199436 127952 199442
rect 127900 199378 127952 199384
rect 127716 197328 127768 197334
rect 127716 197270 127768 197276
rect 127728 140690 127756 197270
rect 127808 196444 127860 196450
rect 127808 196386 127860 196392
rect 127716 140684 127768 140690
rect 127716 140626 127768 140632
rect 127820 140622 127848 196386
rect 127912 144158 127940 199378
rect 127992 197260 128044 197266
rect 127992 197202 128044 197208
rect 128084 197260 128136 197266
rect 128084 197202 128136 197208
rect 127900 144152 127952 144158
rect 127900 144094 127952 144100
rect 128004 142186 128032 197202
rect 128096 197130 128124 197202
rect 128084 197124 128136 197130
rect 128084 197066 128136 197072
rect 128176 197124 128228 197130
rect 128176 197066 128228 197072
rect 128188 196382 128216 197066
rect 128176 196376 128228 196382
rect 128176 196318 128228 196324
rect 128084 196308 128136 196314
rect 128084 196250 128136 196256
rect 128096 142322 128124 196250
rect 128912 148368 128964 148374
rect 128912 148310 128964 148316
rect 128728 143336 128780 143342
rect 128728 143278 128780 143284
rect 128740 142526 128768 143278
rect 128728 142520 128780 142526
rect 128728 142462 128780 142468
rect 128084 142316 128136 142322
rect 128084 142258 128136 142264
rect 127992 142180 128044 142186
rect 127992 142122 128044 142128
rect 127808 140616 127860 140622
rect 127808 140558 127860 140564
rect 127622 140312 127678 140321
rect 127622 140247 127678 140256
rect 128096 139890 128124 142258
rect 128740 139890 128768 142462
rect 128924 139890 128952 148310
rect 129016 140418 129044 200466
rect 131868 200394 131896 200670
rect 132040 200670 132092 200676
rect 180064 200728 180116 200734
rect 180064 200670 180116 200676
rect 180524 200728 180576 200734
rect 180524 200670 180576 200676
rect 131946 200631 132002 200640
rect 131856 200388 131908 200394
rect 131856 200330 131908 200336
rect 129648 200184 129700 200190
rect 129648 200126 129700 200132
rect 129280 199912 129332 199918
rect 129280 199854 129332 199860
rect 129186 198792 129242 198801
rect 129186 198727 129242 198736
rect 129096 196580 129148 196586
rect 129096 196522 129148 196528
rect 129108 140486 129136 196522
rect 129200 144294 129228 198727
rect 129292 198121 129320 199854
rect 129278 198112 129334 198121
rect 129278 198047 129334 198056
rect 129660 195401 129688 200126
rect 130660 199980 130712 199986
rect 130660 199922 130712 199928
rect 129740 196512 129792 196518
rect 129740 196454 129792 196460
rect 129646 195392 129702 195401
rect 129646 195327 129702 195336
rect 129280 195220 129332 195226
rect 129280 195162 129332 195168
rect 129188 144288 129240 144294
rect 129188 144230 129240 144236
rect 129292 143274 129320 195162
rect 129752 193089 129780 196454
rect 130384 194404 130436 194410
rect 130384 194346 130436 194352
rect 129738 193080 129794 193089
rect 129738 193015 129794 193024
rect 129372 192432 129424 192438
rect 129372 192374 129424 192380
rect 129280 143268 129332 143274
rect 129280 143210 129332 143216
rect 129384 141370 129412 192374
rect 129740 146260 129792 146266
rect 129740 146202 129792 146208
rect 129372 141364 129424 141370
rect 129372 141306 129424 141312
rect 129752 140758 129780 146202
rect 130016 146192 130068 146198
rect 130016 146134 130068 146140
rect 129924 142452 129976 142458
rect 129924 142394 129976 142400
rect 129832 142180 129884 142186
rect 129936 142168 129964 142394
rect 130028 142186 130056 146134
rect 130108 145512 130160 145518
rect 130108 145454 130160 145460
rect 130120 142254 130148 145454
rect 130292 144288 130344 144294
rect 130292 144230 130344 144236
rect 130304 144090 130332 144230
rect 130292 144084 130344 144090
rect 130292 144026 130344 144032
rect 130108 142248 130160 142254
rect 130108 142190 130160 142196
rect 129884 142140 129964 142168
rect 130016 142180 130068 142186
rect 129832 142122 129884 142128
rect 130016 142122 130068 142128
rect 129740 140752 129792 140758
rect 129740 140694 129792 140700
rect 129096 140480 129148 140486
rect 129096 140422 129148 140428
rect 129004 140412 129056 140418
rect 129004 140354 129056 140360
rect 129844 139890 129872 142122
rect 130304 139890 130332 144026
rect 130396 140350 130424 194346
rect 130566 193216 130622 193225
rect 130566 193151 130622 193160
rect 130476 192364 130528 192370
rect 130476 192306 130528 192312
rect 130488 141982 130516 192306
rect 130476 141976 130528 141982
rect 130476 141918 130528 141924
rect 130580 140978 130608 193151
rect 130672 148714 130700 199922
rect 131854 199336 131910 199345
rect 131854 199271 131910 199280
rect 131764 196104 131816 196110
rect 131764 196046 131816 196052
rect 130752 192296 130804 192302
rect 130752 192238 130804 192244
rect 130660 148708 130712 148714
rect 130660 148650 130712 148656
rect 130488 140950 130608 140978
rect 130384 140344 130436 140350
rect 130488 140321 130516 140950
rect 130764 140842 130792 192238
rect 131776 151814 131804 196046
rect 131684 151786 131804 151814
rect 131488 144220 131540 144226
rect 131488 144162 131540 144168
rect 130580 140814 130792 140842
rect 130384 140286 130436 140292
rect 130474 140312 130530 140321
rect 130474 140247 130530 140256
rect 127544 139862 127696 139890
rect 128096 139862 128248 139890
rect 128740 139862 128800 139890
rect 128924 139862 129352 139890
rect 129844 139862 129904 139890
rect 130304 139862 130456 139890
rect 130580 139369 130608 140814
rect 130660 140752 130712 140758
rect 130660 140694 130712 140700
rect 130672 139890 130700 140694
rect 131500 139890 131528 144162
rect 131684 140049 131712 151786
rect 131868 148238 131896 199271
rect 131960 148986 131988 200631
rect 132052 200530 132080 200670
rect 132224 200592 132276 200598
rect 132222 200560 132224 200569
rect 132276 200560 132278 200569
rect 132040 200524 132092 200530
rect 132222 200495 132278 200504
rect 132040 200466 132092 200472
rect 177946 200424 178002 200433
rect 177856 200388 177908 200394
rect 177946 200359 178002 200368
rect 177856 200330 177908 200336
rect 132052 200110 132388 200138
rect 132052 193905 132080 200110
rect 132466 199866 132494 200124
rect 132420 199838 132494 199866
rect 132558 199850 132586 200124
rect 132546 199844 132598 199850
rect 132316 199708 132368 199714
rect 132316 199650 132368 199656
rect 132222 198928 132278 198937
rect 132222 198863 132278 198872
rect 132132 198620 132184 198626
rect 132132 198562 132184 198568
rect 132144 198218 132172 198562
rect 132132 198212 132184 198218
rect 132132 198154 132184 198160
rect 132236 196058 132264 198863
rect 132144 196030 132264 196058
rect 132038 193896 132094 193905
rect 132038 193831 132094 193840
rect 132144 190738 132172 196030
rect 132224 194744 132276 194750
rect 132224 194686 132276 194692
rect 132132 190732 132184 190738
rect 132132 190674 132184 190680
rect 132132 190528 132184 190534
rect 132132 190470 132184 190476
rect 132040 190392 132092 190398
rect 132040 190334 132092 190340
rect 131948 148980 132000 148986
rect 131948 148922 132000 148928
rect 131856 148232 131908 148238
rect 131856 148174 131908 148180
rect 131854 146296 131910 146305
rect 131854 146231 131910 146240
rect 131868 143206 131896 146231
rect 132052 144770 132080 190334
rect 132144 148753 132172 190470
rect 132236 190398 132264 194686
rect 132328 190398 132356 199650
rect 132420 198393 132448 199838
rect 132546 199786 132598 199792
rect 132650 199730 132678 200124
rect 132604 199702 132678 199730
rect 132406 198384 132462 198393
rect 132406 198319 132462 198328
rect 132604 196518 132632 199702
rect 132742 199458 132770 200124
rect 132834 199730 132862 200124
rect 132926 199918 132954 200124
rect 133018 199918 133046 200124
rect 133110 199918 133138 200124
rect 132914 199912 132966 199918
rect 132914 199854 132966 199860
rect 133006 199912 133058 199918
rect 133006 199854 133058 199860
rect 133098 199912 133150 199918
rect 133098 199854 133150 199860
rect 133202 199764 133230 200124
rect 133294 199889 133322 200124
rect 133280 199880 133336 199889
rect 133280 199815 133336 199824
rect 133202 199736 133276 199764
rect 132834 199702 132908 199730
rect 132742 199430 132816 199458
rect 132592 196512 132644 196518
rect 132592 196454 132644 196460
rect 132408 195084 132460 195090
rect 132408 195026 132460 195032
rect 132224 190392 132276 190398
rect 132224 190334 132276 190340
rect 132316 190392 132368 190398
rect 132316 190334 132368 190340
rect 132420 188426 132448 195026
rect 132788 191350 132816 199430
rect 132776 191344 132828 191350
rect 132776 191286 132828 191292
rect 132500 190392 132552 190398
rect 132500 190334 132552 190340
rect 132224 188420 132276 188426
rect 132224 188362 132276 188368
rect 132408 188420 132460 188426
rect 132408 188362 132460 188368
rect 132130 148744 132186 148753
rect 132130 148679 132186 148688
rect 132236 146130 132264 188362
rect 132512 183554 132540 190334
rect 132880 187241 132908 199702
rect 133052 197464 133104 197470
rect 133052 197406 133104 197412
rect 132960 196988 133012 196994
rect 132960 196930 133012 196936
rect 132972 196246 133000 196930
rect 132960 196240 133012 196246
rect 132960 196182 133012 196188
rect 133064 195838 133092 197406
rect 133144 196784 133196 196790
rect 133144 196726 133196 196732
rect 133156 196314 133184 196726
rect 133144 196308 133196 196314
rect 133144 196250 133196 196256
rect 133052 195832 133104 195838
rect 133052 195774 133104 195780
rect 133144 195560 133196 195566
rect 133144 195502 133196 195508
rect 133156 194818 133184 195502
rect 133144 194812 133196 194818
rect 133144 194754 133196 194760
rect 133052 191072 133104 191078
rect 133052 191014 133104 191020
rect 132866 187232 132922 187241
rect 132866 187167 132922 187176
rect 132328 183526 132540 183554
rect 132328 148578 132356 183526
rect 133064 151570 133092 191014
rect 133248 187134 133276 199736
rect 133386 199628 133414 200124
rect 133340 199600 133414 199628
rect 133478 199628 133506 200124
rect 133570 199730 133598 200124
rect 133662 199889 133690 200124
rect 133754 199918 133782 200124
rect 133742 199912 133794 199918
rect 133648 199880 133704 199889
rect 133846 199889 133874 200124
rect 133938 199918 133966 200124
rect 134030 199923 134058 200124
rect 133926 199912 133978 199918
rect 133742 199854 133794 199860
rect 133832 199880 133888 199889
rect 133648 199815 133704 199824
rect 133926 199854 133978 199860
rect 134016 199914 134072 199923
rect 134122 199918 134150 200124
rect 134016 199849 134072 199858
rect 134110 199912 134162 199918
rect 134110 199854 134162 199860
rect 133832 199815 133888 199824
rect 133696 199776 133748 199782
rect 133570 199702 133644 199730
rect 133972 199776 134024 199782
rect 133696 199718 133748 199724
rect 133786 199744 133842 199753
rect 133478 199600 133552 199628
rect 133340 191185 133368 199600
rect 133524 195956 133552 199600
rect 133432 195928 133552 195956
rect 133326 191176 133382 191185
rect 133326 191111 133382 191120
rect 133236 187128 133288 187134
rect 133236 187070 133288 187076
rect 133432 180794 133460 195928
rect 133616 191834 133644 199702
rect 133524 191806 133644 191834
rect 133524 187202 133552 191806
rect 133708 191457 133736 199718
rect 133972 199718 134024 199724
rect 134064 199776 134116 199782
rect 134214 199730 134242 200124
rect 134306 199782 134334 200124
rect 134398 199918 134426 200124
rect 134490 199918 134518 200124
rect 134386 199912 134438 199918
rect 134386 199854 134438 199860
rect 134478 199912 134530 199918
rect 134582 199889 134610 200124
rect 134674 199918 134702 200124
rect 134662 199912 134714 199918
rect 134478 199854 134530 199860
rect 134568 199880 134624 199889
rect 134766 199889 134794 200124
rect 134858 199918 134886 200124
rect 134846 199912 134898 199918
rect 134662 199854 134714 199860
rect 134752 199880 134808 199889
rect 134568 199815 134624 199824
rect 134846 199854 134898 199860
rect 134752 199815 134808 199824
rect 134064 199718 134116 199724
rect 133786 199679 133842 199688
rect 133694 191448 133750 191457
rect 133694 191383 133750 191392
rect 133800 191078 133828 199679
rect 133878 199472 133934 199481
rect 133878 199407 133934 199416
rect 133892 192953 133920 199407
rect 133878 192944 133934 192953
rect 133878 192879 133934 192888
rect 133788 191072 133840 191078
rect 133788 191014 133840 191020
rect 133984 187474 134012 199718
rect 134076 193214 134104 199718
rect 134168 199702 134242 199730
rect 134294 199776 134346 199782
rect 134386 199776 134438 199782
rect 134294 199718 134346 199724
rect 134384 199744 134386 199753
rect 134616 199776 134668 199782
rect 134438 199744 134440 199753
rect 134168 196489 134196 199702
rect 134384 199679 134440 199688
rect 134522 199744 134578 199753
rect 134616 199718 134668 199724
rect 134708 199776 134760 199782
rect 134950 199764 134978 200124
rect 134904 199753 134978 199764
rect 134708 199718 134760 199724
rect 134890 199744 134978 199753
rect 134522 199679 134578 199688
rect 134154 196480 134210 196489
rect 134154 196415 134210 196424
rect 134536 193214 134564 199679
rect 134628 195265 134656 199718
rect 134614 195256 134670 195265
rect 134614 195191 134670 195200
rect 134076 193186 134288 193214
rect 134260 191834 134288 193186
rect 134444 193186 134564 193214
rect 134720 193214 134748 199718
rect 134946 199736 134978 199744
rect 135042 199714 135070 200124
rect 135134 199923 135162 200124
rect 135120 199914 135176 199923
rect 135120 199849 135176 199858
rect 135226 199764 135254 200124
rect 135318 199918 135346 200124
rect 135410 199918 135438 200124
rect 135502 199923 135530 200124
rect 135306 199912 135358 199918
rect 135306 199854 135358 199860
rect 135398 199912 135450 199918
rect 135398 199854 135450 199860
rect 135488 199914 135544 199923
rect 135594 199918 135622 200124
rect 135686 199918 135714 200124
rect 135778 199923 135806 200124
rect 135488 199849 135544 199858
rect 135582 199912 135634 199918
rect 135582 199854 135634 199860
rect 135674 199912 135726 199918
rect 135674 199854 135726 199860
rect 135764 199914 135820 199923
rect 135764 199849 135820 199858
rect 135870 199764 135898 200124
rect 135962 199918 135990 200124
rect 136054 199918 136082 200124
rect 136146 199918 136174 200124
rect 135950 199912 136002 199918
rect 135950 199854 136002 199860
rect 136042 199912 136094 199918
rect 136042 199854 136094 199860
rect 136134 199912 136186 199918
rect 136134 199854 136186 199860
rect 135996 199776 136048 199782
rect 135226 199736 135300 199764
rect 135870 199736 135944 199764
rect 134890 199679 134946 199688
rect 135030 199708 135082 199714
rect 135030 199650 135082 199656
rect 135272 199628 135300 199736
rect 135720 199708 135772 199714
rect 135720 199650 135772 199656
rect 135444 199640 135496 199646
rect 135074 199608 135130 199617
rect 135272 199600 135346 199628
rect 135074 199543 135130 199552
rect 134982 199472 135038 199481
rect 134982 199407 135038 199416
rect 134892 197396 134944 197402
rect 134892 197338 134944 197344
rect 134720 193186 134840 193214
rect 134260 191806 134380 191834
rect 133972 187468 134024 187474
rect 133972 187410 134024 187416
rect 134352 187338 134380 191806
rect 134340 187332 134392 187338
rect 134340 187274 134392 187280
rect 134444 187218 134472 193186
rect 133512 187196 133564 187202
rect 133512 187138 133564 187144
rect 134076 187190 134472 187218
rect 133156 180766 133460 180794
rect 133052 151564 133104 151570
rect 133052 151506 133104 151512
rect 133156 151230 133184 180766
rect 133972 154216 134024 154222
rect 133972 154158 134024 154164
rect 133144 151224 133196 151230
rect 133144 151166 133196 151172
rect 132316 148572 132368 148578
rect 132316 148514 132368 148520
rect 132224 146124 132276 146130
rect 132224 146066 132276 146072
rect 132040 144764 132092 144770
rect 132040 144706 132092 144712
rect 132868 143472 132920 143478
rect 132868 143414 132920 143420
rect 131764 143200 131816 143206
rect 131764 143142 131816 143148
rect 131856 143200 131908 143206
rect 131856 143142 131908 143148
rect 131670 140040 131726 140049
rect 131670 139975 131726 139984
rect 131776 139890 131804 143142
rect 132500 142180 132552 142186
rect 132500 142122 132552 142128
rect 132512 139890 132540 142122
rect 132880 139890 132908 143414
rect 133420 143132 133472 143138
rect 133420 143074 133472 143080
rect 133432 139890 133460 143074
rect 133512 142452 133564 142458
rect 133512 142394 133564 142400
rect 133524 142254 133552 142394
rect 133512 142248 133564 142254
rect 133512 142190 133564 142196
rect 133984 139890 134012 154158
rect 134076 151366 134104 187190
rect 134248 186516 134300 186522
rect 134248 186458 134300 186464
rect 134260 151706 134288 186458
rect 134812 186314 134840 193186
rect 134352 186286 134840 186314
rect 134248 151700 134300 151706
rect 134248 151642 134300 151648
rect 134352 151434 134380 186286
rect 134904 180794 134932 197338
rect 134996 192846 135024 199407
rect 134984 192840 135036 192846
rect 134984 192782 135036 192788
rect 135088 186522 135116 199543
rect 135318 199492 135346 199600
rect 135628 199640 135680 199646
rect 135496 199588 135576 199594
rect 135444 199582 135576 199588
rect 135628 199582 135680 199588
rect 135456 199566 135576 199582
rect 135272 199464 135346 199492
rect 135272 199458 135300 199464
rect 135180 199430 135300 199458
rect 135180 192914 135208 199430
rect 135548 197146 135576 199566
rect 135456 197118 135576 197146
rect 135456 196897 135484 197118
rect 135534 197024 135590 197033
rect 135534 196959 135590 196968
rect 135442 196888 135498 196897
rect 135442 196823 135498 196832
rect 135444 196784 135496 196790
rect 135444 196726 135496 196732
rect 135168 192908 135220 192914
rect 135168 192850 135220 192856
rect 135076 186516 135128 186522
rect 135076 186458 135128 186464
rect 135456 186314 135484 196726
rect 135548 194070 135576 196959
rect 135536 194064 135588 194070
rect 135536 194006 135588 194012
rect 135640 187542 135668 199582
rect 135732 191078 135760 199650
rect 135812 199640 135864 199646
rect 135812 199582 135864 199588
rect 135824 196790 135852 199582
rect 135812 196784 135864 196790
rect 135812 196726 135864 196732
rect 135916 196081 135944 199736
rect 136238 199764 136266 200124
rect 136330 199918 136358 200124
rect 136422 199923 136450 200124
rect 136318 199912 136370 199918
rect 136318 199854 136370 199860
rect 136408 199914 136464 199923
rect 136514 199918 136542 200124
rect 136408 199849 136464 199858
rect 136502 199912 136554 199918
rect 136502 199854 136554 199860
rect 135996 199718 136048 199724
rect 136192 199736 136266 199764
rect 136364 199776 136416 199782
rect 136008 198626 136036 199718
rect 136088 199708 136140 199714
rect 136088 199650 136140 199656
rect 135996 198620 136048 198626
rect 135996 198562 136048 198568
rect 135996 197532 136048 197538
rect 135996 197474 136048 197480
rect 135902 196072 135958 196081
rect 135902 196007 135958 196016
rect 135904 195832 135956 195838
rect 135904 195774 135956 195780
rect 135812 195764 135864 195770
rect 135812 195706 135864 195712
rect 135824 195566 135852 195706
rect 135812 195560 135864 195566
rect 135812 195502 135864 195508
rect 135720 191072 135772 191078
rect 135720 191014 135772 191020
rect 135720 187740 135772 187746
rect 135720 187682 135772 187688
rect 135628 187536 135680 187542
rect 135628 187478 135680 187484
rect 135456 186286 135576 186314
rect 134536 180766 134932 180794
rect 134536 154154 134564 180766
rect 134524 154148 134576 154154
rect 134524 154090 134576 154096
rect 134340 151428 134392 151434
rect 134340 151370 134392 151376
rect 134064 151360 134116 151366
rect 134064 151302 134116 151308
rect 135548 151162 135576 186286
rect 135536 151156 135588 151162
rect 135536 151098 135588 151104
rect 135732 147150 135760 187682
rect 135916 186314 135944 195774
rect 136008 193866 136036 197474
rect 135996 193860 136048 193866
rect 135996 193802 136048 193808
rect 136100 191834 136128 199650
rect 136192 195945 136220 199736
rect 136364 199718 136416 199724
rect 136454 199744 136510 199753
rect 136376 196761 136404 199718
rect 136606 199730 136634 200124
rect 136698 199918 136726 200124
rect 136790 199923 136818 200124
rect 136686 199912 136738 199918
rect 136686 199854 136738 199860
rect 136776 199914 136832 199923
rect 136776 199849 136832 199858
rect 136732 199776 136784 199782
rect 136510 199702 136634 199730
rect 136730 199744 136732 199753
rect 136784 199744 136786 199753
rect 136882 199730 136910 200124
rect 136454 199679 136510 199688
rect 136730 199679 136786 199688
rect 136836 199702 136910 199730
rect 136974 199730 137002 200124
rect 137066 199918 137094 200124
rect 137054 199912 137106 199918
rect 137054 199854 137106 199860
rect 137158 199850 137186 200124
rect 137146 199844 137198 199850
rect 137146 199786 137198 199792
rect 136974 199702 137048 199730
rect 136548 199640 136600 199646
rect 136732 199640 136784 199646
rect 136548 199582 136600 199588
rect 136638 199608 136694 199617
rect 136454 198384 136510 198393
rect 136454 198319 136510 198328
rect 136362 196752 136418 196761
rect 136362 196687 136418 196696
rect 136178 195936 136234 195945
rect 136178 195871 136234 195880
rect 136468 191834 136496 198319
rect 136008 191806 136128 191834
rect 136376 191806 136496 191834
rect 136008 189990 136036 191806
rect 136088 191072 136140 191078
rect 136088 191014 136140 191020
rect 135996 189984 136048 189990
rect 135996 189926 136048 189932
rect 135824 186286 135944 186314
rect 135824 151638 135852 186286
rect 135812 151632 135864 151638
rect 135812 151574 135864 151580
rect 136100 151298 136128 191014
rect 136376 190194 136404 191806
rect 136364 190188 136416 190194
rect 136364 190130 136416 190136
rect 136560 187746 136588 199582
rect 136732 199582 136784 199588
rect 136638 199543 136694 199552
rect 136652 191834 136680 199543
rect 136744 195838 136772 199582
rect 136836 198937 136864 199702
rect 136916 199640 136968 199646
rect 136916 199582 136968 199588
rect 136822 198928 136878 198937
rect 136822 198863 136878 198872
rect 136824 198620 136876 198626
rect 136824 198562 136876 198568
rect 136836 196654 136864 198562
rect 136928 198082 136956 199582
rect 136916 198076 136968 198082
rect 136916 198018 136968 198024
rect 136824 196648 136876 196654
rect 136824 196590 136876 196596
rect 136732 195832 136784 195838
rect 136732 195774 136784 195780
rect 136652 191806 136864 191834
rect 136836 190233 136864 191806
rect 137020 190369 137048 199702
rect 137100 199708 137152 199714
rect 137100 199650 137152 199656
rect 137006 190360 137062 190369
rect 137006 190295 137062 190304
rect 136822 190224 136878 190233
rect 136822 190159 136878 190168
rect 137112 190074 137140 199650
rect 137250 199628 137278 200124
rect 137342 199918 137370 200124
rect 137434 199923 137462 200124
rect 137330 199912 137382 199918
rect 137330 199854 137382 199860
rect 137420 199914 137476 199923
rect 137420 199849 137476 199858
rect 137376 199776 137428 199782
rect 137526 199764 137554 200124
rect 137376 199718 137428 199724
rect 137480 199736 137554 199764
rect 137204 199600 137278 199628
rect 137204 190262 137232 199600
rect 137388 196761 137416 199718
rect 137374 196752 137430 196761
rect 137374 196687 137430 196696
rect 137376 196648 137428 196654
rect 137376 196590 137428 196596
rect 137192 190256 137244 190262
rect 137192 190198 137244 190204
rect 137388 190210 137416 196590
rect 137480 191282 137508 199736
rect 137618 199696 137646 200124
rect 137710 199923 137738 200124
rect 137696 199914 137752 199923
rect 137696 199849 137752 199858
rect 137802 199764 137830 200124
rect 137894 199918 137922 200124
rect 137986 199918 138014 200124
rect 137882 199912 137934 199918
rect 137882 199854 137934 199860
rect 137974 199912 138026 199918
rect 137974 199854 138026 199860
rect 138078 199764 138106 200124
rect 137572 199668 137646 199696
rect 137756 199736 137830 199764
rect 138032 199736 138106 199764
rect 138170 199764 138198 200124
rect 138262 199918 138290 200124
rect 138354 199918 138382 200124
rect 138250 199912 138302 199918
rect 138250 199854 138302 199860
rect 138342 199912 138394 199918
rect 138342 199854 138394 199860
rect 138170 199736 138244 199764
rect 137468 191276 137520 191282
rect 137468 191218 137520 191224
rect 137388 190182 137508 190210
rect 137112 190046 137416 190074
rect 137284 189984 137336 189990
rect 137284 189926 137336 189932
rect 137192 188692 137244 188698
rect 137192 188634 137244 188640
rect 136548 187740 136600 187746
rect 136548 187682 136600 187688
rect 136088 151292 136140 151298
rect 136088 151234 136140 151240
rect 137204 147286 137232 188634
rect 137192 147280 137244 147286
rect 137192 147222 137244 147228
rect 135720 147144 135772 147150
rect 135720 147086 135772 147092
rect 137296 147082 137324 189926
rect 137388 151502 137416 190046
rect 137480 189990 137508 190182
rect 137468 189984 137520 189990
rect 137468 189926 137520 189932
rect 137572 188698 137600 199668
rect 137650 199608 137706 199617
rect 137650 199543 137706 199552
rect 137664 197062 137692 199543
rect 137652 197056 137704 197062
rect 137652 196998 137704 197004
rect 137756 193214 137784 199736
rect 137928 199708 137980 199714
rect 137928 199650 137980 199656
rect 137836 199640 137888 199646
rect 137836 199582 137888 199588
rect 137848 196654 137876 199582
rect 137940 197470 137968 199650
rect 138032 198937 138060 199736
rect 138112 199640 138164 199646
rect 138110 199608 138112 199617
rect 138164 199608 138166 199617
rect 138110 199543 138166 199552
rect 138018 198928 138074 198937
rect 138018 198863 138074 198872
rect 137928 197464 137980 197470
rect 137928 197406 137980 197412
rect 138216 197402 138244 199736
rect 138446 199696 138474 200124
rect 138538 199918 138566 200124
rect 138630 199923 138658 200124
rect 138526 199912 138578 199918
rect 138526 199854 138578 199860
rect 138616 199914 138672 199923
rect 138616 199849 138672 199858
rect 138572 199776 138624 199782
rect 138722 199764 138750 200124
rect 138814 199918 138842 200124
rect 138802 199912 138854 199918
rect 138802 199854 138854 199860
rect 138676 199753 138750 199764
rect 138572 199718 138624 199724
rect 138662 199744 138750 199753
rect 138400 199668 138474 199696
rect 138296 199640 138348 199646
rect 138296 199582 138348 199588
rect 138204 197396 138256 197402
rect 138204 197338 138256 197344
rect 137836 196648 137888 196654
rect 137836 196590 137888 196596
rect 138020 195764 138072 195770
rect 138020 195706 138072 195712
rect 138032 195566 138060 195706
rect 138020 195560 138072 195566
rect 138020 195502 138072 195508
rect 137664 193186 137784 193214
rect 137664 191554 137692 193186
rect 137652 191548 137704 191554
rect 137652 191490 137704 191496
rect 137560 188692 137612 188698
rect 137560 188634 137612 188640
rect 138308 187270 138336 199582
rect 138400 193214 138428 199668
rect 138478 198656 138534 198665
rect 138478 198591 138534 198600
rect 138492 194750 138520 198591
rect 138584 198393 138612 199718
rect 138718 199736 138750 199744
rect 138906 199764 138934 200124
rect 138998 199923 139026 200124
rect 138984 199914 139040 199923
rect 138984 199849 139040 199858
rect 138906 199736 138980 199764
rect 138662 199679 138718 199688
rect 138664 199640 138716 199646
rect 138664 199582 138716 199588
rect 138756 199640 138808 199646
rect 138756 199582 138808 199588
rect 138676 198626 138704 199582
rect 138664 198620 138716 198626
rect 138664 198562 138716 198568
rect 138570 198384 138626 198393
rect 138570 198319 138626 198328
rect 138572 198280 138624 198286
rect 138572 198222 138624 198228
rect 138584 197810 138612 198222
rect 138572 197804 138624 197810
rect 138572 197746 138624 197752
rect 138480 194744 138532 194750
rect 138480 194686 138532 194692
rect 138400 193186 138612 193214
rect 138388 191140 138440 191146
rect 138388 191082 138440 191088
rect 138296 187264 138348 187270
rect 138296 187206 138348 187212
rect 137376 151496 137428 151502
rect 137376 151438 137428 151444
rect 137284 147076 137336 147082
rect 137284 147018 137336 147024
rect 135352 144900 135404 144906
rect 135352 144842 135404 144848
rect 134524 142180 134576 142186
rect 134524 142122 134576 142128
rect 134536 139890 134564 142122
rect 135364 139890 135392 144842
rect 136180 144832 136232 144838
rect 136180 144774 136232 144780
rect 135628 141908 135680 141914
rect 135628 141850 135680 141856
rect 135640 139890 135668 141850
rect 136192 139890 136220 144774
rect 138020 144696 138072 144702
rect 138020 144638 138072 144644
rect 137284 144628 137336 144634
rect 137284 144570 137336 144576
rect 137008 142520 137060 142526
rect 137008 142462 137060 142468
rect 137020 142186 137048 142462
rect 137008 142180 137060 142186
rect 137008 142122 137060 142128
rect 136730 141400 136786 141409
rect 136730 141335 136786 141344
rect 136744 139890 136772 141335
rect 137296 139890 137324 144570
rect 138032 139890 138060 144638
rect 138400 142154 138428 191082
rect 138584 147354 138612 193186
rect 138768 191834 138796 199582
rect 138846 198928 138902 198937
rect 138846 198863 138902 198872
rect 138860 196314 138888 198863
rect 138848 196308 138900 196314
rect 138848 196250 138900 196256
rect 138952 196110 138980 199736
rect 139090 199730 139118 200124
rect 139182 199923 139210 200124
rect 139168 199914 139224 199923
rect 139274 199918 139302 200124
rect 139366 199918 139394 200124
rect 139458 199918 139486 200124
rect 139550 199918 139578 200124
rect 139168 199849 139224 199858
rect 139262 199912 139314 199918
rect 139262 199854 139314 199860
rect 139354 199912 139406 199918
rect 139354 199854 139406 199860
rect 139446 199912 139498 199918
rect 139446 199854 139498 199860
rect 139538 199912 139590 199918
rect 139538 199854 139590 199860
rect 139216 199776 139268 199782
rect 139090 199702 139164 199730
rect 139492 199776 139544 199782
rect 139216 199718 139268 199724
rect 139398 199744 139454 199753
rect 139030 199608 139086 199617
rect 139030 199543 139086 199552
rect 138940 196104 138992 196110
rect 138940 196046 138992 196052
rect 138676 191806 138796 191834
rect 138676 147665 138704 191806
rect 139044 186314 139072 199543
rect 139136 194818 139164 199702
rect 139124 194812 139176 194818
rect 139124 194754 139176 194760
rect 139228 191146 139256 199718
rect 139308 199708 139360 199714
rect 139642 199764 139670 200124
rect 139734 199918 139762 200124
rect 139826 199923 139854 200124
rect 139722 199912 139774 199918
rect 139722 199854 139774 199860
rect 139812 199914 139868 199923
rect 139918 199918 139946 200124
rect 140010 199918 140038 200124
rect 139812 199849 139868 199858
rect 139906 199912 139958 199918
rect 139906 199854 139958 199860
rect 139998 199912 140050 199918
rect 139998 199854 140050 199860
rect 139768 199776 139820 199782
rect 139642 199736 139716 199764
rect 139492 199718 139544 199724
rect 139398 199679 139400 199688
rect 139308 199650 139360 199656
rect 139452 199679 139454 199688
rect 139400 199650 139452 199656
rect 139320 193934 139348 199650
rect 139398 199608 139454 199617
rect 139398 199543 139454 199552
rect 139412 198490 139440 199543
rect 139400 198484 139452 198490
rect 139400 198426 139452 198432
rect 139400 196784 139452 196790
rect 139400 196726 139452 196732
rect 139308 193928 139360 193934
rect 139308 193870 139360 193876
rect 139412 191593 139440 196726
rect 139398 191584 139454 191593
rect 139398 191519 139454 191528
rect 139504 191486 139532 199718
rect 139582 199472 139638 199481
rect 139582 199407 139638 199416
rect 139492 191480 139544 191486
rect 139492 191422 139544 191428
rect 139216 191140 139268 191146
rect 139216 191082 139268 191088
rect 139596 186314 139624 199407
rect 139688 196761 139716 199736
rect 139768 199718 139820 199724
rect 139860 199776 139912 199782
rect 139860 199718 139912 199724
rect 139952 199776 140004 199782
rect 140102 199764 140130 200124
rect 140194 199923 140222 200124
rect 140180 199914 140236 199923
rect 140286 199918 140314 200124
rect 140180 199849 140236 199858
rect 140274 199912 140326 199918
rect 140274 199854 140326 199860
rect 140378 199850 140406 200124
rect 140470 199923 140498 200124
rect 140456 199914 140512 199923
rect 140366 199844 140418 199850
rect 140456 199849 140512 199858
rect 140366 199786 140418 199792
rect 140102 199736 140176 199764
rect 139952 199718 140004 199724
rect 139780 196790 139808 199718
rect 139768 196784 139820 196790
rect 139674 196752 139730 196761
rect 139768 196726 139820 196732
rect 139872 196722 139900 199718
rect 139674 196687 139730 196696
rect 139860 196716 139912 196722
rect 139860 196658 139912 196664
rect 139964 187406 139992 199718
rect 140042 197024 140098 197033
rect 140042 196959 140098 196968
rect 140056 196450 140084 196959
rect 140044 196444 140096 196450
rect 140044 196386 140096 196392
rect 140148 191834 140176 199736
rect 140226 199744 140282 199753
rect 140410 199744 140466 199753
rect 140226 199679 140282 199688
rect 140332 199702 140410 199730
rect 140240 196081 140268 199679
rect 140226 196072 140282 196081
rect 140226 196007 140282 196016
rect 140228 195900 140280 195906
rect 140228 195842 140280 195848
rect 140240 195702 140268 195842
rect 140228 195696 140280 195702
rect 140228 195638 140280 195644
rect 140332 194206 140360 199702
rect 140562 199696 140590 200124
rect 140654 199923 140682 200124
rect 140640 199914 140696 199923
rect 140746 199918 140774 200124
rect 140838 199918 140866 200124
rect 140930 199923 140958 200124
rect 140640 199849 140696 199858
rect 140734 199912 140786 199918
rect 140734 199854 140786 199860
rect 140826 199912 140878 199918
rect 140826 199854 140878 199860
rect 140916 199914 140972 199923
rect 141022 199918 141050 200124
rect 140916 199849 140972 199858
rect 141010 199912 141062 199918
rect 141010 199854 141062 199860
rect 140688 199776 140740 199782
rect 140688 199718 140740 199724
rect 140964 199776 141016 199782
rect 141114 199730 141142 200124
rect 140964 199718 141016 199724
rect 140410 199679 140466 199688
rect 140516 199668 140590 199696
rect 140412 199640 140464 199646
rect 140412 199582 140464 199588
rect 140424 196897 140452 199582
rect 140410 196888 140466 196897
rect 140410 196823 140466 196832
rect 140516 195158 140544 199668
rect 140594 196888 140650 196897
rect 140594 196823 140650 196832
rect 140504 195152 140556 195158
rect 140504 195094 140556 195100
rect 140320 194200 140372 194206
rect 140320 194142 140372 194148
rect 140148 191806 140360 191834
rect 140228 191140 140280 191146
rect 140228 191082 140280 191088
rect 139952 187400 140004 187406
rect 139952 187342 140004 187348
rect 139044 186286 139348 186314
rect 139596 186286 140176 186314
rect 139320 151094 139348 186286
rect 139308 151088 139360 151094
rect 139308 151030 139360 151036
rect 138662 147656 138718 147665
rect 138662 147591 138718 147600
rect 138572 147348 138624 147354
rect 138572 147290 138624 147296
rect 140148 146946 140176 186286
rect 140240 154086 140268 191082
rect 140332 186314 140360 191806
rect 140608 191146 140636 196823
rect 140700 194342 140728 199718
rect 140780 199708 140832 199714
rect 140780 199650 140832 199656
rect 140872 199708 140924 199714
rect 140872 199650 140924 199656
rect 140792 196489 140820 199650
rect 140884 196722 140912 199650
rect 140872 196716 140924 196722
rect 140872 196658 140924 196664
rect 140976 196654 141004 199718
rect 141068 199702 141142 199730
rect 140964 196648 141016 196654
rect 140964 196590 141016 196596
rect 140778 196480 140834 196489
rect 140778 196415 140834 196424
rect 140872 195832 140924 195838
rect 140872 195774 140924 195780
rect 140884 195226 140912 195774
rect 140872 195220 140924 195226
rect 140872 195162 140924 195168
rect 141068 194546 141096 199702
rect 141206 199594 141234 200124
rect 141298 199696 141326 200124
rect 141390 199764 141418 200124
rect 141482 199923 141510 200124
rect 141468 199914 141524 199923
rect 141468 199849 141524 199858
rect 141574 199850 141602 200124
rect 141666 199923 141694 200124
rect 141652 199914 141708 199923
rect 141758 199918 141786 200124
rect 141850 199918 141878 200124
rect 141562 199844 141614 199850
rect 141652 199849 141708 199858
rect 141746 199912 141798 199918
rect 141746 199854 141798 199860
rect 141838 199912 141890 199918
rect 141838 199854 141890 199860
rect 141562 199786 141614 199792
rect 141390 199736 141464 199764
rect 141298 199668 141372 199696
rect 141206 199566 141280 199594
rect 141252 196314 141280 199566
rect 141240 196308 141292 196314
rect 141240 196250 141292 196256
rect 141056 194540 141108 194546
rect 141056 194482 141108 194488
rect 140688 194336 140740 194342
rect 140688 194278 140740 194284
rect 141344 193866 141372 199668
rect 141332 193860 141384 193866
rect 141332 193802 141384 193808
rect 141436 191834 141464 199736
rect 141942 199730 141970 200124
rect 142034 199918 142062 200124
rect 142126 199918 142154 200124
rect 142218 199918 142246 200124
rect 142310 199918 142338 200124
rect 142402 199918 142430 200124
rect 142022 199912 142074 199918
rect 142022 199854 142074 199860
rect 142114 199912 142166 199918
rect 142114 199854 142166 199860
rect 142206 199912 142258 199918
rect 142206 199854 142258 199860
rect 142298 199912 142350 199918
rect 142298 199854 142350 199860
rect 142390 199912 142442 199918
rect 142390 199854 142442 199860
rect 142252 199776 142304 199782
rect 141516 199708 141568 199714
rect 141516 199650 141568 199656
rect 141896 199702 141970 199730
rect 142066 199744 142122 199753
rect 141528 196897 141556 199650
rect 141608 199640 141660 199646
rect 141608 199582 141660 199588
rect 141792 199640 141844 199646
rect 141792 199582 141844 199588
rect 141620 199481 141648 199582
rect 141606 199472 141662 199481
rect 141606 199407 141662 199416
rect 141698 198248 141754 198257
rect 141698 198183 141754 198192
rect 141514 196888 141570 196897
rect 141514 196823 141570 196832
rect 141712 191834 141740 198183
rect 141804 196874 141832 199582
rect 141896 197538 141924 199702
rect 142066 199679 142122 199688
rect 142250 199744 142252 199753
rect 142304 199744 142306 199753
rect 142250 199679 142306 199688
rect 142494 199696 142522 200124
rect 142586 199764 142614 200124
rect 142678 199923 142706 200124
rect 142664 199914 142720 199923
rect 142770 199918 142798 200124
rect 142862 199923 142890 200124
rect 142664 199849 142720 199858
rect 142758 199912 142810 199918
rect 142758 199854 142810 199860
rect 142848 199914 142904 199923
rect 142848 199849 142904 199858
rect 142712 199776 142764 199782
rect 142586 199736 142660 199764
rect 141976 199640 142028 199646
rect 141976 199582 142028 199588
rect 141884 197532 141936 197538
rect 141884 197474 141936 197480
rect 141884 197260 141936 197266
rect 141884 197202 141936 197208
rect 141896 197062 141924 197202
rect 141884 197056 141936 197062
rect 141884 196998 141936 197004
rect 141804 196846 141924 196874
rect 141792 196716 141844 196722
rect 141792 196658 141844 196664
rect 141068 191806 141464 191834
rect 141620 191806 141740 191834
rect 141068 191622 141096 191806
rect 141056 191616 141108 191622
rect 141056 191558 141108 191564
rect 140596 191140 140648 191146
rect 140596 191082 140648 191088
rect 141620 187066 141648 191806
rect 141608 187060 141660 187066
rect 141608 187002 141660 187008
rect 141804 186946 141832 196658
rect 141896 194206 141924 196846
rect 141884 194200 141936 194206
rect 141884 194142 141936 194148
rect 140976 186918 141832 186946
rect 140332 186286 140452 186314
rect 140228 154080 140280 154086
rect 140228 154022 140280 154028
rect 140424 154018 140452 186286
rect 140412 154012 140464 154018
rect 140412 153954 140464 153960
rect 140976 151774 141004 186918
rect 141988 186314 142016 199582
rect 142080 197266 142108 199679
rect 142494 199668 142568 199696
rect 142252 199640 142304 199646
rect 142252 199582 142304 199588
rect 142158 199336 142214 199345
rect 142158 199271 142160 199280
rect 142212 199271 142214 199280
rect 142160 199242 142212 199248
rect 142158 199200 142214 199209
rect 142158 199135 142214 199144
rect 142172 198694 142200 199135
rect 142160 198688 142212 198694
rect 142160 198630 142212 198636
rect 142264 198014 142292 199582
rect 142344 199572 142396 199578
rect 142344 199514 142396 199520
rect 142356 198150 142384 199514
rect 142344 198144 142396 198150
rect 142344 198086 142396 198092
rect 142252 198008 142304 198014
rect 142252 197950 142304 197956
rect 142068 197260 142120 197266
rect 142068 197202 142120 197208
rect 142160 196648 142212 196654
rect 142160 196590 142212 196596
rect 142068 196308 142120 196314
rect 142068 196250 142120 196256
rect 141620 186286 142016 186314
rect 140964 151768 141016 151774
rect 140964 151710 141016 151716
rect 140136 146940 140188 146946
rect 140136 146882 140188 146888
rect 138940 144492 138992 144498
rect 138940 144434 138992 144440
rect 138308 142126 138428 142154
rect 138308 140078 138336 142126
rect 138388 141840 138440 141846
rect 138388 141782 138440 141788
rect 138296 140072 138348 140078
rect 138296 140014 138348 140020
rect 138400 139890 138428 141782
rect 138952 139890 138980 144434
rect 141148 143200 141200 143206
rect 141148 143142 141200 143148
rect 140044 142996 140096 143002
rect 140044 142938 140096 142944
rect 139490 141536 139546 141545
rect 139490 141471 139546 141480
rect 139504 139890 139532 141471
rect 140056 139890 140084 142938
rect 140780 142928 140832 142934
rect 140780 142870 140832 142876
rect 140792 139890 140820 142870
rect 141160 139890 141188 143142
rect 141620 141778 141648 186286
rect 142080 180794 142108 196250
rect 141896 180766 142108 180794
rect 141896 150958 141924 180766
rect 141884 150952 141936 150958
rect 141884 150894 141936 150900
rect 142172 147121 142200 196590
rect 142540 191026 142568 199668
rect 142632 192710 142660 199736
rect 142954 199764 142982 200124
rect 143046 199923 143074 200124
rect 143032 199914 143088 199923
rect 143138 199918 143166 200124
rect 143230 199918 143258 200124
rect 143032 199849 143088 199858
rect 143126 199912 143178 199918
rect 143126 199854 143178 199860
rect 143218 199912 143270 199918
rect 143218 199854 143270 199860
rect 143322 199850 143350 200124
rect 143414 199918 143442 200124
rect 143506 199918 143534 200124
rect 143402 199912 143454 199918
rect 143402 199854 143454 199860
rect 143494 199912 143546 199918
rect 143494 199854 143546 199860
rect 143310 199844 143362 199850
rect 143310 199786 143362 199792
rect 142712 199718 142764 199724
rect 142908 199736 142982 199764
rect 143448 199776 143500 199782
rect 142724 196625 142752 199718
rect 142802 197432 142858 197441
rect 142802 197367 142858 197376
rect 142710 196616 142766 196625
rect 142710 196551 142766 196560
rect 142816 192778 142844 197367
rect 142908 195634 142936 199736
rect 143598 199764 143626 200124
rect 143690 199918 143718 200124
rect 143782 199918 143810 200124
rect 143874 199923 143902 200124
rect 143678 199912 143730 199918
rect 143678 199854 143730 199860
rect 143770 199912 143822 199918
rect 143770 199854 143822 199860
rect 143860 199914 143916 199923
rect 143966 199918 143994 200124
rect 144058 199918 144086 200124
rect 144150 199918 144178 200124
rect 144242 199918 144270 200124
rect 144334 199918 144362 200124
rect 144426 199923 144454 200124
rect 143860 199849 143916 199858
rect 143954 199912 144006 199918
rect 143954 199854 144006 199860
rect 144046 199912 144098 199918
rect 144046 199854 144098 199860
rect 144138 199912 144190 199918
rect 144138 199854 144190 199860
rect 144230 199912 144282 199918
rect 144230 199854 144282 199860
rect 144322 199912 144374 199918
rect 144322 199854 144374 199860
rect 144412 199914 144468 199923
rect 144412 199849 144468 199858
rect 143448 199718 143500 199724
rect 143552 199736 143626 199764
rect 143816 199776 143868 199782
rect 143080 199640 143132 199646
rect 143080 199582 143132 199588
rect 143354 199608 143410 199617
rect 142986 197432 143042 197441
rect 142986 197367 143042 197376
rect 142896 195628 142948 195634
rect 142896 195570 142948 195576
rect 142804 192772 142856 192778
rect 142804 192714 142856 192720
rect 142620 192704 142672 192710
rect 142620 192646 142672 192652
rect 142540 190998 142752 191026
rect 142620 190936 142672 190942
rect 142620 190878 142672 190884
rect 142528 188420 142580 188426
rect 142528 188362 142580 188368
rect 142540 148918 142568 188362
rect 142528 148912 142580 148918
rect 142528 148854 142580 148860
rect 142632 148782 142660 190878
rect 142724 186314 142752 190998
rect 143000 190942 143028 197367
rect 143092 196246 143120 199582
rect 143172 199572 143224 199578
rect 143172 199514 143224 199520
rect 143264 199572 143316 199578
rect 143354 199543 143410 199552
rect 143264 199514 143316 199520
rect 143080 196240 143132 196246
rect 143080 196182 143132 196188
rect 143184 194002 143212 199514
rect 143172 193996 143224 194002
rect 143172 193938 143224 193944
rect 142988 190936 143040 190942
rect 142988 190878 143040 190884
rect 143276 188426 143304 199514
rect 143368 198354 143396 199543
rect 143356 198348 143408 198354
rect 143356 198290 143408 198296
rect 143356 198076 143408 198082
rect 143356 198018 143408 198024
rect 143368 195673 143396 198018
rect 143460 195906 143488 199718
rect 143448 195900 143500 195906
rect 143448 195842 143500 195848
rect 143354 195664 143410 195673
rect 143354 195599 143410 195608
rect 143552 195242 143580 199736
rect 143816 199718 143868 199724
rect 143908 199776 143960 199782
rect 143908 199718 143960 199724
rect 144276 199776 144328 199782
rect 144276 199718 144328 199724
rect 144368 199776 144420 199782
rect 144518 199764 144546 200124
rect 144368 199718 144420 199724
rect 144472 199736 144546 199764
rect 144610 199764 144638 200124
rect 144702 199923 144730 200124
rect 144688 199914 144744 199923
rect 144794 199918 144822 200124
rect 144688 199849 144744 199858
rect 144782 199912 144834 199918
rect 144782 199854 144834 199860
rect 144736 199776 144788 199782
rect 144610 199736 144684 199764
rect 143632 199640 143684 199646
rect 143632 199582 143684 199588
rect 143644 199209 143672 199582
rect 143722 199472 143778 199481
rect 143722 199407 143724 199416
rect 143776 199407 143778 199416
rect 143724 199378 143776 199384
rect 143630 199200 143686 199209
rect 143630 199135 143686 199144
rect 143630 199064 143686 199073
rect 143630 198999 143686 199008
rect 143644 198626 143672 198999
rect 143632 198620 143684 198626
rect 143632 198562 143684 198568
rect 143552 195214 143764 195242
rect 143632 195152 143684 195158
rect 143632 195094 143684 195100
rect 143540 194540 143592 194546
rect 143540 194482 143592 194488
rect 143264 188420 143316 188426
rect 143264 188362 143316 188368
rect 142724 186286 142936 186314
rect 142908 152522 142936 186286
rect 142896 152516 142948 152522
rect 142896 152458 142948 152464
rect 142620 148776 142672 148782
rect 142620 148718 142672 148724
rect 143552 147393 143580 194482
rect 143538 147384 143594 147393
rect 143538 147319 143594 147328
rect 142158 147112 142214 147121
rect 142158 147047 142214 147056
rect 143644 147014 143672 195094
rect 143736 193186 143764 195214
rect 143724 193180 143776 193186
rect 143724 193122 143776 193128
rect 143828 192574 143856 199718
rect 143920 197354 143948 199718
rect 144000 199708 144052 199714
rect 144000 199650 144052 199656
rect 144012 197878 144040 199650
rect 144182 199472 144238 199481
rect 144182 199407 144238 199416
rect 144000 197872 144052 197878
rect 144000 197814 144052 197820
rect 144196 197810 144224 199407
rect 144184 197804 144236 197810
rect 144184 197746 144236 197752
rect 144288 197354 144316 199718
rect 144380 198422 144408 199718
rect 144472 198744 144500 199736
rect 144552 199572 144604 199578
rect 144552 199514 144604 199520
rect 144564 198937 144592 199514
rect 144550 198928 144606 198937
rect 144550 198863 144606 198872
rect 144472 198716 144592 198744
rect 144368 198416 144420 198422
rect 144368 198358 144420 198364
rect 143920 197326 144132 197354
rect 144000 196308 144052 196314
rect 144000 196250 144052 196256
rect 143908 193860 143960 193866
rect 143908 193802 143960 193808
rect 143816 192568 143868 192574
rect 143816 192510 143868 192516
rect 143920 189922 143948 193802
rect 143908 189916 143960 189922
rect 143908 189858 143960 189864
rect 144012 147218 144040 196250
rect 144104 190058 144132 197326
rect 144196 197326 144316 197354
rect 144196 195090 144224 197326
rect 144274 196072 144330 196081
rect 144274 196007 144330 196016
rect 144288 195294 144316 196007
rect 144276 195288 144328 195294
rect 144276 195230 144328 195236
rect 144184 195084 144236 195090
rect 144184 195026 144236 195032
rect 144564 190126 144592 198716
rect 144656 198558 144684 199736
rect 144886 199764 144914 200124
rect 144978 199918 145006 200124
rect 144966 199912 145018 199918
rect 144966 199854 145018 199860
rect 145070 199764 145098 200124
rect 145162 199782 145190 200124
rect 144736 199718 144788 199724
rect 144840 199736 144914 199764
rect 145024 199753 145098 199764
rect 145010 199744 145098 199753
rect 144644 198552 144696 198558
rect 144644 198494 144696 198500
rect 144748 196314 144776 199718
rect 144736 196308 144788 196314
rect 144736 196250 144788 196256
rect 144552 190120 144604 190126
rect 144552 190062 144604 190068
rect 144092 190052 144144 190058
rect 144092 189994 144144 190000
rect 144840 189854 144868 199736
rect 145066 199736 145098 199744
rect 145150 199776 145202 199782
rect 145150 199718 145202 199724
rect 145010 199679 145066 199688
rect 145104 199640 145156 199646
rect 145254 199628 145282 200124
rect 145104 199582 145156 199588
rect 145208 199600 145282 199628
rect 145012 199572 145064 199578
rect 145012 199514 145064 199520
rect 144920 199504 144972 199510
rect 144920 199446 144972 199452
rect 144932 199209 144960 199446
rect 144918 199200 144974 199209
rect 144918 199135 144974 199144
rect 145024 198082 145052 199514
rect 145012 198076 145064 198082
rect 145012 198018 145064 198024
rect 144920 197260 144972 197266
rect 144920 197202 144972 197208
rect 144828 189848 144880 189854
rect 144828 189790 144880 189796
rect 144932 151026 144960 197202
rect 145116 191834 145144 199582
rect 145208 195809 145236 199600
rect 145346 199560 145374 200124
rect 145438 199923 145466 200124
rect 145424 199914 145480 199923
rect 145530 199918 145558 200124
rect 145622 199918 145650 200124
rect 145714 199918 145742 200124
rect 145806 199918 145834 200124
rect 145898 199923 145926 200124
rect 145424 199849 145480 199858
rect 145518 199912 145570 199918
rect 145518 199854 145570 199860
rect 145610 199912 145662 199918
rect 145610 199854 145662 199860
rect 145702 199912 145754 199918
rect 145702 199854 145754 199860
rect 145794 199912 145846 199918
rect 145794 199854 145846 199860
rect 145884 199914 145940 199923
rect 145884 199849 145940 199858
rect 145990 199782 146018 200124
rect 146082 199923 146110 200124
rect 146068 199914 146124 199923
rect 146068 199849 146124 199858
rect 146174 199782 146202 200124
rect 146266 199918 146294 200124
rect 146358 199918 146386 200124
rect 146254 199912 146306 199918
rect 146254 199854 146306 199860
rect 146346 199912 146398 199918
rect 146346 199854 146398 199860
rect 145472 199776 145524 199782
rect 145978 199776 146030 199782
rect 145472 199718 145524 199724
rect 145746 199744 145802 199753
rect 145300 199532 145374 199560
rect 145194 195800 145250 195809
rect 145194 195735 145250 195744
rect 145300 193118 145328 199532
rect 145378 199200 145434 199209
rect 145378 199135 145380 199144
rect 145432 199135 145434 199144
rect 145380 199106 145432 199112
rect 145288 193112 145340 193118
rect 145288 193054 145340 193060
rect 145116 191806 145420 191834
rect 145392 186998 145420 191806
rect 145380 186992 145432 186998
rect 145380 186934 145432 186940
rect 145484 186314 145512 199718
rect 145564 199708 145616 199714
rect 145564 199650 145616 199656
rect 145656 199708 145708 199714
rect 145978 199718 146030 199724
rect 146162 199776 146214 199782
rect 146162 199718 146214 199724
rect 146450 199730 146478 200124
rect 146542 199923 146570 200124
rect 146528 199914 146584 199923
rect 146528 199849 146584 199858
rect 146634 199764 146662 200124
rect 146726 199918 146754 200124
rect 146714 199912 146766 199918
rect 146714 199854 146766 199860
rect 146818 199764 146846 200124
rect 146910 199923 146938 200124
rect 146896 199914 146952 199923
rect 147002 199918 147030 200124
rect 146896 199849 146952 199858
rect 146990 199912 147042 199918
rect 146990 199854 147042 199860
rect 147094 199764 147122 200124
rect 146588 199753 146662 199764
rect 146574 199744 146662 199753
rect 146450 199714 146524 199730
rect 145746 199679 145802 199688
rect 145840 199708 145892 199714
rect 145656 199650 145708 199656
rect 145576 195498 145604 199650
rect 145668 196858 145696 199650
rect 145760 199646 145788 199679
rect 146450 199708 146536 199714
rect 146450 199702 146484 199708
rect 145840 199650 145892 199656
rect 146630 199736 146662 199744
rect 146772 199736 146846 199764
rect 147048 199736 147122 199764
rect 146574 199679 146630 199688
rect 146484 199650 146536 199656
rect 145748 199640 145800 199646
rect 145748 199582 145800 199588
rect 145748 199504 145800 199510
rect 145748 199446 145800 199452
rect 145760 198762 145788 199446
rect 145748 198756 145800 198762
rect 145748 198698 145800 198704
rect 145746 198656 145802 198665
rect 145746 198591 145802 198600
rect 145760 197062 145788 198591
rect 145748 197056 145800 197062
rect 145748 196998 145800 197004
rect 145656 196852 145708 196858
rect 145656 196794 145708 196800
rect 145852 195974 145880 199650
rect 145932 199640 145984 199646
rect 145932 199582 145984 199588
rect 146024 199640 146076 199646
rect 146024 199582 146076 199588
rect 146208 199640 146260 199646
rect 146392 199640 146444 199646
rect 146208 199582 146260 199588
rect 146312 199588 146392 199594
rect 146668 199640 146720 199646
rect 146312 199582 146444 199588
rect 146482 199608 146538 199617
rect 145840 195968 145892 195974
rect 145840 195910 145892 195916
rect 145564 195492 145616 195498
rect 145564 195434 145616 195440
rect 145944 195362 145972 199582
rect 146036 198830 146064 199582
rect 146114 199200 146170 199209
rect 146114 199135 146170 199144
rect 146128 199102 146156 199135
rect 146116 199096 146168 199102
rect 146116 199038 146168 199044
rect 146024 198824 146076 198830
rect 146024 198766 146076 198772
rect 145932 195356 145984 195362
rect 145932 195298 145984 195304
rect 146220 192982 146248 199582
rect 146312 199566 146432 199582
rect 146312 196722 146340 199566
rect 146668 199582 146720 199588
rect 146482 199543 146538 199552
rect 146576 199572 146628 199578
rect 146392 199504 146444 199510
rect 146392 199446 146444 199452
rect 146300 196716 146352 196722
rect 146300 196658 146352 196664
rect 146208 192976 146260 192982
rect 146208 192918 146260 192924
rect 145300 186286 145512 186314
rect 146404 186314 146432 199446
rect 146496 195702 146524 199543
rect 146576 199514 146628 199520
rect 146588 199481 146616 199514
rect 146574 199472 146630 199481
rect 146574 199407 146630 199416
rect 146484 195696 146536 195702
rect 146484 195638 146536 195644
rect 146680 193214 146708 199582
rect 146772 199034 146800 199736
rect 147048 199730 147076 199736
rect 147002 199702 147076 199730
rect 147002 199696 147030 199702
rect 146956 199668 147030 199696
rect 146956 199560 146984 199668
rect 147186 199594 147214 200124
rect 147278 199923 147306 200124
rect 147264 199914 147320 199923
rect 147264 199849 147320 199858
rect 147370 199782 147398 200124
rect 147358 199776 147410 199782
rect 147358 199718 147410 199724
rect 147140 199578 147214 199594
rect 147312 199640 147364 199646
rect 147462 199628 147490 200124
rect 147554 199764 147582 200124
rect 147646 199918 147674 200124
rect 147738 199918 147766 200124
rect 147830 199918 147858 200124
rect 147922 199918 147950 200124
rect 147634 199912 147686 199918
rect 147634 199854 147686 199860
rect 147726 199912 147778 199918
rect 147726 199854 147778 199860
rect 147818 199912 147870 199918
rect 147818 199854 147870 199860
rect 147910 199912 147962 199918
rect 147910 199854 147962 199860
rect 147554 199753 147628 199764
rect 147554 199744 147642 199753
rect 147554 199736 147586 199744
rect 148014 199730 148042 200124
rect 148106 199918 148134 200124
rect 148198 199918 148226 200124
rect 148290 199918 148318 200124
rect 148094 199912 148146 199918
rect 148094 199854 148146 199860
rect 148186 199912 148238 199918
rect 148186 199854 148238 199860
rect 148278 199912 148330 199918
rect 148278 199854 148330 199860
rect 148382 199850 148410 200124
rect 148370 199844 148422 199850
rect 148370 199786 148422 199792
rect 148140 199776 148192 199782
rect 147586 199679 147642 199688
rect 147772 199708 147824 199714
rect 147772 199650 147824 199656
rect 147864 199708 147916 199714
rect 148014 199702 148088 199730
rect 148140 199718 148192 199724
rect 148232 199776 148284 199782
rect 148232 199718 148284 199724
rect 147864 199650 147916 199656
rect 147680 199640 147732 199646
rect 147462 199600 147536 199628
rect 147312 199582 147364 199588
rect 146864 199532 146984 199560
rect 147128 199572 147214 199578
rect 146864 199306 146892 199532
rect 147180 199566 147214 199572
rect 147128 199514 147180 199520
rect 147126 199472 147182 199481
rect 146944 199436 146996 199442
rect 147126 199407 147182 199416
rect 146944 199378 146996 199384
rect 146852 199300 146904 199306
rect 146852 199242 146904 199248
rect 146760 199028 146812 199034
rect 146760 198970 146812 198976
rect 146956 196840 146984 199378
rect 146588 193186 146708 193214
rect 146772 196812 146984 196840
rect 146588 192642 146616 193186
rect 146576 192636 146628 192642
rect 146576 192578 146628 192584
rect 146772 191214 146800 196812
rect 146852 196716 146904 196722
rect 146852 196658 146904 196664
rect 147036 196716 147088 196722
rect 147036 196658 147088 196664
rect 146760 191208 146812 191214
rect 146760 191150 146812 191156
rect 146864 191078 146892 196658
rect 146944 195288 146996 195294
rect 146944 195230 146996 195236
rect 146852 191072 146904 191078
rect 146852 191014 146904 191020
rect 146404 186286 146892 186314
rect 145300 153950 145328 186286
rect 145288 153944 145340 153950
rect 145288 153886 145340 153892
rect 144920 151020 144972 151026
rect 144920 150962 144972 150968
rect 144000 147212 144052 147218
rect 144000 147154 144052 147160
rect 143632 147008 143684 147014
rect 143632 146950 143684 146956
rect 142250 146160 142306 146169
rect 142250 146095 142306 146104
rect 142160 145988 142212 145994
rect 142160 145930 142212 145936
rect 141700 143064 141752 143070
rect 141700 143006 141752 143012
rect 141608 141772 141660 141778
rect 141608 141714 141660 141720
rect 141712 139890 141740 143006
rect 142172 140758 142200 145930
rect 142160 140752 142212 140758
rect 142160 140694 142212 140700
rect 142264 139890 142292 146095
rect 144366 146024 144422 146033
rect 144366 145959 144422 145968
rect 143908 144356 143960 144362
rect 143908 144298 143960 144304
rect 143540 142860 143592 142866
rect 143540 142802 143592 142808
rect 142804 140752 142856 140758
rect 142804 140694 142856 140700
rect 142816 139890 142844 140694
rect 143552 139890 143580 142802
rect 143920 139890 143948 144298
rect 144380 139890 144408 145959
rect 146758 145888 146814 145897
rect 146758 145823 146814 145832
rect 146298 145616 146354 145625
rect 146298 145551 146354 145560
rect 145562 144800 145618 144809
rect 145562 144735 145618 144744
rect 145102 143440 145158 143449
rect 145102 143375 145158 143384
rect 145116 139890 145144 143375
rect 145576 139890 145604 144735
rect 146312 139890 146340 145551
rect 146666 143032 146722 143041
rect 146666 142967 146722 142976
rect 146680 139890 146708 142967
rect 146772 140740 146800 145823
rect 146864 141642 146892 186286
rect 146956 143313 146984 195230
rect 147048 149054 147076 196658
rect 147140 151814 147168 199407
rect 147324 198898 147352 199582
rect 147312 198892 147364 198898
rect 147312 198834 147364 198840
rect 147508 196654 147536 199600
rect 147680 199582 147732 199588
rect 147588 199572 147640 199578
rect 147588 199514 147640 199520
rect 147496 196648 147548 196654
rect 147496 196590 147548 196596
rect 147494 196480 147550 196489
rect 147494 196415 147550 196424
rect 147508 192302 147536 196415
rect 147600 195786 147628 199514
rect 147692 199345 147720 199582
rect 147678 199336 147734 199345
rect 147678 199271 147734 199280
rect 147600 195758 147720 195786
rect 147586 195664 147642 195673
rect 147586 195599 147642 195608
rect 147496 192296 147548 192302
rect 147496 192238 147548 192244
rect 147600 186425 147628 195599
rect 147692 194410 147720 195758
rect 147784 194478 147812 199650
rect 147876 199481 147904 199650
rect 147956 199640 148008 199646
rect 147956 199582 148008 199588
rect 147862 199472 147918 199481
rect 147862 199407 147918 199416
rect 147968 195838 147996 199582
rect 147956 195832 148008 195838
rect 147956 195774 148008 195780
rect 147772 194472 147824 194478
rect 147772 194414 147824 194420
rect 147680 194404 147732 194410
rect 147680 194346 147732 194352
rect 147956 194268 148008 194274
rect 147956 194210 148008 194216
rect 147586 186416 147642 186425
rect 147586 186351 147642 186360
rect 147140 151786 147260 151814
rect 147036 149048 147088 149054
rect 147036 148990 147088 148996
rect 146942 143304 146998 143313
rect 146942 143239 146998 143248
rect 147232 141710 147260 151786
rect 147968 148306 147996 194210
rect 148060 149734 148088 199702
rect 148152 198529 148180 199718
rect 148244 199238 148272 199718
rect 148474 199696 148502 200124
rect 148566 199918 148594 200124
rect 148554 199912 148606 199918
rect 148554 199854 148606 199860
rect 148658 199753 148686 200124
rect 148750 199764 148778 200124
rect 148842 199918 148870 200124
rect 148830 199912 148882 199918
rect 148830 199854 148882 199860
rect 148934 199764 148962 200124
rect 148428 199668 148502 199696
rect 148644 199744 148700 199753
rect 148750 199736 148824 199764
rect 148888 199753 148962 199764
rect 148644 199679 148700 199688
rect 148324 199572 148376 199578
rect 148324 199514 148376 199520
rect 148232 199232 148284 199238
rect 148232 199174 148284 199180
rect 148138 198520 148194 198529
rect 148138 198455 148194 198464
rect 148336 196704 148364 199514
rect 148428 196926 148456 199668
rect 148600 199640 148652 199646
rect 148600 199582 148652 199588
rect 148692 199640 148744 199646
rect 148692 199582 148744 199588
rect 148416 196920 148468 196926
rect 148416 196862 148468 196868
rect 148152 196676 148364 196704
rect 148048 149728 148100 149734
rect 148048 149670 148100 149676
rect 147956 148300 148008 148306
rect 147956 148242 148008 148248
rect 147772 144560 147824 144566
rect 147772 144502 147824 144508
rect 147220 141704 147272 141710
rect 147220 141646 147272 141652
rect 146852 141636 146904 141642
rect 146852 141578 146904 141584
rect 146772 140712 147168 140740
rect 147140 139890 147168 140712
rect 147784 139890 147812 144502
rect 148152 140214 148180 196676
rect 148232 194472 148284 194478
rect 148232 194414 148284 194420
rect 148244 141506 148272 194414
rect 148612 194274 148640 199582
rect 148600 194268 148652 194274
rect 148600 194210 148652 194216
rect 148704 193214 148732 199582
rect 148796 195430 148824 199736
rect 148874 199744 148962 199753
rect 148930 199736 148962 199744
rect 148874 199679 148930 199688
rect 149026 199560 149054 200124
rect 149118 199696 149146 200124
rect 149210 199918 149238 200124
rect 149198 199912 149250 199918
rect 149198 199854 149250 199860
rect 149302 199782 149330 200124
rect 149394 199918 149422 200124
rect 149486 199918 149514 200124
rect 149578 199918 149606 200124
rect 149670 199918 149698 200124
rect 149382 199912 149434 199918
rect 149382 199854 149434 199860
rect 149474 199912 149526 199918
rect 149474 199854 149526 199860
rect 149566 199912 149618 199918
rect 149566 199854 149618 199860
rect 149658 199912 149710 199918
rect 149658 199854 149710 199860
rect 149762 199850 149790 200124
rect 149854 199918 149882 200124
rect 149842 199912 149894 199918
rect 149842 199854 149894 199860
rect 149946 199850 149974 200124
rect 150038 199918 150066 200124
rect 150130 199918 150158 200124
rect 150026 199912 150078 199918
rect 150026 199854 150078 199860
rect 150118 199912 150170 199918
rect 150118 199854 150170 199860
rect 149750 199844 149802 199850
rect 149750 199786 149802 199792
rect 149934 199844 149986 199850
rect 149934 199786 149986 199792
rect 149290 199776 149342 199782
rect 150222 199730 150250 200124
rect 149290 199718 149342 199724
rect 149612 199708 149664 199714
rect 149118 199668 149192 199696
rect 149026 199532 149100 199560
rect 148876 199504 148928 199510
rect 148876 199446 148928 199452
rect 148784 195424 148836 195430
rect 148784 195366 148836 195372
rect 148888 193214 148916 199446
rect 149072 195770 149100 199532
rect 149164 197130 149192 199668
rect 149612 199650 149664 199656
rect 149704 199708 149756 199714
rect 149704 199650 149756 199656
rect 149796 199708 149848 199714
rect 149796 199650 149848 199656
rect 149888 199708 149940 199714
rect 149888 199650 149940 199656
rect 150176 199702 150250 199730
rect 149336 199572 149388 199578
rect 149336 199514 149388 199520
rect 149520 199572 149572 199578
rect 149520 199514 149572 199520
rect 149348 198393 149376 199514
rect 149428 199436 149480 199442
rect 149428 199378 149480 199384
rect 149334 198384 149390 198393
rect 149334 198319 149390 198328
rect 149152 197124 149204 197130
rect 149152 197066 149204 197072
rect 149336 196784 149388 196790
rect 149336 196726 149388 196732
rect 149060 195764 149112 195770
rect 149060 195706 149112 195712
rect 148704 193186 148824 193214
rect 148888 193186 149192 193214
rect 148796 180794 148824 193186
rect 149164 192370 149192 193186
rect 149152 192364 149204 192370
rect 149152 192306 149204 192312
rect 148428 180766 148824 180794
rect 148428 145654 148456 180766
rect 149348 148510 149376 196726
rect 149336 148504 149388 148510
rect 149336 148446 149388 148452
rect 149244 146056 149296 146062
rect 149244 145998 149296 146004
rect 149060 145920 149112 145926
rect 149060 145862 149112 145868
rect 148416 145648 148468 145654
rect 148416 145590 148468 145596
rect 148322 143168 148378 143177
rect 148322 143103 148378 143112
rect 148232 141500 148284 141506
rect 148232 141442 148284 141448
rect 148140 140208 148192 140214
rect 148140 140150 148192 140156
rect 148336 139890 148364 143103
rect 149072 139890 149100 145862
rect 149256 140758 149284 145998
rect 149244 140752 149296 140758
rect 149244 140694 149296 140700
rect 130672 139862 131008 139890
rect 131500 139862 131560 139890
rect 131776 139862 132112 139890
rect 132512 139862 132664 139890
rect 132880 139862 133216 139890
rect 133432 139862 133768 139890
rect 133984 139862 134320 139890
rect 134536 139862 134872 139890
rect 135364 139862 135424 139890
rect 135640 139862 135976 139890
rect 136192 139862 136528 139890
rect 136744 139862 137080 139890
rect 137296 139862 137632 139890
rect 138032 139862 138184 139890
rect 138400 139862 138736 139890
rect 138952 139862 139288 139890
rect 139504 139862 139840 139890
rect 140056 139862 140392 139890
rect 140792 139862 140944 139890
rect 141160 139862 141496 139890
rect 141712 139862 142048 139890
rect 142264 139862 142600 139890
rect 142816 139862 143152 139890
rect 143552 139862 143704 139890
rect 143920 139862 144256 139890
rect 144380 139862 144808 139890
rect 145116 139862 145360 139890
rect 145576 139862 145912 139890
rect 146312 139862 146464 139890
rect 146680 139862 147016 139890
rect 147140 139862 147568 139890
rect 147784 139862 148120 139890
rect 148336 139862 148672 139890
rect 149072 139862 149224 139890
rect 149440 139369 149468 199378
rect 149532 196058 149560 199514
rect 149624 198966 149652 199650
rect 149612 198960 149664 198966
rect 149612 198902 149664 198908
rect 149716 196722 149744 199650
rect 149704 196716 149756 196722
rect 149704 196658 149756 196664
rect 149532 196030 149744 196058
rect 149520 195424 149572 195430
rect 149520 195366 149572 195372
rect 149532 189786 149560 195366
rect 149612 195356 149664 195362
rect 149612 195298 149664 195304
rect 149520 189780 149572 189786
rect 149520 189722 149572 189728
rect 149624 141574 149652 195298
rect 149716 145858 149744 196030
rect 149808 191418 149836 199650
rect 149900 196790 149928 199650
rect 149980 199504 150032 199510
rect 149980 199446 150032 199452
rect 149888 196784 149940 196790
rect 149888 196726 149940 196732
rect 149992 195430 150020 199446
rect 149980 195424 150032 195430
rect 149980 195366 150032 195372
rect 150176 195362 150204 199702
rect 150314 199628 150342 200124
rect 150406 199918 150434 200124
rect 150498 199918 150526 200124
rect 150590 199923 150618 200124
rect 150394 199912 150446 199918
rect 150394 199854 150446 199860
rect 150486 199912 150538 199918
rect 150486 199854 150538 199860
rect 150576 199914 150632 199923
rect 150576 199849 150632 199858
rect 150578 199776 150630 199782
rect 150452 199753 150578 199764
rect 150438 199744 150578 199753
rect 150494 199736 150578 199744
rect 150578 199718 150630 199724
rect 150438 199679 150494 199688
rect 150682 199696 150710 200124
rect 150774 199764 150802 200124
rect 150866 199918 150894 200124
rect 150958 199918 150986 200124
rect 151050 199918 151078 200124
rect 151142 199918 151170 200124
rect 150854 199912 150906 199918
rect 150854 199854 150906 199860
rect 150946 199912 150998 199918
rect 150946 199854 150998 199860
rect 151038 199912 151090 199918
rect 151038 199854 151090 199860
rect 151130 199912 151182 199918
rect 151130 199854 151182 199860
rect 150992 199776 151044 199782
rect 150774 199736 150848 199764
rect 150682 199668 150756 199696
rect 150268 199600 150342 199628
rect 150440 199640 150492 199646
rect 150164 195356 150216 195362
rect 150164 195298 150216 195304
rect 150268 192438 150296 199600
rect 150440 199582 150492 199588
rect 150532 199640 150584 199646
rect 150532 199582 150584 199588
rect 150452 197130 150480 199582
rect 150440 197124 150492 197130
rect 150440 197066 150492 197072
rect 150544 196858 150572 199582
rect 150624 199436 150676 199442
rect 150624 199378 150676 199384
rect 150532 196852 150584 196858
rect 150532 196794 150584 196800
rect 150348 196784 150400 196790
rect 150348 196726 150400 196732
rect 150256 192432 150308 192438
rect 150256 192374 150308 192380
rect 149796 191412 149848 191418
rect 149796 191354 149848 191360
rect 149704 145852 149756 145858
rect 149704 145794 149756 145800
rect 150360 145654 150388 196726
rect 150636 196704 150664 199378
rect 150544 196676 150664 196704
rect 150544 192506 150572 196676
rect 150728 196586 150756 199668
rect 150820 198626 150848 199736
rect 151234 199764 151262 200124
rect 151326 199918 151354 200124
rect 151418 199918 151446 200124
rect 151510 199923 151538 200124
rect 151314 199912 151366 199918
rect 151314 199854 151366 199860
rect 151406 199912 151458 199918
rect 151406 199854 151458 199860
rect 151496 199914 151552 199923
rect 151602 199918 151630 200124
rect 151694 199918 151722 200124
rect 151496 199849 151552 199858
rect 151590 199912 151642 199918
rect 151590 199854 151642 199860
rect 151682 199912 151734 199918
rect 151682 199854 151734 199860
rect 150992 199718 151044 199724
rect 151188 199736 151262 199764
rect 151360 199776 151412 199782
rect 150900 199572 150952 199578
rect 150900 199514 150952 199520
rect 150808 198620 150860 198626
rect 150808 198562 150860 198568
rect 150912 198121 150940 199514
rect 150898 198112 150954 198121
rect 150898 198047 150954 198056
rect 150808 196852 150860 196858
rect 150808 196794 150860 196800
rect 150716 196580 150768 196586
rect 150716 196522 150768 196528
rect 150820 196466 150848 196794
rect 150636 196438 150848 196466
rect 150532 192500 150584 192506
rect 150532 192442 150584 192448
rect 150348 145648 150400 145654
rect 150348 145590 150400 145596
rect 150532 144424 150584 144430
rect 150532 144366 150584 144372
rect 149978 142896 150034 142905
rect 149978 142831 150034 142840
rect 149612 141568 149664 141574
rect 149612 141510 149664 141516
rect 149520 140752 149572 140758
rect 149520 140694 149572 140700
rect 149532 139890 149560 140694
rect 149992 139890 150020 142831
rect 150544 139890 150572 144366
rect 150636 142866 150664 196438
rect 150716 196376 150768 196382
rect 150716 196318 150768 196324
rect 150728 145722 150756 196318
rect 151004 180794 151032 199718
rect 151084 199708 151136 199714
rect 151084 199650 151136 199656
rect 151096 199442 151124 199650
rect 151084 199436 151136 199442
rect 151084 199378 151136 199384
rect 151084 198348 151136 198354
rect 151084 198290 151136 198296
rect 151096 190330 151124 198290
rect 151188 197334 151216 199736
rect 151544 199776 151596 199782
rect 151360 199718 151412 199724
rect 151450 199744 151506 199753
rect 151268 199436 151320 199442
rect 151268 199378 151320 199384
rect 151176 197328 151228 197334
rect 151176 197270 151228 197276
rect 151280 197198 151308 199378
rect 151268 197192 151320 197198
rect 151268 197134 151320 197140
rect 151176 197124 151228 197130
rect 151176 197066 151228 197072
rect 151084 190324 151136 190330
rect 151084 190266 151136 190272
rect 150820 180766 151032 180794
rect 150820 148617 150848 180766
rect 150806 148608 150862 148617
rect 150806 148543 150862 148552
rect 150716 145716 150768 145722
rect 150716 145658 150768 145664
rect 151082 144664 151138 144673
rect 151082 144599 151138 144608
rect 150624 142860 150676 142866
rect 150624 142802 150676 142808
rect 151096 139890 151124 144599
rect 151188 140282 151216 197066
rect 151372 193214 151400 199718
rect 151786 199764 151814 200124
rect 151878 199918 151906 200124
rect 151866 199912 151918 199918
rect 151866 199854 151918 199860
rect 151786 199736 151860 199764
rect 151544 199718 151596 199724
rect 151450 199679 151506 199688
rect 151464 199442 151492 199679
rect 151452 199436 151504 199442
rect 151452 199378 151504 199384
rect 151556 196382 151584 199718
rect 151636 199708 151688 199714
rect 151636 199650 151688 199656
rect 151544 196376 151596 196382
rect 151544 196318 151596 196324
rect 151280 193186 151400 193214
rect 151176 140276 151228 140282
rect 151176 140218 151228 140224
rect 151280 140146 151308 193186
rect 151648 189553 151676 199650
rect 151728 199368 151780 199374
rect 151728 199310 151780 199316
rect 151740 195401 151768 199310
rect 151832 199238 151860 199736
rect 151970 199730 151998 200124
rect 152062 199918 152090 200124
rect 152154 199918 152182 200124
rect 152246 199918 152274 200124
rect 152050 199912 152102 199918
rect 152050 199854 152102 199860
rect 152142 199912 152194 199918
rect 152142 199854 152194 199860
rect 152234 199912 152286 199918
rect 152234 199854 152286 199860
rect 151970 199702 152044 199730
rect 151912 199572 151964 199578
rect 151912 199514 151964 199520
rect 151820 199232 151872 199238
rect 151820 199174 151872 199180
rect 151818 197024 151874 197033
rect 151818 196959 151874 196968
rect 151726 195392 151782 195401
rect 151726 195327 151782 195336
rect 151832 193934 151860 196959
rect 151924 195498 151952 199514
rect 151912 195492 151964 195498
rect 151912 195434 151964 195440
rect 151912 194744 151964 194750
rect 151912 194686 151964 194692
rect 151820 193928 151872 193934
rect 151820 193870 151872 193876
rect 151634 189544 151690 189553
rect 151634 189479 151690 189488
rect 151820 145784 151872 145790
rect 151820 145726 151872 145732
rect 151832 140758 151860 145726
rect 151924 144401 151952 194686
rect 151910 144392 151966 144401
rect 151910 144327 151966 144336
rect 152016 144129 152044 199702
rect 152096 199708 152148 199714
rect 152096 199650 152148 199656
rect 152188 199708 152240 199714
rect 152338 199696 152366 200124
rect 152430 199918 152458 200124
rect 152522 199918 152550 200124
rect 152614 199923 152642 200124
rect 152418 199912 152470 199918
rect 152418 199854 152470 199860
rect 152510 199912 152562 199918
rect 152510 199854 152562 199860
rect 152600 199914 152656 199923
rect 152706 199918 152734 200124
rect 152798 199918 152826 200124
rect 152890 199918 152918 200124
rect 152600 199849 152656 199858
rect 152694 199912 152746 199918
rect 152694 199854 152746 199860
rect 152786 199912 152838 199918
rect 152786 199854 152838 199860
rect 152878 199912 152930 199918
rect 152878 199854 152930 199860
rect 152464 199776 152516 199782
rect 152464 199718 152516 199724
rect 152556 199776 152608 199782
rect 152556 199718 152608 199724
rect 152648 199776 152700 199782
rect 152648 199718 152700 199724
rect 152740 199776 152792 199782
rect 152740 199718 152792 199724
rect 152338 199668 152412 199696
rect 152188 199650 152240 199656
rect 152108 195906 152136 199650
rect 152200 196466 152228 199650
rect 152384 198801 152412 199668
rect 152370 198792 152426 198801
rect 152370 198727 152426 198736
rect 152200 196438 152320 196466
rect 152096 195900 152148 195906
rect 152096 195842 152148 195848
rect 152096 195492 152148 195498
rect 152096 195434 152148 195440
rect 152108 148442 152136 195434
rect 152188 195084 152240 195090
rect 152188 195026 152240 195032
rect 152200 148646 152228 195026
rect 152292 158030 152320 196438
rect 152372 195900 152424 195906
rect 152372 195842 152424 195848
rect 152384 186998 152412 195842
rect 152372 186992 152424 186998
rect 152372 186934 152424 186940
rect 152372 158296 152424 158302
rect 152372 158238 152424 158244
rect 152280 158024 152332 158030
rect 152280 157966 152332 157972
rect 152188 148640 152240 148646
rect 152188 148582 152240 148588
rect 152096 148436 152148 148442
rect 152096 148378 152148 148384
rect 152002 144120 152058 144129
rect 152002 144055 152058 144064
rect 151820 140752 151872 140758
rect 151820 140694 151872 140700
rect 151268 140140 151320 140146
rect 151268 140082 151320 140088
rect 152384 139890 152412 158238
rect 152476 144265 152504 199718
rect 152568 195265 152596 199718
rect 152554 195256 152610 195265
rect 152554 195191 152610 195200
rect 152660 194750 152688 199718
rect 152752 195294 152780 199718
rect 152832 199708 152884 199714
rect 152982 199696 153010 200124
rect 153074 199923 153102 200124
rect 153060 199914 153116 199923
rect 153166 199918 153194 200124
rect 153258 199918 153286 200124
rect 153060 199849 153116 199858
rect 153154 199912 153206 199918
rect 153154 199854 153206 199860
rect 153246 199912 153298 199918
rect 153246 199854 153298 199860
rect 153350 199764 153378 200124
rect 153442 199923 153470 200124
rect 153428 199914 153484 199923
rect 153534 199918 153562 200124
rect 153428 199849 153484 199858
rect 153522 199912 153574 199918
rect 153522 199854 153574 199860
rect 153350 199736 153424 199764
rect 152832 199650 152884 199656
rect 152936 199668 153010 199696
rect 152740 195288 152792 195294
rect 152740 195230 152792 195236
rect 152648 194744 152700 194750
rect 152648 194686 152700 194692
rect 152844 186969 152872 199650
rect 152936 195090 152964 199668
rect 153108 199640 153160 199646
rect 153108 199582 153160 199588
rect 153292 199640 153344 199646
rect 153292 199582 153344 199588
rect 153120 195537 153148 199582
rect 153200 199572 153252 199578
rect 153200 199514 153252 199520
rect 153212 199374 153240 199514
rect 153200 199368 153252 199374
rect 153200 199310 153252 199316
rect 153200 196852 153252 196858
rect 153200 196794 153252 196800
rect 153106 195528 153162 195537
rect 153106 195463 153162 195472
rect 152924 195084 152976 195090
rect 152924 195026 152976 195032
rect 153212 193050 153240 196794
rect 153200 193044 153252 193050
rect 153200 192986 153252 192992
rect 153304 192982 153332 199582
rect 153396 196722 153424 199736
rect 153626 199696 153654 200124
rect 153580 199668 153654 199696
rect 153476 199640 153528 199646
rect 153476 199582 153528 199588
rect 153384 196716 153436 196722
rect 153384 196658 153436 196664
rect 153488 195922 153516 199582
rect 153396 195894 153516 195922
rect 153292 192976 153344 192982
rect 153292 192918 153344 192924
rect 153292 191548 153344 191554
rect 153292 191490 153344 191496
rect 152830 186960 152886 186969
rect 152830 186895 152886 186904
rect 153304 145761 153332 191490
rect 153396 148481 153424 195894
rect 153476 192976 153528 192982
rect 153476 192918 153528 192924
rect 153488 148850 153516 192918
rect 153580 192817 153608 199668
rect 153718 199594 153746 200124
rect 153810 199764 153838 200124
rect 153902 199923 153930 200124
rect 153888 199914 153944 199923
rect 153888 199849 153944 199858
rect 153994 199764 154022 200124
rect 154086 199918 154114 200124
rect 154178 199918 154206 200124
rect 154270 199918 154298 200124
rect 154362 199923 154390 200124
rect 154074 199912 154126 199918
rect 154074 199854 154126 199860
rect 154166 199912 154218 199918
rect 154166 199854 154218 199860
rect 154258 199912 154310 199918
rect 154258 199854 154310 199860
rect 154348 199914 154404 199923
rect 154454 199918 154482 200124
rect 154546 199918 154574 200124
rect 154348 199849 154404 199858
rect 154442 199912 154494 199918
rect 154442 199854 154494 199860
rect 154534 199912 154586 199918
rect 154534 199854 154586 199860
rect 153810 199736 153884 199764
rect 153718 199566 153792 199594
rect 153660 199504 153712 199510
rect 153660 199446 153712 199452
rect 153672 196858 153700 199446
rect 153660 196852 153712 196858
rect 153660 196794 153712 196800
rect 153660 196648 153712 196654
rect 153660 196590 153712 196596
rect 153566 192808 153622 192817
rect 153566 192743 153622 192752
rect 153568 151088 153620 151094
rect 153568 151030 153620 151036
rect 153476 148844 153528 148850
rect 153476 148786 153528 148792
rect 153382 148472 153438 148481
rect 153382 148407 153438 148416
rect 153290 145752 153346 145761
rect 153290 145687 153346 145696
rect 152462 144256 152518 144265
rect 152462 144191 152518 144200
rect 152646 144120 152702 144129
rect 152646 144055 152702 144064
rect 152660 139890 152688 144055
rect 152740 140752 152792 140758
rect 152740 140694 152792 140700
rect 149532 139862 149776 139890
rect 149992 139862 150328 139890
rect 150544 139862 150880 139890
rect 151096 139862 151432 139890
rect 151984 139862 152412 139890
rect 152536 139862 152688 139890
rect 152752 139890 152780 140694
rect 153580 139890 153608 151030
rect 153672 141438 153700 196590
rect 153764 187377 153792 199566
rect 153856 198694 153884 199736
rect 153948 199736 154022 199764
rect 154212 199776 154264 199782
rect 154118 199744 154174 199753
rect 153948 199578 153976 199736
rect 154396 199776 154448 199782
rect 154212 199718 154264 199724
rect 154302 199744 154358 199753
rect 154118 199679 154174 199688
rect 154028 199640 154080 199646
rect 154028 199582 154080 199588
rect 153936 199572 153988 199578
rect 153936 199514 153988 199520
rect 153936 199368 153988 199374
rect 153936 199310 153988 199316
rect 153844 198688 153896 198694
rect 153844 198630 153896 198636
rect 153948 196625 153976 199310
rect 154040 196790 154068 199582
rect 154028 196784 154080 196790
rect 154028 196726 154080 196732
rect 153934 196616 153990 196625
rect 153934 196551 153990 196560
rect 154028 195968 154080 195974
rect 154028 195910 154080 195916
rect 153750 187368 153806 187377
rect 153750 187303 153806 187312
rect 153660 141432 153712 141438
rect 153660 141374 153712 141380
rect 154040 140185 154068 195910
rect 154132 192953 154160 199679
rect 154224 199510 154252 199718
rect 154396 199718 154448 199724
rect 154488 199776 154540 199782
rect 154638 199764 154666 200124
rect 154730 199918 154758 200124
rect 154822 199923 154850 200124
rect 154718 199912 154770 199918
rect 154718 199854 154770 199860
rect 154808 199914 154864 199923
rect 154914 199918 154942 200124
rect 155006 199918 155034 200124
rect 155098 199923 155126 200124
rect 154808 199849 154864 199858
rect 154902 199912 154954 199918
rect 154902 199854 154954 199860
rect 154994 199912 155046 199918
rect 154994 199854 155046 199860
rect 155084 199914 155140 199923
rect 155190 199918 155218 200124
rect 155084 199849 155140 199858
rect 155178 199912 155230 199918
rect 155178 199854 155230 199860
rect 154488 199718 154540 199724
rect 154592 199736 154666 199764
rect 154856 199776 154908 199782
rect 154762 199744 154818 199753
rect 154302 199679 154358 199688
rect 154212 199504 154264 199510
rect 154212 199446 154264 199452
rect 154118 192944 154174 192953
rect 154118 192879 154174 192888
rect 154316 191554 154344 199679
rect 154408 193361 154436 199718
rect 154500 199034 154528 199718
rect 154592 199646 154620 199736
rect 154856 199718 154908 199724
rect 154948 199776 155000 199782
rect 154948 199718 155000 199724
rect 155132 199776 155184 199782
rect 155282 199764 155310 200124
rect 155374 199918 155402 200124
rect 155362 199912 155414 199918
rect 155362 199854 155414 199860
rect 155132 199718 155184 199724
rect 155236 199736 155310 199764
rect 154762 199679 154818 199688
rect 154580 199640 154632 199646
rect 154580 199582 154632 199588
rect 154672 199640 154724 199646
rect 154672 199582 154724 199588
rect 154488 199028 154540 199034
rect 154488 198970 154540 198976
rect 154684 195974 154712 199582
rect 154776 199102 154804 199679
rect 154764 199096 154816 199102
rect 154764 199038 154816 199044
rect 154868 198558 154896 199718
rect 154856 198552 154908 198558
rect 154856 198494 154908 198500
rect 154960 198354 154988 199718
rect 155040 199708 155092 199714
rect 155040 199650 155092 199656
rect 155052 198762 155080 199650
rect 155040 198756 155092 198762
rect 155040 198698 155092 198704
rect 154948 198348 155000 198354
rect 154948 198290 155000 198296
rect 154856 197124 154908 197130
rect 154856 197066 154908 197072
rect 154672 195968 154724 195974
rect 154672 195910 154724 195916
rect 154764 195968 154816 195974
rect 154764 195910 154816 195916
rect 154672 195764 154724 195770
rect 154672 195706 154724 195712
rect 154394 193352 154450 193361
rect 154394 193287 154450 193296
rect 154304 191548 154356 191554
rect 154304 191490 154356 191496
rect 154578 144392 154634 144401
rect 154578 144327 154634 144336
rect 154302 144256 154358 144265
rect 154302 144191 154358 144200
rect 154026 140176 154082 140185
rect 154026 140111 154082 140120
rect 154316 139890 154344 144191
rect 152752 139862 153088 139890
rect 153580 139862 153640 139890
rect 154192 139862 154344 139890
rect 154592 139890 154620 144327
rect 154684 141438 154712 195706
rect 154776 141574 154804 195910
rect 154868 194041 154896 197066
rect 154854 194032 154910 194041
rect 154854 193967 154910 193976
rect 155144 193214 155172 199718
rect 154868 193186 155172 193214
rect 154868 143002 154896 193186
rect 155236 192506 155264 199736
rect 155466 199730 155494 200124
rect 155420 199702 155494 199730
rect 155316 199640 155368 199646
rect 155316 199582 155368 199588
rect 155328 197198 155356 199582
rect 155316 197192 155368 197198
rect 155316 197134 155368 197140
rect 155224 192500 155276 192506
rect 155224 192442 155276 192448
rect 155420 192386 155448 199702
rect 155558 199594 155586 200124
rect 154960 192358 155448 192386
rect 155512 199566 155586 199594
rect 155650 199594 155678 200124
rect 155742 199696 155770 200124
rect 155834 199764 155862 200124
rect 155926 199918 155954 200124
rect 156018 199918 156046 200124
rect 156110 199923 156138 200124
rect 155914 199912 155966 199918
rect 155914 199854 155966 199860
rect 156006 199912 156058 199918
rect 156006 199854 156058 199860
rect 156096 199914 156152 199923
rect 156202 199918 156230 200124
rect 156096 199849 156152 199858
rect 156190 199912 156242 199918
rect 156190 199854 156242 199860
rect 155960 199776 156012 199782
rect 155834 199736 155908 199764
rect 155742 199668 155816 199696
rect 155650 199566 155724 199594
rect 154960 152522 154988 192358
rect 155512 190466 155540 199566
rect 155592 199504 155644 199510
rect 155592 199446 155644 199452
rect 155604 199345 155632 199446
rect 155590 199336 155646 199345
rect 155590 199271 155646 199280
rect 155696 198694 155724 199566
rect 155684 198688 155736 198694
rect 155684 198630 155736 198636
rect 155500 190460 155552 190466
rect 155500 190402 155552 190408
rect 154948 152516 155000 152522
rect 154948 152458 155000 152464
rect 154948 151156 155000 151162
rect 154948 151098 155000 151104
rect 154856 142996 154908 143002
rect 154856 142938 154908 142944
rect 154764 141568 154816 141574
rect 154764 141510 154816 141516
rect 154672 141432 154724 141438
rect 154672 141374 154724 141380
rect 154960 139890 154988 151098
rect 155684 144492 155736 144498
rect 155684 144434 155736 144440
rect 155696 139890 155724 144434
rect 155788 140146 155816 199668
rect 155880 195974 155908 199736
rect 156294 199764 156322 200124
rect 155960 199718 156012 199724
rect 156050 199744 156106 199753
rect 155868 195968 155920 195974
rect 155868 195910 155920 195916
rect 155972 195770 156000 199718
rect 156050 199679 156106 199688
rect 156248 199736 156322 199764
rect 156386 199764 156414 200124
rect 156478 199918 156506 200124
rect 156466 199912 156518 199918
rect 156466 199854 156518 199860
rect 156386 199736 156460 199764
rect 155960 195764 156012 195770
rect 155960 195706 156012 195712
rect 156064 195650 156092 199679
rect 156248 195922 156276 199736
rect 156326 199608 156382 199617
rect 156326 199543 156382 199552
rect 156340 199170 156368 199543
rect 156328 199164 156380 199170
rect 156328 199106 156380 199112
rect 156432 197130 156460 199736
rect 156570 199730 156598 200124
rect 156662 199764 156690 200124
rect 156754 199918 156782 200124
rect 156846 199918 156874 200124
rect 156938 199918 156966 200124
rect 157030 199918 157058 200124
rect 157122 199923 157150 200124
rect 156742 199912 156794 199918
rect 156742 199854 156794 199860
rect 156834 199912 156886 199918
rect 156834 199854 156886 199860
rect 156926 199912 156978 199918
rect 156926 199854 156978 199860
rect 157018 199912 157070 199918
rect 157018 199854 157070 199860
rect 157108 199914 157164 199923
rect 157214 199918 157242 200124
rect 157306 199918 157334 200124
rect 157108 199849 157164 199858
rect 157202 199912 157254 199918
rect 157202 199854 157254 199860
rect 157294 199912 157346 199918
rect 157294 199854 157346 199860
rect 156788 199776 156840 199782
rect 156662 199736 156736 199764
rect 156524 199702 156598 199730
rect 156420 197124 156472 197130
rect 156420 197066 156472 197072
rect 155880 195622 156092 195650
rect 156156 195894 156276 195922
rect 155880 144430 155908 195622
rect 156052 195356 156104 195362
rect 156052 195298 156104 195304
rect 155868 144424 155920 144430
rect 155868 144366 155920 144372
rect 156064 143070 156092 195298
rect 156156 147082 156184 195894
rect 156236 195764 156288 195770
rect 156236 195706 156288 195712
rect 156248 153134 156276 195706
rect 156524 195362 156552 199702
rect 156604 199640 156656 199646
rect 156604 199582 156656 199588
rect 156616 199238 156644 199582
rect 156604 199232 156656 199238
rect 156604 199174 156656 199180
rect 156512 195356 156564 195362
rect 156512 195298 156564 195304
rect 156708 195242 156736 199736
rect 156788 199718 156840 199724
rect 156880 199776 156932 199782
rect 157398 199764 157426 200124
rect 157490 199918 157518 200124
rect 157582 199918 157610 200124
rect 157674 199918 157702 200124
rect 157766 199923 157794 200124
rect 157478 199912 157530 199918
rect 157478 199854 157530 199860
rect 157570 199912 157622 199918
rect 157570 199854 157622 199860
rect 157662 199912 157714 199918
rect 157662 199854 157714 199860
rect 157752 199914 157808 199923
rect 157858 199918 157886 200124
rect 157950 199918 157978 200124
rect 158042 199923 158070 200124
rect 157752 199849 157808 199858
rect 157846 199912 157898 199918
rect 157846 199854 157898 199860
rect 157938 199912 157990 199918
rect 157938 199854 157990 199860
rect 158028 199914 158084 199923
rect 158028 199849 158084 199858
rect 157892 199776 157944 199782
rect 157016 199744 157072 199753
rect 156932 199724 157016 199730
rect 156880 199718 157016 199724
rect 156432 195214 156736 195242
rect 156328 194880 156380 194886
rect 156328 194822 156380 194828
rect 156340 187134 156368 194822
rect 156432 189786 156460 195214
rect 156512 193384 156564 193390
rect 156512 193326 156564 193332
rect 156524 189854 156552 193326
rect 156800 191834 156828 199718
rect 156892 199702 157016 199718
rect 157398 199736 157472 199764
rect 157016 199679 157072 199688
rect 156880 199640 156932 199646
rect 156880 199582 156932 199588
rect 156972 199640 157024 199646
rect 157248 199640 157300 199646
rect 156972 199582 157024 199588
rect 157062 199608 157118 199617
rect 156892 198121 156920 199582
rect 156878 198112 156934 198121
rect 156878 198047 156934 198056
rect 156984 194886 157012 199582
rect 157248 199582 157300 199588
rect 157062 199543 157118 199552
rect 157156 199572 157208 199578
rect 157076 195770 157104 199543
rect 157156 199514 157208 199520
rect 157168 198830 157196 199514
rect 157156 198824 157208 198830
rect 157156 198766 157208 198772
rect 157064 195764 157116 195770
rect 157064 195706 157116 195712
rect 156972 194880 157024 194886
rect 156972 194822 157024 194828
rect 157260 193390 157288 199582
rect 157340 198824 157392 198830
rect 157340 198766 157392 198772
rect 157352 196110 157380 198766
rect 157340 196104 157392 196110
rect 157340 196046 157392 196052
rect 157340 195968 157392 195974
rect 157340 195910 157392 195916
rect 157248 193384 157300 193390
rect 157248 193326 157300 193332
rect 157352 191834 157380 195910
rect 156708 191806 156828 191834
rect 157260 191806 157380 191834
rect 156708 190454 156736 191806
rect 156708 190426 157012 190454
rect 156512 189848 156564 189854
rect 156512 189790 156564 189796
rect 156420 189780 156472 189786
rect 156420 189722 156472 189728
rect 156328 187128 156380 187134
rect 156328 187070 156380 187076
rect 156236 153128 156288 153134
rect 156236 153070 156288 153076
rect 156144 147076 156196 147082
rect 156144 147018 156196 147024
rect 156696 144628 156748 144634
rect 156696 144570 156748 144576
rect 156052 143064 156104 143070
rect 156052 143006 156104 143012
rect 155776 140140 155828 140146
rect 155776 140082 155828 140088
rect 156708 139890 156736 144570
rect 156984 141710 157012 190426
rect 157260 145722 157288 191806
rect 157444 152454 157472 199736
rect 158134 199764 158162 200124
rect 158226 199918 158254 200124
rect 158318 199923 158346 200124
rect 158214 199912 158266 199918
rect 158214 199854 158266 199860
rect 158304 199914 158360 199923
rect 158304 199849 158360 199858
rect 157892 199718 157944 199724
rect 157982 199744 158038 199753
rect 157524 199708 157576 199714
rect 157524 199650 157576 199656
rect 157616 199708 157668 199714
rect 157616 199650 157668 199656
rect 157536 195974 157564 199650
rect 157524 195968 157576 195974
rect 157524 195910 157576 195916
rect 157524 195832 157576 195838
rect 157524 195774 157576 195780
rect 157536 152726 157564 195774
rect 157628 153066 157656 199650
rect 157708 199640 157760 199646
rect 157708 199582 157760 199588
rect 157798 199608 157854 199617
rect 157720 196722 157748 199582
rect 157798 199543 157854 199552
rect 157708 196716 157760 196722
rect 157708 196658 157760 196664
rect 157812 196246 157840 199543
rect 157904 196518 157932 199718
rect 157982 199679 158038 199688
rect 158088 199736 158162 199764
rect 158260 199776 158312 199782
rect 157892 196512 157944 196518
rect 157892 196454 157944 196460
rect 157996 196330 158024 199679
rect 158088 197130 158116 199736
rect 158410 199753 158438 200124
rect 158502 199918 158530 200124
rect 158594 199918 158622 200124
rect 158686 199923 158714 200124
rect 158490 199912 158542 199918
rect 158490 199854 158542 199860
rect 158582 199912 158634 199918
rect 158582 199854 158634 199860
rect 158672 199914 158728 199923
rect 158672 199849 158728 199858
rect 158628 199776 158680 199782
rect 158260 199718 158312 199724
rect 158396 199744 158452 199753
rect 158076 197124 158128 197130
rect 158076 197066 158128 197072
rect 157904 196302 158024 196330
rect 157800 196240 157852 196246
rect 157800 196182 157852 196188
rect 157798 196072 157854 196081
rect 157798 196007 157854 196016
rect 157708 193180 157760 193186
rect 157708 193122 157760 193128
rect 157720 155514 157748 193122
rect 157812 189990 157840 196007
rect 157904 190126 157932 196302
rect 157984 196240 158036 196246
rect 157984 196182 158036 196188
rect 157892 190120 157944 190126
rect 157892 190062 157944 190068
rect 157800 189984 157852 189990
rect 157800 189926 157852 189932
rect 157996 189922 158024 196182
rect 158272 193186 158300 199718
rect 158778 199730 158806 200124
rect 158870 199764 158898 200124
rect 158962 199918 158990 200124
rect 159054 199918 159082 200124
rect 159146 199918 159174 200124
rect 159238 199918 159266 200124
rect 159330 199923 159358 200124
rect 158950 199912 159002 199918
rect 158950 199854 159002 199860
rect 159042 199912 159094 199918
rect 159042 199854 159094 199860
rect 159134 199912 159186 199918
rect 159134 199854 159186 199860
rect 159226 199912 159278 199918
rect 159226 199854 159278 199860
rect 159316 199914 159372 199923
rect 159316 199849 159372 199858
rect 158996 199776 159048 199782
rect 158870 199736 158944 199764
rect 158628 199718 158680 199724
rect 158396 199679 158452 199688
rect 158444 199640 158496 199646
rect 158444 199582 158496 199588
rect 158456 195838 158484 199582
rect 158536 196716 158588 196722
rect 158536 196658 158588 196664
rect 158444 195832 158496 195838
rect 158444 195774 158496 195780
rect 158260 193180 158312 193186
rect 158260 193122 158312 193128
rect 157984 189916 158036 189922
rect 157984 189858 158036 189864
rect 157708 155508 157760 155514
rect 157708 155450 157760 155456
rect 158548 153202 158576 196658
rect 158640 192545 158668 199718
rect 158732 199702 158806 199730
rect 158732 198150 158760 199702
rect 158810 199608 158866 199617
rect 158810 199543 158866 199552
rect 158720 198144 158772 198150
rect 158720 198086 158772 198092
rect 158824 197878 158852 199543
rect 158812 197872 158864 197878
rect 158812 197814 158864 197820
rect 158720 195492 158772 195498
rect 158720 195434 158772 195440
rect 158626 192536 158682 192545
rect 158626 192471 158682 192480
rect 158536 153196 158588 153202
rect 158536 153138 158588 153144
rect 157616 153060 157668 153066
rect 157616 153002 157668 153008
rect 157524 152720 157576 152726
rect 157524 152662 157576 152668
rect 158732 152590 158760 195434
rect 158916 195378 158944 199736
rect 159272 199776 159324 199782
rect 158996 199718 159048 199724
rect 159086 199744 159142 199753
rect 159008 195945 159036 199718
rect 159422 199764 159450 200124
rect 159514 199918 159542 200124
rect 159606 199918 159634 200124
rect 159502 199912 159554 199918
rect 159502 199854 159554 199860
rect 159594 199912 159646 199918
rect 159594 199854 159646 199860
rect 159548 199776 159600 199782
rect 159422 199736 159496 199764
rect 159272 199718 159324 199724
rect 159086 199679 159142 199688
rect 159180 199708 159232 199714
rect 159100 198393 159128 199679
rect 159180 199650 159232 199656
rect 159086 198384 159142 198393
rect 159086 198319 159142 198328
rect 158994 195936 159050 195945
rect 158994 195871 159050 195880
rect 158916 195350 159036 195378
rect 158904 195288 158956 195294
rect 158904 195230 158956 195236
rect 158812 193996 158864 194002
rect 158812 193938 158864 193944
rect 158824 155582 158852 193938
rect 158916 187066 158944 195230
rect 159008 194070 159036 195350
rect 158996 194064 159048 194070
rect 158996 194006 159048 194012
rect 159192 191834 159220 199650
rect 159284 196926 159312 199718
rect 159364 199640 159416 199646
rect 159364 199582 159416 199588
rect 159376 199306 159404 199582
rect 159364 199300 159416 199306
rect 159364 199242 159416 199248
rect 159272 196920 159324 196926
rect 159272 196862 159324 196868
rect 159468 193225 159496 199736
rect 159698 199764 159726 200124
rect 159790 199918 159818 200124
rect 159882 199918 159910 200124
rect 159778 199912 159830 199918
rect 159778 199854 159830 199860
rect 159870 199912 159922 199918
rect 159870 199854 159922 199860
rect 159974 199850 160002 200124
rect 160066 199923 160094 200124
rect 160052 199914 160108 199923
rect 160158 199918 160186 200124
rect 159962 199844 160014 199850
rect 160052 199849 160108 199858
rect 160146 199912 160198 199918
rect 160146 199854 160198 199860
rect 159962 199786 160014 199792
rect 160250 199764 160278 200124
rect 159548 199718 159600 199724
rect 159652 199736 159726 199764
rect 160204 199736 160278 199764
rect 160342 199764 160370 200124
rect 160434 199923 160462 200124
rect 160420 199914 160476 199923
rect 160420 199849 160476 199858
rect 160342 199736 160416 199764
rect 159560 194002 159588 199718
rect 159548 193996 159600 194002
rect 159548 193938 159600 193944
rect 159454 193216 159510 193225
rect 159454 193151 159510 193160
rect 159008 191806 159220 191834
rect 159008 190058 159036 191806
rect 158996 190052 159048 190058
rect 158996 189994 159048 190000
rect 159652 189718 159680 199736
rect 159824 199708 159876 199714
rect 159824 199650 159876 199656
rect 159732 199572 159784 199578
rect 159732 199514 159784 199520
rect 159744 195566 159772 199514
rect 159732 195560 159784 195566
rect 159732 195502 159784 195508
rect 159836 195498 159864 199650
rect 159916 199640 159968 199646
rect 159916 199582 159968 199588
rect 159824 195492 159876 195498
rect 159824 195434 159876 195440
rect 159928 195294 159956 199582
rect 160008 199572 160060 199578
rect 160008 199514 160060 199520
rect 160020 197985 160048 199514
rect 160100 199504 160152 199510
rect 160100 199446 160152 199452
rect 160112 199073 160140 199446
rect 160098 199064 160154 199073
rect 160098 198999 160154 199008
rect 160006 197976 160062 197985
rect 160006 197911 160062 197920
rect 160204 196704 160232 199736
rect 160284 199640 160336 199646
rect 160284 199582 160336 199588
rect 160296 196994 160324 199582
rect 160284 196988 160336 196994
rect 160284 196930 160336 196936
rect 160282 196888 160338 196897
rect 160282 196823 160338 196832
rect 160020 196676 160232 196704
rect 159916 195288 159968 195294
rect 159916 195230 159968 195236
rect 159640 189712 159692 189718
rect 159640 189654 159692 189660
rect 158904 187060 158956 187066
rect 158904 187002 158956 187008
rect 158812 155576 158864 155582
rect 158812 155518 158864 155524
rect 158720 152584 158772 152590
rect 158720 152526 158772 152532
rect 157432 152448 157484 152454
rect 157432 152390 157484 152396
rect 160020 148510 160048 196676
rect 160192 194948 160244 194954
rect 160192 194890 160244 194896
rect 160204 152998 160232 194890
rect 160192 152992 160244 152998
rect 160192 152934 160244 152940
rect 160296 152658 160324 196823
rect 160388 195362 160416 199736
rect 160526 199696 160554 200124
rect 160618 199918 160646 200124
rect 160710 199918 160738 200124
rect 160802 199918 160830 200124
rect 160606 199912 160658 199918
rect 160606 199854 160658 199860
rect 160698 199912 160750 199918
rect 160698 199854 160750 199860
rect 160790 199912 160842 199918
rect 160790 199854 160842 199860
rect 160744 199776 160796 199782
rect 160744 199718 160796 199724
rect 160526 199668 160692 199696
rect 160468 199572 160520 199578
rect 160468 199514 160520 199520
rect 160376 195356 160428 195362
rect 160376 195298 160428 195304
rect 160480 195242 160508 199514
rect 160388 195214 160508 195242
rect 160388 187338 160416 195214
rect 160468 195152 160520 195158
rect 160468 195094 160520 195100
rect 160480 187406 160508 195094
rect 160664 191834 160692 199668
rect 160756 194954 160784 199718
rect 160894 199696 160922 200124
rect 160986 199918 161014 200124
rect 161078 199923 161106 200124
rect 160974 199912 161026 199918
rect 160974 199854 161026 199860
rect 161064 199914 161120 199923
rect 161170 199918 161198 200124
rect 161064 199849 161120 199858
rect 161158 199912 161210 199918
rect 161262 199889 161290 200124
rect 161158 199854 161210 199860
rect 161248 199880 161304 199889
rect 161248 199815 161304 199824
rect 161020 199776 161072 199782
rect 161020 199718 161072 199724
rect 161112 199776 161164 199782
rect 161112 199718 161164 199724
rect 160848 199668 160922 199696
rect 160848 197169 160876 199668
rect 160928 199572 160980 199578
rect 160928 199514 160980 199520
rect 160940 198801 160968 199514
rect 161032 199442 161060 199718
rect 161020 199436 161072 199442
rect 161020 199378 161072 199384
rect 160926 198792 160982 198801
rect 160926 198727 160982 198736
rect 160834 197160 160890 197169
rect 160834 197095 160890 197104
rect 161124 196897 161152 199718
rect 161354 199696 161382 200124
rect 161446 199918 161474 200124
rect 161434 199912 161486 199918
rect 161434 199854 161486 199860
rect 161538 199764 161566 200124
rect 161630 199918 161658 200124
rect 161722 199918 161750 200124
rect 161618 199912 161670 199918
rect 161618 199854 161670 199860
rect 161710 199912 161762 199918
rect 161710 199854 161762 199860
rect 161664 199776 161716 199782
rect 161538 199753 161612 199764
rect 161538 199744 161626 199753
rect 161538 199736 161570 199744
rect 161308 199668 161382 199696
rect 161814 199764 161842 200124
rect 161664 199718 161716 199724
rect 161768 199736 161842 199764
rect 161570 199679 161626 199688
rect 161204 199640 161256 199646
rect 161204 199582 161256 199588
rect 161110 196888 161166 196897
rect 161110 196823 161166 196832
rect 161112 196784 161164 196790
rect 160926 196752 160982 196761
rect 161112 196726 161164 196732
rect 160926 196687 160982 196696
rect 160744 194948 160796 194954
rect 160744 194890 160796 194896
rect 160940 191834 160968 196687
rect 160664 191806 160876 191834
rect 160940 191806 161060 191834
rect 160848 191350 160876 191806
rect 160836 191344 160888 191350
rect 160836 191286 160888 191292
rect 160468 187400 160520 187406
rect 160468 187342 160520 187348
rect 160376 187332 160428 187338
rect 160376 187274 160428 187280
rect 160284 152652 160336 152658
rect 160284 152594 160336 152600
rect 161032 148850 161060 191806
rect 161124 190454 161152 196726
rect 161216 195430 161244 199582
rect 161204 195424 161256 195430
rect 161204 195366 161256 195372
rect 161308 195158 161336 199668
rect 161480 199640 161532 199646
rect 161480 199582 161532 199588
rect 161388 199572 161440 199578
rect 161388 199514 161440 199520
rect 161400 195838 161428 199514
rect 161492 197062 161520 199582
rect 161572 199572 161624 199578
rect 161572 199514 161624 199520
rect 161480 197056 161532 197062
rect 161480 196998 161532 197004
rect 161480 196716 161532 196722
rect 161480 196658 161532 196664
rect 161388 195832 161440 195838
rect 161388 195774 161440 195780
rect 161296 195152 161348 195158
rect 161296 195094 161348 195100
rect 161492 191834 161520 196658
rect 161584 196602 161612 199514
rect 161676 196790 161704 199718
rect 161664 196784 161716 196790
rect 161664 196726 161716 196732
rect 161584 196574 161704 196602
rect 161570 195936 161626 195945
rect 161570 195871 161626 195880
rect 161400 191806 161520 191834
rect 161124 190426 161336 190454
rect 161020 148844 161072 148850
rect 161020 148786 161072 148792
rect 161308 148782 161336 190426
rect 161296 148776 161348 148782
rect 161296 148718 161348 148724
rect 160008 148504 160060 148510
rect 160008 148446 160060 148452
rect 157340 147212 157392 147218
rect 157340 147154 157392 147160
rect 157248 145716 157300 145722
rect 157248 145658 157300 145664
rect 157246 142896 157302 142905
rect 157246 142831 157302 142840
rect 156972 141704 157024 141710
rect 156972 141646 157024 141652
rect 157260 139890 157288 142831
rect 157352 140758 157380 147154
rect 161400 146946 161428 191806
rect 161388 146940 161440 146946
rect 161388 146882 161440 146888
rect 157616 145852 157668 145858
rect 157616 145794 157668 145800
rect 157432 141636 157484 141642
rect 157432 141578 157484 141584
rect 157340 140752 157392 140758
rect 157340 140694 157392 140700
rect 154592 139862 154744 139890
rect 154960 139862 155296 139890
rect 155696 139862 155848 139890
rect 156400 139862 156736 139890
rect 156952 139862 157288 139890
rect 157444 139754 157472 141578
rect 157628 139890 157656 145794
rect 161584 145790 161612 195871
rect 161676 145926 161704 196574
rect 161768 148986 161796 199736
rect 161906 199696 161934 200124
rect 161998 199764 162026 200124
rect 162090 199918 162118 200124
rect 162078 199912 162130 199918
rect 162182 199889 162210 200124
rect 162274 199918 162302 200124
rect 162262 199912 162314 199918
rect 162078 199854 162130 199860
rect 162168 199880 162224 199889
rect 162262 199854 162314 199860
rect 162168 199815 162224 199824
rect 161998 199736 162072 199764
rect 161906 199668 161980 199696
rect 161848 196784 161900 196790
rect 161848 196726 161900 196732
rect 161860 155854 161888 196726
rect 161952 187474 161980 199668
rect 162044 198529 162072 199736
rect 162214 199744 162270 199753
rect 162214 199679 162270 199688
rect 162366 199696 162394 200124
rect 162458 199764 162486 200124
rect 162550 199918 162578 200124
rect 162642 199918 162670 200124
rect 162734 199923 162762 200124
rect 162538 199912 162590 199918
rect 162538 199854 162590 199860
rect 162630 199912 162682 199918
rect 162630 199854 162682 199860
rect 162720 199914 162776 199923
rect 162826 199918 162854 200124
rect 162720 199849 162776 199858
rect 162814 199912 162866 199918
rect 162814 199854 162866 199860
rect 162458 199736 162532 199764
rect 162228 199084 162256 199679
rect 162366 199668 162440 199696
rect 162306 199608 162362 199617
rect 162306 199543 162362 199552
rect 162136 199056 162256 199084
rect 162030 198520 162086 198529
rect 162030 198455 162086 198464
rect 162136 194002 162164 199056
rect 162320 198830 162348 199543
rect 162308 198824 162360 198830
rect 162308 198766 162360 198772
rect 162412 196790 162440 199668
rect 162400 196784 162452 196790
rect 162400 196726 162452 196732
rect 162306 195664 162362 195673
rect 162306 195599 162308 195608
rect 162360 195599 162362 195608
rect 162308 195570 162360 195576
rect 162124 193996 162176 194002
rect 162124 193938 162176 193944
rect 162504 192574 162532 199736
rect 162582 199744 162638 199753
rect 162918 199730 162946 200124
rect 163010 199918 163038 200124
rect 163102 199918 163130 200124
rect 163194 199923 163222 200124
rect 162998 199912 163050 199918
rect 162998 199854 163050 199860
rect 163090 199912 163142 199918
rect 163090 199854 163142 199860
rect 163180 199914 163236 199923
rect 163180 199849 163236 199858
rect 163286 199764 163314 200124
rect 163378 199918 163406 200124
rect 163366 199912 163418 199918
rect 163366 199854 163418 199860
rect 163470 199764 163498 200124
rect 162582 199679 162638 199688
rect 162676 199708 162728 199714
rect 162596 197810 162624 199679
rect 162676 199650 162728 199656
rect 162780 199702 162946 199730
rect 163134 199744 163190 199753
rect 163044 199708 163096 199714
rect 162584 197804 162636 197810
rect 162584 197746 162636 197752
rect 162492 192568 162544 192574
rect 162492 192510 162544 192516
rect 161940 187468 161992 187474
rect 161940 187410 161992 187416
rect 161848 155848 161900 155854
rect 161848 155790 161900 155796
rect 161756 148980 161808 148986
rect 161756 148922 161808 148928
rect 161664 145920 161716 145926
rect 161664 145862 161716 145868
rect 161572 145784 161624 145790
rect 161572 145726 161624 145732
rect 159456 144560 159508 144566
rect 159456 144502 159508 144508
rect 158260 140752 158312 140758
rect 158260 140694 158312 140700
rect 158272 139890 158300 140694
rect 159468 139890 159496 144502
rect 160008 144356 160060 144362
rect 160008 144298 160060 144304
rect 160020 139890 160048 144298
rect 162214 143168 162270 143177
rect 160560 143132 160612 143138
rect 162214 143103 162270 143112
rect 160560 143074 160612 143080
rect 160572 139890 160600 143074
rect 161110 141400 161166 141409
rect 161110 141335 161166 141344
rect 161124 139890 161152 141335
rect 162228 139890 162256 143103
rect 162688 141545 162716 199650
rect 162780 148918 162808 199702
rect 163134 199679 163190 199688
rect 163240 199736 163314 199764
rect 163424 199736 163498 199764
rect 163044 199650 163096 199656
rect 162860 199640 162912 199646
rect 162860 199582 162912 199588
rect 162952 199640 163004 199646
rect 162952 199582 163004 199588
rect 162872 196897 162900 199582
rect 162858 196888 162914 196897
rect 162858 196823 162914 196832
rect 162964 196722 162992 199582
rect 163056 197266 163084 199650
rect 163044 197260 163096 197266
rect 163044 197202 163096 197208
rect 162952 196716 163004 196722
rect 162952 196658 163004 196664
rect 162952 196104 163004 196110
rect 162952 196046 163004 196052
rect 162964 155786 162992 196046
rect 163148 193214 163176 199679
rect 163056 193186 163176 193214
rect 163056 155922 163084 193186
rect 163136 193112 163188 193118
rect 163136 193054 163188 193060
rect 163148 158098 163176 193054
rect 163240 191146 163268 199736
rect 163320 199504 163372 199510
rect 163320 199446 163372 199452
rect 163332 198937 163360 199446
rect 163318 198928 163374 198937
rect 163318 198863 163374 198872
rect 163424 196110 163452 199736
rect 163562 199696 163590 200124
rect 163654 199918 163682 200124
rect 163642 199912 163694 199918
rect 163642 199854 163694 199860
rect 163746 199764 163774 200124
rect 163838 199918 163866 200124
rect 163930 199918 163958 200124
rect 163826 199912 163878 199918
rect 163826 199854 163878 199860
rect 163918 199912 163970 199918
rect 164022 199889 164050 200124
rect 164114 199918 164142 200124
rect 164206 199918 164234 200124
rect 164102 199912 164154 199918
rect 163918 199854 163970 199860
rect 164008 199880 164064 199889
rect 164102 199854 164154 199860
rect 164194 199912 164246 199918
rect 164194 199854 164246 199860
rect 164008 199815 164064 199824
rect 163872 199776 163924 199782
rect 163746 199736 163820 199764
rect 163562 199668 163636 199696
rect 163504 199572 163556 199578
rect 163504 199514 163556 199520
rect 163516 196858 163544 199514
rect 163608 197402 163636 199668
rect 163688 199640 163740 199646
rect 163792 199617 163820 199736
rect 163872 199718 163924 199724
rect 163964 199776 164016 199782
rect 163964 199718 164016 199724
rect 164146 199744 164202 199753
rect 163688 199582 163740 199588
rect 163778 199608 163834 199617
rect 163596 197396 163648 197402
rect 163596 197338 163648 197344
rect 163700 197033 163728 199582
rect 163778 199543 163834 199552
rect 163780 199504 163832 199510
rect 163780 199446 163832 199452
rect 163686 197024 163742 197033
rect 163686 196959 163742 196968
rect 163504 196852 163556 196858
rect 163504 196794 163556 196800
rect 163688 196512 163740 196518
rect 163688 196454 163740 196460
rect 163412 196104 163464 196110
rect 163412 196046 163464 196052
rect 163228 191140 163280 191146
rect 163228 191082 163280 191088
rect 163700 190454 163728 196454
rect 163792 195809 163820 199446
rect 163884 197538 163912 199718
rect 163872 197532 163924 197538
rect 163872 197474 163924 197480
rect 163872 197192 163924 197198
rect 163872 197134 163924 197140
rect 163778 195800 163834 195809
rect 163778 195735 163834 195744
rect 163700 190426 163820 190454
rect 163136 158092 163188 158098
rect 163136 158034 163188 158040
rect 163044 155916 163096 155922
rect 163044 155858 163096 155864
rect 162952 155780 163004 155786
rect 162952 155722 163004 155728
rect 162952 153944 163004 153950
rect 162952 153886 163004 153892
rect 162768 148912 162820 148918
rect 162768 148854 162820 148860
rect 162766 144528 162822 144537
rect 162766 144463 162822 144472
rect 162674 141536 162730 141545
rect 162674 141471 162730 141480
rect 162780 139890 162808 144463
rect 157628 139862 158056 139890
rect 158272 139862 158608 139890
rect 159160 139862 159496 139890
rect 159712 139862 160048 139890
rect 160264 139862 160600 139890
rect 160816 139862 161152 139890
rect 161920 139862 162256 139890
rect 162472 139862 162808 139890
rect 162964 139890 162992 153886
rect 163792 141506 163820 190426
rect 163884 187270 163912 197134
rect 163976 193118 164004 199718
rect 164056 199708 164108 199714
rect 164298 199730 164326 200124
rect 164390 199918 164418 200124
rect 164482 199918 164510 200124
rect 164378 199912 164430 199918
rect 164378 199854 164430 199860
rect 164470 199912 164522 199918
rect 164470 199854 164522 199860
rect 164146 199679 164202 199688
rect 164252 199702 164326 199730
rect 164424 199776 164476 199782
rect 164574 199764 164602 200124
rect 164666 199918 164694 200124
rect 164758 199923 164786 200124
rect 164654 199912 164706 199918
rect 164654 199854 164706 199860
rect 164744 199914 164800 199923
rect 164744 199849 164800 199858
rect 164424 199718 164476 199724
rect 164528 199736 164602 199764
rect 164056 199650 164108 199656
rect 164068 196790 164096 199650
rect 164056 196784 164108 196790
rect 164056 196726 164108 196732
rect 163964 193112 164016 193118
rect 163964 193054 164016 193060
rect 164160 191834 164188 199679
rect 163976 191806 164188 191834
rect 163872 187264 163924 187270
rect 163872 187206 163924 187212
rect 163976 145897 164004 191806
rect 164252 148714 164280 199702
rect 164436 199617 164464 199718
rect 164422 199608 164478 199617
rect 164422 199543 164478 199552
rect 164424 199436 164476 199442
rect 164424 199378 164476 199384
rect 164436 199238 164464 199378
rect 164424 199232 164476 199238
rect 164424 199174 164476 199180
rect 164528 196704 164556 199736
rect 164850 199696 164878 200124
rect 164942 199918 164970 200124
rect 164930 199912 164982 199918
rect 164930 199854 164982 199860
rect 165034 199764 165062 200124
rect 165126 199918 165154 200124
rect 165114 199912 165166 199918
rect 165114 199854 165166 199860
rect 165218 199764 165246 200124
rect 165310 199923 165338 200124
rect 165296 199914 165352 199923
rect 165296 199849 165352 199858
rect 165402 199764 165430 200124
rect 165494 199923 165522 200124
rect 165480 199914 165536 199923
rect 165586 199918 165614 200124
rect 165678 199918 165706 200124
rect 165770 199918 165798 200124
rect 165480 199849 165536 199858
rect 165574 199912 165626 199918
rect 165574 199854 165626 199860
rect 165666 199912 165718 199918
rect 165666 199854 165718 199860
rect 165758 199912 165810 199918
rect 165862 199889 165890 200124
rect 165758 199854 165810 199860
rect 165848 199880 165904 199889
rect 165848 199815 165904 199824
rect 165034 199736 165108 199764
rect 165218 199736 165292 199764
rect 165356 199753 165430 199764
rect 164850 199668 164924 199696
rect 164700 199640 164752 199646
rect 164700 199582 164752 199588
rect 164608 199300 164660 199306
rect 164608 199242 164660 199248
rect 164620 199209 164648 199242
rect 164606 199200 164662 199209
rect 164606 199135 164662 199144
rect 164436 196676 164556 196704
rect 164332 194812 164384 194818
rect 164332 194754 164384 194760
rect 164344 155718 164372 194754
rect 164332 155712 164384 155718
rect 164332 155654 164384 155660
rect 164436 155174 164464 196676
rect 164516 195968 164568 195974
rect 164516 195910 164568 195916
rect 164528 155242 164556 195910
rect 164712 191834 164740 199582
rect 164792 199572 164844 199578
rect 164792 199514 164844 199520
rect 164804 195974 164832 199514
rect 164792 195968 164844 195974
rect 164792 195910 164844 195916
rect 164896 194818 164924 199668
rect 164976 199640 165028 199646
rect 164976 199582 165028 199588
rect 164884 194812 164936 194818
rect 164884 194754 164936 194760
rect 164988 192438 165016 199582
rect 165080 195498 165108 199736
rect 165158 199608 165214 199617
rect 165158 199543 165214 199552
rect 165172 199374 165200 199543
rect 165160 199368 165212 199374
rect 165160 199310 165212 199316
rect 165160 199232 165212 199238
rect 165160 199174 165212 199180
rect 165172 198626 165200 199174
rect 165160 198620 165212 198626
rect 165160 198562 165212 198568
rect 165068 195492 165120 195498
rect 165068 195434 165120 195440
rect 164976 192432 165028 192438
rect 164976 192374 165028 192380
rect 165264 191834 165292 199736
rect 165342 199744 165430 199753
rect 165398 199736 165430 199744
rect 165804 199776 165856 199782
rect 165804 199718 165856 199724
rect 165342 199679 165398 199688
rect 165712 199708 165764 199714
rect 165712 199650 165764 199656
rect 165344 199640 165396 199646
rect 165344 199582 165396 199588
rect 165356 196518 165384 199582
rect 165620 199572 165672 199578
rect 165620 199514 165672 199520
rect 165528 199436 165580 199442
rect 165528 199378 165580 199384
rect 165436 199368 165488 199374
rect 165436 199310 165488 199316
rect 165448 199238 165476 199310
rect 165436 199232 165488 199238
rect 165436 199174 165488 199180
rect 165344 196512 165396 196518
rect 165344 196454 165396 196460
rect 165540 195974 165568 199378
rect 165632 198966 165660 199514
rect 165620 198960 165672 198966
rect 165620 198902 165672 198908
rect 165724 196722 165752 199650
rect 165816 198898 165844 199718
rect 165954 199696 165982 200124
rect 166046 199918 166074 200124
rect 166138 199918 166166 200124
rect 166230 199918 166258 200124
rect 166034 199912 166086 199918
rect 166034 199854 166086 199860
rect 166126 199912 166178 199918
rect 166126 199854 166178 199860
rect 166218 199912 166270 199918
rect 166218 199854 166270 199860
rect 166218 199776 166270 199782
rect 165908 199668 165982 199696
rect 166092 199724 166218 199730
rect 166322 199764 166350 200124
rect 166414 199918 166442 200124
rect 166506 199918 166534 200124
rect 166402 199912 166454 199918
rect 166402 199854 166454 199860
rect 166494 199912 166546 199918
rect 166494 199854 166546 199860
rect 166598 199764 166626 200124
rect 166690 199918 166718 200124
rect 166678 199912 166730 199918
rect 166678 199854 166730 199860
rect 166782 199764 166810 200124
rect 166874 199889 166902 200124
rect 166860 199880 166916 199889
rect 166860 199815 166916 199824
rect 166966 199764 166994 200124
rect 167058 199918 167086 200124
rect 167150 199918 167178 200124
rect 167046 199912 167098 199918
rect 167046 199854 167098 199860
rect 167138 199912 167190 199918
rect 167138 199854 167190 199860
rect 166322 199736 166396 199764
rect 166092 199718 166270 199724
rect 166092 199702 166258 199718
rect 165908 199617 165936 199668
rect 165894 199608 165950 199617
rect 166092 199594 166120 199702
rect 166368 199594 166396 199736
rect 165894 199543 165950 199552
rect 166000 199566 166120 199594
rect 166276 199566 166396 199594
rect 166552 199736 166626 199764
rect 166736 199736 166810 199764
rect 166920 199736 166994 199764
rect 166448 199572 166500 199578
rect 165804 198892 165856 198898
rect 165804 198834 165856 198840
rect 165712 196716 165764 196722
rect 165712 196658 165764 196664
rect 166000 196602 166028 199566
rect 166080 199504 166132 199510
rect 166080 199446 166132 199452
rect 166092 197606 166120 199446
rect 166080 197600 166132 197606
rect 166080 197542 166132 197548
rect 166276 197418 166304 199566
rect 166448 199514 166500 199520
rect 166356 199504 166408 199510
rect 166356 199446 166408 199452
rect 165620 196580 165672 196586
rect 165620 196522 165672 196528
rect 165816 196574 166028 196602
rect 166092 197390 166304 197418
rect 165528 195968 165580 195974
rect 165528 195910 165580 195916
rect 165528 194540 165580 194546
rect 165528 194482 165580 194488
rect 164620 191806 164740 191834
rect 165172 191806 165292 191834
rect 164620 158166 164648 191806
rect 165172 180794 165200 191806
rect 164712 180766 165200 180794
rect 164712 158234 164740 180766
rect 164792 158704 164844 158710
rect 164792 158646 164844 158652
rect 164700 158228 164752 158234
rect 164700 158170 164752 158176
rect 164608 158160 164660 158166
rect 164608 158102 164660 158108
rect 164516 155236 164568 155242
rect 164516 155178 164568 155184
rect 164424 155168 164476 155174
rect 164424 155110 164476 155116
rect 164240 148708 164292 148714
rect 164240 148650 164292 148656
rect 163962 145888 164018 145897
rect 163962 145823 164018 145832
rect 164146 144664 164202 144673
rect 164146 144599 164202 144608
rect 163870 143032 163926 143041
rect 163870 142967 163926 142976
rect 163780 141500 163832 141506
rect 163780 141442 163832 141448
rect 163884 139890 163912 142967
rect 164160 140162 164188 144599
rect 162964 139862 163024 139890
rect 163576 139862 163912 139890
rect 164114 140134 164188 140162
rect 164114 139876 164142 140134
rect 164804 139890 164832 158646
rect 165540 145994 165568 194482
rect 165632 148442 165660 196522
rect 165712 196036 165764 196042
rect 165712 195978 165764 195984
rect 165724 155310 165752 195978
rect 165816 155378 165844 196574
rect 165896 196512 165948 196518
rect 165896 196454 165948 196460
rect 165908 155446 165936 196454
rect 165986 196344 166042 196353
rect 165986 196279 166042 196288
rect 166000 158574 166028 196279
rect 165988 158568 166040 158574
rect 165988 158510 166040 158516
rect 166092 158370 166120 197390
rect 166368 196874 166396 199446
rect 166460 197674 166488 199514
rect 166448 197668 166500 197674
rect 166448 197610 166500 197616
rect 166368 196846 166488 196874
rect 166356 196716 166408 196722
rect 166356 196658 166408 196664
rect 166172 195968 166224 195974
rect 166172 195910 166224 195916
rect 166184 187542 166212 195910
rect 166368 191214 166396 196658
rect 166460 196586 166488 196846
rect 166448 196580 166500 196586
rect 166448 196522 166500 196528
rect 166552 195226 166580 199736
rect 166632 199640 166684 199646
rect 166632 199582 166684 199588
rect 166540 195220 166592 195226
rect 166540 195162 166592 195168
rect 166644 194954 166672 199582
rect 166736 196042 166764 199736
rect 166816 199640 166868 199646
rect 166814 199608 166816 199617
rect 166868 199608 166870 199617
rect 166814 199543 166870 199552
rect 166816 199368 166868 199374
rect 166816 199310 166868 199316
rect 166828 199209 166856 199310
rect 166814 199200 166870 199209
rect 166814 199135 166870 199144
rect 166920 198734 166948 199736
rect 167000 199640 167052 199646
rect 167242 199628 167270 200124
rect 167334 199918 167362 200124
rect 167322 199912 167374 199918
rect 167322 199854 167374 199860
rect 167426 199764 167454 200124
rect 167000 199582 167052 199588
rect 167196 199600 167270 199628
rect 167380 199736 167454 199764
rect 166828 198706 166948 198734
rect 166724 196036 166776 196042
rect 166724 195978 166776 195984
rect 166632 194948 166684 194954
rect 166632 194890 166684 194896
rect 166828 193186 166856 198706
rect 167012 198665 167040 199582
rect 167092 199572 167144 199578
rect 167092 199514 167144 199520
rect 166998 198656 167054 198665
rect 166998 198591 167054 198600
rect 166816 193180 166868 193186
rect 166816 193122 166868 193128
rect 167104 191350 167132 199514
rect 167196 196722 167224 199600
rect 167276 199504 167328 199510
rect 167276 199446 167328 199452
rect 167184 196716 167236 196722
rect 167184 196658 167236 196664
rect 167288 195945 167316 199446
rect 167274 195936 167330 195945
rect 167274 195871 167330 195880
rect 167380 194546 167408 199736
rect 167518 199696 167546 200124
rect 167472 199668 167546 199696
rect 167610 199696 167638 200124
rect 167702 199764 167730 200124
rect 167794 199918 167822 200124
rect 167886 199918 167914 200124
rect 167782 199912 167834 199918
rect 167782 199854 167834 199860
rect 167874 199912 167926 199918
rect 167978 199889 168006 200124
rect 168070 199918 168098 200124
rect 168058 199912 168110 199918
rect 167874 199854 167926 199860
rect 167964 199880 168020 199889
rect 168058 199854 168110 199860
rect 167964 199815 168020 199824
rect 167702 199736 167776 199764
rect 167610 199668 167684 199696
rect 167368 194540 167420 194546
rect 167368 194482 167420 194488
rect 167472 193118 167500 199668
rect 167552 199572 167604 199578
rect 167552 199514 167604 199520
rect 167564 199073 167592 199514
rect 167550 199064 167606 199073
rect 167550 198999 167606 199008
rect 167460 193112 167512 193118
rect 167460 193054 167512 193060
rect 167092 191344 167144 191350
rect 167092 191286 167144 191292
rect 167184 191276 167236 191282
rect 167184 191218 167236 191224
rect 166356 191208 166408 191214
rect 166356 191150 166408 191156
rect 167092 191004 167144 191010
rect 167092 190946 167144 190952
rect 166172 187536 166224 187542
rect 166172 187478 166224 187484
rect 166080 158364 166132 158370
rect 166080 158306 166132 158312
rect 165896 155440 165948 155446
rect 165896 155382 165948 155388
rect 165804 155372 165856 155378
rect 165804 155314 165856 155320
rect 165712 155304 165764 155310
rect 165712 155246 165764 155252
rect 165712 154012 165764 154018
rect 165712 153954 165764 153960
rect 165724 151814 165752 153954
rect 165724 151786 165936 151814
rect 165620 148436 165672 148442
rect 165620 148378 165672 148384
rect 165528 145988 165580 145994
rect 165528 145930 165580 145936
rect 165804 144696 165856 144702
rect 165804 144638 165856 144644
rect 165528 143200 165580 143206
rect 165528 143142 165580 143148
rect 165540 139890 165568 143142
rect 165816 140162 165844 144638
rect 164680 139862 164832 139890
rect 165232 139862 165568 139890
rect 165770 140134 165844 140162
rect 165770 139876 165798 140134
rect 165908 139890 165936 151786
rect 167104 148617 167132 190946
rect 167196 151201 167224 191218
rect 167656 190942 167684 199668
rect 167748 198665 167776 199736
rect 167918 199744 167974 199753
rect 167828 199708 167880 199714
rect 167918 199679 167974 199688
rect 168012 199708 168064 199714
rect 167828 199650 167880 199656
rect 167734 198656 167790 198665
rect 167734 198591 167790 198600
rect 167840 198150 167868 199650
rect 167932 198734 167960 199679
rect 168162 199696 168190 200124
rect 168254 199923 168282 200124
rect 168240 199914 168296 199923
rect 168240 199849 168296 199858
rect 168012 199650 168064 199656
rect 168116 199668 168190 199696
rect 168024 199510 168052 199650
rect 168012 199504 168064 199510
rect 168012 199446 168064 199452
rect 167932 198706 168052 198734
rect 167828 198144 167880 198150
rect 167828 198086 167880 198092
rect 167736 198008 167788 198014
rect 167736 197950 167788 197956
rect 167748 197826 167776 197950
rect 167748 197798 167960 197826
rect 167828 197056 167880 197062
rect 167828 196998 167880 197004
rect 167840 191078 167868 196998
rect 167828 191072 167880 191078
rect 167828 191014 167880 191020
rect 167644 190936 167696 190942
rect 167644 190878 167696 190884
rect 167276 151224 167328 151230
rect 167182 151192 167238 151201
rect 167276 151166 167328 151172
rect 167182 151127 167238 151136
rect 167090 148608 167146 148617
rect 167090 148543 167146 148552
rect 166998 145752 167054 145761
rect 166998 145687 167054 145696
rect 166816 141772 166868 141778
rect 166816 141714 166868 141720
rect 165908 139862 166336 139890
rect 166828 139754 166856 141714
rect 167012 140758 167040 145687
rect 167000 140752 167052 140758
rect 167000 140694 167052 140700
rect 167288 139890 167316 151166
rect 167932 146062 167960 197798
rect 168024 191282 168052 198706
rect 168012 191276 168064 191282
rect 168012 191218 168064 191224
rect 168012 191072 168064 191078
rect 168012 191014 168064 191020
rect 168024 158438 168052 191014
rect 168116 191010 168144 199668
rect 168346 199628 168374 200124
rect 168438 199764 168466 200124
rect 168530 199918 168558 200124
rect 168622 199923 168650 200124
rect 168518 199912 168570 199918
rect 168518 199854 168570 199860
rect 168608 199914 168664 199923
rect 168714 199918 168742 200124
rect 168608 199849 168664 199858
rect 168702 199912 168754 199918
rect 168702 199854 168754 199860
rect 168564 199776 168616 199782
rect 168438 199736 168512 199764
rect 168194 199608 168250 199617
rect 168194 199543 168250 199552
rect 168300 199600 168374 199628
rect 168104 191004 168156 191010
rect 168104 190946 168156 190952
rect 168208 187202 168236 199543
rect 168300 197334 168328 199600
rect 168380 199436 168432 199442
rect 168380 199378 168432 199384
rect 168392 198626 168420 199378
rect 168380 198620 168432 198626
rect 168380 198562 168432 198568
rect 168288 197328 168340 197334
rect 168288 197270 168340 197276
rect 168380 195152 168432 195158
rect 168380 195094 168432 195100
rect 168288 190936 168340 190942
rect 168288 190878 168340 190884
rect 168196 187196 168248 187202
rect 168196 187138 168248 187144
rect 168012 158432 168064 158438
rect 168012 158374 168064 158380
rect 168300 148646 168328 190878
rect 168288 148640 168340 148646
rect 168288 148582 168340 148588
rect 167920 146056 167972 146062
rect 167920 145998 167972 146004
rect 168392 142934 168420 195094
rect 168484 191834 168512 199736
rect 168656 199776 168708 199782
rect 168564 199718 168616 199724
rect 168654 199744 168656 199753
rect 168806 199764 168834 200124
rect 168898 199923 168926 200124
rect 168884 199914 168940 199923
rect 168990 199918 169018 200124
rect 168884 199849 168940 199858
rect 168978 199912 169030 199918
rect 168978 199854 169030 199860
rect 169082 199764 169110 200124
rect 169174 199923 169202 200124
rect 169160 199914 169216 199923
rect 169266 199918 169294 200124
rect 169358 199918 169386 200124
rect 169450 199923 169478 200124
rect 169160 199849 169216 199858
rect 169254 199912 169306 199918
rect 169254 199854 169306 199860
rect 169346 199912 169398 199918
rect 169346 199854 169398 199860
rect 169436 199914 169492 199923
rect 169436 199849 169492 199858
rect 168708 199744 168710 199753
rect 168806 199736 168880 199764
rect 168576 199594 168604 199718
rect 168654 199679 168710 199688
rect 168576 199566 168696 199594
rect 168564 199504 168616 199510
rect 168564 199446 168616 199452
rect 168576 195974 168604 199446
rect 168668 197062 168696 199566
rect 168852 198014 168880 199736
rect 168930 199744 168986 199753
rect 169082 199736 169156 199764
rect 168930 199679 168986 199688
rect 168840 198008 168892 198014
rect 168840 197950 168892 197956
rect 168746 197704 168802 197713
rect 168746 197639 168802 197648
rect 168760 197198 168788 197639
rect 168748 197192 168800 197198
rect 168748 197134 168800 197140
rect 168656 197056 168708 197062
rect 168656 196998 168708 197004
rect 168564 195968 168616 195974
rect 168564 195910 168616 195916
rect 168944 192817 168972 199679
rect 169128 199646 169156 199736
rect 169542 199730 169570 200124
rect 169634 199764 169662 200124
rect 169726 199918 169754 200124
rect 169714 199912 169766 199918
rect 169714 199854 169766 199860
rect 169634 199736 169708 199764
rect 169496 199702 169570 199730
rect 169116 199640 169168 199646
rect 169116 199582 169168 199588
rect 169300 199572 169352 199578
rect 169300 199514 169352 199520
rect 169392 199572 169444 199578
rect 169392 199514 169444 199520
rect 169024 199504 169076 199510
rect 169024 199446 169076 199452
rect 169116 199504 169168 199510
rect 169116 199446 169168 199452
rect 169036 193214 169064 199446
rect 169128 198937 169156 199446
rect 169114 198928 169170 198937
rect 169114 198863 169170 198872
rect 169206 198656 169262 198665
rect 169206 198591 169262 198600
rect 169036 193186 169156 193214
rect 168930 192808 168986 192817
rect 168930 192743 168986 192752
rect 169128 191834 169156 193186
rect 169220 192982 169248 198591
rect 169208 192976 169260 192982
rect 169208 192918 169260 192924
rect 168484 191806 168604 191834
rect 168576 188426 168604 191806
rect 168852 191806 169156 191834
rect 169312 191834 169340 199514
rect 169404 198665 169432 199514
rect 169390 198656 169446 198665
rect 169390 198591 169446 198600
rect 169392 198416 169444 198422
rect 169392 198358 169444 198364
rect 169404 195158 169432 198358
rect 169392 195152 169444 195158
rect 169392 195094 169444 195100
rect 169496 191834 169524 199702
rect 169576 199640 169628 199646
rect 169576 199582 169628 199588
rect 169588 193866 169616 199582
rect 169576 193860 169628 193866
rect 169576 193802 169628 193808
rect 169312 191806 169432 191834
rect 169496 191806 169616 191834
rect 168852 188578 168880 191806
rect 168668 188550 168880 188578
rect 168564 188420 168616 188426
rect 168564 188362 168616 188368
rect 168472 188148 168524 188154
rect 168472 188090 168524 188096
rect 168484 144838 168512 188090
rect 168668 151298 168696 188550
rect 168748 188420 168800 188426
rect 168748 188362 168800 188368
rect 168760 158506 168788 188362
rect 169404 187105 169432 191806
rect 169390 187096 169446 187105
rect 169390 187031 169446 187040
rect 169588 186314 169616 191806
rect 169680 188154 169708 199736
rect 169818 199730 169846 200124
rect 169772 199702 169846 199730
rect 169772 191834 169800 199702
rect 169910 199628 169938 200124
rect 170002 199918 170030 200124
rect 170094 199923 170122 200124
rect 169990 199912 170042 199918
rect 169990 199854 170042 199860
rect 170080 199914 170136 199923
rect 170080 199849 170136 199858
rect 170186 199764 170214 200124
rect 170140 199736 170214 199764
rect 169864 199600 169938 199628
rect 170036 199640 170088 199646
rect 169864 193214 169892 199600
rect 170036 199582 170088 199588
rect 170048 198490 170076 199582
rect 170036 198484 170088 198490
rect 170036 198426 170088 198432
rect 170036 197600 170088 197606
rect 170036 197542 170088 197548
rect 170048 195838 170076 197542
rect 170036 195832 170088 195838
rect 170036 195774 170088 195780
rect 169864 193186 169984 193214
rect 169956 192914 169984 193186
rect 169944 192908 169996 192914
rect 169944 192850 169996 192856
rect 170140 192778 170168 199736
rect 170278 199560 170306 200124
rect 170370 199764 170398 200124
rect 170462 199918 170490 200124
rect 170554 199923 170582 200124
rect 170450 199912 170502 199918
rect 170450 199854 170502 199860
rect 170540 199914 170596 199923
rect 170646 199918 170674 200124
rect 170540 199849 170596 199858
rect 170634 199912 170686 199918
rect 170634 199854 170686 199860
rect 170496 199776 170548 199782
rect 170370 199736 170444 199764
rect 170232 199532 170306 199560
rect 170232 198286 170260 199532
rect 170416 199458 170444 199736
rect 170496 199718 170548 199724
rect 170588 199776 170640 199782
rect 170738 199764 170766 200124
rect 170830 199918 170858 200124
rect 170818 199912 170870 199918
rect 170818 199854 170870 199860
rect 170588 199718 170640 199724
rect 170692 199736 170766 199764
rect 170324 199430 170444 199458
rect 170220 198280 170272 198286
rect 170220 198222 170272 198228
rect 170128 192772 170180 192778
rect 170128 192714 170180 192720
rect 169772 191806 169892 191834
rect 169760 191072 169812 191078
rect 169760 191014 169812 191020
rect 169668 188148 169720 188154
rect 169668 188090 169720 188096
rect 169588 186286 169708 186314
rect 168748 158500 168800 158506
rect 168748 158442 168800 158448
rect 168840 157956 168892 157962
rect 168840 157898 168892 157904
rect 168656 151292 168708 151298
rect 168656 151234 168708 151240
rect 168472 144832 168524 144838
rect 168472 144774 168524 144780
rect 168380 142928 168432 142934
rect 168380 142870 168432 142876
rect 168748 141840 168800 141846
rect 168748 141782 168800 141788
rect 167644 140752 167696 140758
rect 167644 140694 167696 140700
rect 167656 139890 167684 140694
rect 168760 139890 168788 141782
rect 168852 140758 168880 157898
rect 168932 157888 168984 157894
rect 168932 157830 168984 157836
rect 168840 140752 168892 140758
rect 168840 140694 168892 140700
rect 167288 139862 167440 139890
rect 167656 139862 167992 139890
rect 168544 139862 168788 139890
rect 168944 139890 168972 157830
rect 169680 148578 169708 186286
rect 169668 148572 169720 148578
rect 169668 148514 169720 148520
rect 169772 140758 169800 191014
rect 169864 147286 169892 191806
rect 170324 186314 170352 199430
rect 170508 198734 170536 199718
rect 170416 198706 170536 198734
rect 170416 193050 170444 198706
rect 170496 198144 170548 198150
rect 170496 198086 170548 198092
rect 170508 197470 170536 198086
rect 170496 197464 170548 197470
rect 170496 197406 170548 197412
rect 170404 193044 170456 193050
rect 170404 192986 170456 192992
rect 169956 186286 170352 186314
rect 169956 147393 169984 186286
rect 170600 180794 170628 199718
rect 170692 192710 170720 199736
rect 170922 199696 170950 200124
rect 171014 199923 171042 200124
rect 171000 199914 171056 199923
rect 171000 199849 171056 199858
rect 171106 199764 171134 200124
rect 171198 199923 171226 200124
rect 171184 199914 171240 199923
rect 171290 199918 171318 200124
rect 171382 199918 171410 200124
rect 171474 199918 171502 200124
rect 171184 199849 171240 199858
rect 171278 199912 171330 199918
rect 171278 199854 171330 199860
rect 171370 199912 171422 199918
rect 171370 199854 171422 199860
rect 171462 199912 171514 199918
rect 171462 199854 171514 199860
rect 171566 199764 171594 200124
rect 171658 199923 171686 200124
rect 171644 199914 171700 199923
rect 171644 199849 171700 199858
rect 171750 199764 171778 200124
rect 171106 199736 171180 199764
rect 170876 199668 170950 199696
rect 170772 199640 170824 199646
rect 170772 199582 170824 199588
rect 170784 197878 170812 199582
rect 170772 197872 170824 197878
rect 170772 197814 170824 197820
rect 170680 192704 170732 192710
rect 170680 192646 170732 192652
rect 170876 191078 170904 199668
rect 170954 199608 171010 199617
rect 170954 199543 171010 199552
rect 171048 199572 171100 199578
rect 170968 195945 170996 199543
rect 171048 199514 171100 199520
rect 171060 198422 171088 199514
rect 171048 198416 171100 198422
rect 171048 198358 171100 198364
rect 171152 198121 171180 199736
rect 171520 199736 171594 199764
rect 171704 199736 171778 199764
rect 171842 199764 171870 200124
rect 171934 199918 171962 200124
rect 172026 199918 172054 200124
rect 171922 199912 171974 199918
rect 171922 199854 171974 199860
rect 172014 199912 172066 199918
rect 172014 199854 172066 199860
rect 171842 199736 172008 199764
rect 171416 199640 171468 199646
rect 171416 199582 171468 199588
rect 171324 199572 171376 199578
rect 171324 199514 171376 199520
rect 171138 198112 171194 198121
rect 171138 198047 171194 198056
rect 171048 197804 171100 197810
rect 171048 197746 171100 197752
rect 170954 195936 171010 195945
rect 170954 195871 171010 195880
rect 170864 191072 170916 191078
rect 170864 191014 170916 191020
rect 170048 180766 170628 180794
rect 169942 147384 169998 147393
rect 170048 147354 170076 180766
rect 170128 153876 170180 153882
rect 170128 153818 170180 153824
rect 169942 147319 169998 147328
rect 170036 147348 170088 147354
rect 170036 147290 170088 147296
rect 169852 147280 169904 147286
rect 169852 147222 169904 147228
rect 169300 140752 169352 140758
rect 169300 140694 169352 140700
rect 169760 140752 169812 140758
rect 169760 140694 169812 140700
rect 169312 139890 169340 140694
rect 170140 139890 170168 153818
rect 171060 149054 171088 197746
rect 171138 196480 171194 196489
rect 171138 196415 171194 196424
rect 171152 193089 171180 196415
rect 171232 196036 171284 196042
rect 171232 195978 171284 195984
rect 171138 193080 171194 193089
rect 171138 193015 171194 193024
rect 171140 191072 171192 191078
rect 171140 191014 171192 191020
rect 171048 149048 171100 149054
rect 171048 148990 171100 148996
rect 171152 147014 171180 191014
rect 171244 147529 171272 195978
rect 171336 195242 171364 199514
rect 171428 196042 171456 199582
rect 171416 196036 171468 196042
rect 171416 195978 171468 195984
rect 171336 195214 171456 195242
rect 171324 195152 171376 195158
rect 171324 195094 171376 195100
rect 171336 149870 171364 195094
rect 171428 192681 171456 195214
rect 171520 192846 171548 199736
rect 171704 199560 171732 199736
rect 171876 199640 171928 199646
rect 171876 199582 171928 199588
rect 171704 199532 171824 199560
rect 171690 199472 171746 199481
rect 171690 199407 171746 199416
rect 171704 199209 171732 199407
rect 171690 199200 171746 199209
rect 171690 199135 171746 199144
rect 171796 196704 171824 199532
rect 171888 198150 171916 199582
rect 171876 198144 171928 198150
rect 171876 198086 171928 198092
rect 171704 196676 171824 196704
rect 171600 195764 171652 195770
rect 171600 195706 171652 195712
rect 171612 195634 171640 195706
rect 171600 195628 171652 195634
rect 171600 195570 171652 195576
rect 171600 193928 171652 193934
rect 171600 193870 171652 193876
rect 171508 192840 171560 192846
rect 171508 192782 171560 192788
rect 171414 192672 171470 192681
rect 171414 192607 171470 192616
rect 171416 191276 171468 191282
rect 171416 191218 171468 191224
rect 171324 149864 171376 149870
rect 171324 149806 171376 149812
rect 171428 149734 171456 191218
rect 171612 186314 171640 193870
rect 171704 191078 171732 196676
rect 171782 196072 171838 196081
rect 171782 196007 171838 196016
rect 171796 192370 171824 196007
rect 171980 194177 172008 199736
rect 172118 199696 172146 200124
rect 172210 199923 172238 200124
rect 172196 199914 172252 199923
rect 172302 199918 172330 200124
rect 172394 199923 172422 200124
rect 172196 199849 172252 199858
rect 172290 199912 172342 199918
rect 172290 199854 172342 199860
rect 172380 199914 172436 199923
rect 172486 199918 172514 200124
rect 172380 199849 172436 199858
rect 172474 199912 172526 199918
rect 172474 199854 172526 199860
rect 172426 199744 172482 199753
rect 172118 199668 172192 199696
rect 172426 199679 172482 199688
rect 172060 199572 172112 199578
rect 172060 199514 172112 199520
rect 172072 198257 172100 199514
rect 172058 198248 172114 198257
rect 172058 198183 172114 198192
rect 172060 197532 172112 197538
rect 172060 197474 172112 197480
rect 171966 194168 172022 194177
rect 171966 194103 172022 194112
rect 171968 192568 172020 192574
rect 171968 192510 172020 192516
rect 171784 192364 171836 192370
rect 171784 192306 171836 192312
rect 171692 191072 171744 191078
rect 171692 191014 171744 191020
rect 171980 186314 172008 192510
rect 171612 186286 171732 186314
rect 171508 155644 171560 155650
rect 171508 155586 171560 155592
rect 171416 149728 171468 149734
rect 171416 149670 171468 149676
rect 171230 147520 171286 147529
rect 171230 147455 171286 147464
rect 171140 147008 171192 147014
rect 171140 146950 171192 146956
rect 171048 144764 171100 144770
rect 171048 144706 171100 144712
rect 171060 139890 171088 144706
rect 171416 143336 171468 143342
rect 171416 143278 171468 143284
rect 171428 139890 171456 143278
rect 168944 139862 169096 139890
rect 169312 139862 169648 139890
rect 170140 139862 170200 139890
rect 170752 139862 171088 139890
rect 171304 139862 171456 139890
rect 171520 139890 171548 155586
rect 171704 152425 171732 186286
rect 171796 186286 172008 186314
rect 171690 152416 171746 152425
rect 171690 152351 171746 152360
rect 171796 146033 171824 186286
rect 172072 180794 172100 197474
rect 172164 192642 172192 199668
rect 172244 199640 172296 199646
rect 172244 199582 172296 199588
rect 172336 199640 172388 199646
rect 172336 199582 172388 199588
rect 172256 195158 172284 199582
rect 172244 195152 172296 195158
rect 172244 195094 172296 195100
rect 172152 192636 172204 192642
rect 172152 192578 172204 192584
rect 172348 191834 172376 199582
rect 172440 197577 172468 199679
rect 172578 199594 172606 200124
rect 172670 199764 172698 200124
rect 172762 199918 172790 200124
rect 172854 199918 172882 200124
rect 172750 199912 172802 199918
rect 172750 199854 172802 199860
rect 172842 199912 172894 199918
rect 172946 199889 172974 200124
rect 173038 199918 173066 200124
rect 173130 199918 173158 200124
rect 173026 199912 173078 199918
rect 172842 199854 172894 199860
rect 172932 199880 172988 199889
rect 173026 199854 173078 199860
rect 173118 199912 173170 199918
rect 173118 199854 173170 199860
rect 173222 199850 173250 200124
rect 172932 199815 172988 199824
rect 173210 199844 173262 199850
rect 173210 199786 173262 199792
rect 172980 199776 173032 199782
rect 172670 199753 172744 199764
rect 172670 199744 172758 199753
rect 172670 199736 172702 199744
rect 173032 199736 173112 199764
rect 172980 199718 173032 199724
rect 172702 199679 172758 199688
rect 172796 199708 172848 199714
rect 172796 199650 172848 199656
rect 172578 199566 172744 199594
rect 172426 197568 172482 197577
rect 172426 197503 172482 197512
rect 172256 191806 172376 191834
rect 172256 191282 172284 191806
rect 172244 191276 172296 191282
rect 172244 191218 172296 191224
rect 172612 191072 172664 191078
rect 172612 191014 172664 191020
rect 172520 187604 172572 187610
rect 172520 187546 172572 187552
rect 171888 180766 172100 180794
rect 171888 150346 171916 180766
rect 171968 151360 172020 151366
rect 171968 151302 172020 151308
rect 171876 150340 171928 150346
rect 171876 150282 171928 150288
rect 171782 146024 171838 146033
rect 171782 145959 171838 145968
rect 171980 139890 172008 151302
rect 172532 147150 172560 187546
rect 172624 149705 172652 191014
rect 172716 150074 172744 199566
rect 172704 150068 172756 150074
rect 172704 150010 172756 150016
rect 172808 149841 172836 199650
rect 172888 199640 172940 199646
rect 172888 199582 172940 199588
rect 172978 199608 173034 199617
rect 172900 150210 172928 199582
rect 173084 199578 173112 199736
rect 173314 199730 173342 200124
rect 173406 199782 173434 200124
rect 173498 199850 173526 200124
rect 173590 199923 173618 200124
rect 173576 199914 173632 199923
rect 173682 199918 173710 200124
rect 173774 199923 173802 200124
rect 173486 199844 173538 199850
rect 173576 199849 173632 199858
rect 173670 199912 173722 199918
rect 173670 199854 173722 199860
rect 173760 199914 173816 199923
rect 173866 199918 173894 200124
rect 173760 199849 173816 199858
rect 173854 199912 173906 199918
rect 173854 199854 173906 199860
rect 173486 199786 173538 199792
rect 173268 199702 173342 199730
rect 173394 199776 173446 199782
rect 173958 199764 173986 200124
rect 174050 199918 174078 200124
rect 174142 199923 174170 200124
rect 174038 199912 174090 199918
rect 174038 199854 174090 199860
rect 174128 199914 174184 199923
rect 174128 199849 174184 199858
rect 174084 199776 174136 199782
rect 173958 199753 174032 199764
rect 173958 199744 174046 199753
rect 173958 199736 173990 199744
rect 173394 199718 173446 199724
rect 173624 199708 173676 199714
rect 173164 199640 173216 199646
rect 173164 199582 173216 199588
rect 172978 199543 173034 199552
rect 173072 199572 173124 199578
rect 172992 192574 173020 199543
rect 173072 199514 173124 199520
rect 173176 194410 173204 199582
rect 173268 198422 173296 199702
rect 174234 199764 174262 200124
rect 174326 199923 174354 200124
rect 174312 199914 174368 199923
rect 174312 199849 174368 199858
rect 174084 199718 174136 199724
rect 174188 199736 174262 199764
rect 173990 199679 174046 199688
rect 173624 199650 173676 199656
rect 173348 199640 173400 199646
rect 173348 199582 173400 199588
rect 173532 199640 173584 199646
rect 173532 199582 173584 199588
rect 173256 198416 173308 198422
rect 173256 198358 173308 198364
rect 173164 194404 173216 194410
rect 173164 194346 173216 194352
rect 172980 192568 173032 192574
rect 172980 192510 173032 192516
rect 173360 187610 173388 199582
rect 173544 194449 173572 199582
rect 173530 194440 173586 194449
rect 173530 194375 173586 194384
rect 173636 191078 173664 199650
rect 173900 199640 173952 199646
rect 173806 199608 173862 199617
rect 173900 199582 173952 199588
rect 173806 199543 173862 199552
rect 173714 199200 173770 199209
rect 173714 199135 173770 199144
rect 173624 191072 173676 191078
rect 173624 191014 173676 191020
rect 173728 190398 173756 199135
rect 173820 197538 173848 199543
rect 173808 197532 173860 197538
rect 173808 197474 173860 197480
rect 173808 197396 173860 197402
rect 173808 197338 173860 197344
rect 173716 190392 173768 190398
rect 173716 190334 173768 190340
rect 173348 187604 173400 187610
rect 173348 187546 173400 187552
rect 173820 180794 173848 197338
rect 173912 193905 173940 199582
rect 173992 199572 174044 199578
rect 173992 199514 174044 199520
rect 174004 198626 174032 199514
rect 173992 198620 174044 198626
rect 173992 198562 174044 198568
rect 174096 194138 174124 199718
rect 174084 194132 174136 194138
rect 174084 194074 174136 194080
rect 173898 193896 173954 193905
rect 173898 193831 173954 193840
rect 174188 191834 174216 199736
rect 174418 199730 174446 200124
rect 174510 199918 174538 200124
rect 174498 199912 174550 199918
rect 174498 199854 174550 199860
rect 174602 199764 174630 200124
rect 174694 199923 174722 200124
rect 174680 199914 174736 199923
rect 174786 199918 174814 200124
rect 174680 199849 174736 199858
rect 174774 199912 174826 199918
rect 174774 199854 174826 199860
rect 174878 199764 174906 200124
rect 174372 199702 174446 199730
rect 174556 199736 174630 199764
rect 174832 199736 174906 199764
rect 174268 199572 174320 199578
rect 174268 199514 174320 199520
rect 174280 194324 174308 199514
rect 174372 199209 174400 199702
rect 174450 199608 174506 199617
rect 174450 199543 174452 199552
rect 174504 199543 174506 199552
rect 174452 199514 174504 199520
rect 174556 199458 174584 199736
rect 174728 199708 174780 199714
rect 174728 199650 174780 199656
rect 174634 199608 174690 199617
rect 174634 199543 174690 199552
rect 174464 199430 174584 199458
rect 174358 199200 174414 199209
rect 174358 199135 174414 199144
rect 174464 196246 174492 199430
rect 174648 198734 174676 199543
rect 174556 198706 174676 198734
rect 174452 196240 174504 196246
rect 174452 196182 174504 196188
rect 174452 195628 174504 195634
rect 174452 195570 174504 195576
rect 174280 194296 174400 194324
rect 174188 191806 174308 191834
rect 174280 191162 174308 191806
rect 173728 180766 173848 180794
rect 173912 191134 174308 191162
rect 173728 153882 173756 180766
rect 173716 153876 173768 153882
rect 173716 153818 173768 153824
rect 172888 150204 172940 150210
rect 172888 150146 172940 150152
rect 173912 150006 173940 191134
rect 174372 191026 174400 194296
rect 174004 190998 174400 191026
rect 173900 150000 173952 150006
rect 173900 149942 173952 149948
rect 174004 149938 174032 190998
rect 174176 190936 174228 190942
rect 174176 190878 174228 190884
rect 174188 150142 174216 190878
rect 174464 190330 174492 195570
rect 174556 193934 174584 198706
rect 174636 197464 174688 197470
rect 174636 197406 174688 197412
rect 174544 193928 174596 193934
rect 174544 193870 174596 193876
rect 174648 192438 174676 197406
rect 174544 192432 174596 192438
rect 174544 192374 174596 192380
rect 174636 192432 174688 192438
rect 174636 192374 174688 192380
rect 174452 190324 174504 190330
rect 174452 190266 174504 190272
rect 174556 151434 174584 192374
rect 174740 190942 174768 199650
rect 174832 195634 174860 199736
rect 174970 199628 174998 200124
rect 175062 199918 175090 200124
rect 175154 199923 175182 200124
rect 175050 199912 175102 199918
rect 175050 199854 175102 199860
rect 175140 199914 175196 199923
rect 175140 199849 175196 199858
rect 175246 199764 175274 200124
rect 174924 199600 174998 199628
rect 175200 199736 175274 199764
rect 174924 195945 174952 199600
rect 175096 199572 175148 199578
rect 175096 199514 175148 199520
rect 175002 198520 175058 198529
rect 175002 198455 175058 198464
rect 175016 198082 175044 198455
rect 175004 198076 175056 198082
rect 175004 198018 175056 198024
rect 174910 195936 174966 195945
rect 174910 195871 174966 195880
rect 174820 195628 174872 195634
rect 174820 195570 174872 195576
rect 175108 194342 175136 199514
rect 175200 195537 175228 199736
rect 175338 199696 175366 200124
rect 175430 199918 175458 200124
rect 175522 199918 175550 200124
rect 175418 199912 175470 199918
rect 175418 199854 175470 199860
rect 175510 199912 175562 199918
rect 175510 199854 175562 199860
rect 175614 199764 175642 200124
rect 175706 199918 175734 200124
rect 175798 199918 175826 200124
rect 175890 199918 175918 200124
rect 175982 199923 176010 200124
rect 175694 199912 175746 199918
rect 175694 199854 175746 199860
rect 175786 199912 175838 199918
rect 175786 199854 175838 199860
rect 175878 199912 175930 199918
rect 175878 199854 175930 199860
rect 175968 199914 176024 199923
rect 176074 199918 176102 200124
rect 176166 199918 176194 200124
rect 176258 199923 176286 200124
rect 175968 199849 176024 199858
rect 176062 199912 176114 199918
rect 176062 199854 176114 199860
rect 176154 199912 176206 199918
rect 176154 199854 176206 199860
rect 176244 199914 176300 199923
rect 176244 199849 176300 199858
rect 176350 199850 176378 200124
rect 176442 199850 176470 200124
rect 176338 199844 176390 199850
rect 176338 199786 176390 199792
rect 176430 199844 176482 199850
rect 176430 199786 176482 199792
rect 175832 199776 175884 199782
rect 175614 199736 175688 199764
rect 175292 199668 175366 199696
rect 175186 195528 175242 195537
rect 175186 195463 175242 195472
rect 175188 195356 175240 195362
rect 175188 195298 175240 195304
rect 175096 194336 175148 194342
rect 175096 194278 175148 194284
rect 174820 193996 174872 194002
rect 174820 193938 174872 193944
rect 174728 190936 174780 190942
rect 174728 190878 174780 190884
rect 174832 186314 174860 193938
rect 174832 186286 174952 186314
rect 174924 180794 174952 186286
rect 174740 180766 174952 180794
rect 174740 151814 174768 180766
rect 174740 151786 175044 151814
rect 174544 151428 174596 151434
rect 174544 151370 174596 151376
rect 174176 150136 174228 150142
rect 174176 150078 174228 150084
rect 173992 149932 174044 149938
rect 173992 149874 174044 149880
rect 172794 149832 172850 149841
rect 172794 149767 172850 149776
rect 172610 149696 172666 149705
rect 172610 149631 172666 149640
rect 172520 147144 172572 147150
rect 172520 147086 172572 147092
rect 174360 144900 174412 144906
rect 174360 144842 174412 144848
rect 173808 141976 173860 141982
rect 173808 141918 173860 141924
rect 173820 139890 173848 141918
rect 174372 139890 174400 144842
rect 174912 143540 174964 143546
rect 174912 143482 174964 143488
rect 174924 139890 174952 143482
rect 171520 139862 171856 139890
rect 171980 139862 172408 139890
rect 173512 139862 173848 139890
rect 174064 139862 174400 139890
rect 174616 139862 174952 139890
rect 157444 139726 157504 139754
rect 166828 139726 166888 139754
rect 172960 139738 173296 139754
rect 172960 139732 173308 139738
rect 172960 139726 173256 139732
rect 173256 139674 173308 139680
rect 161480 139664 161532 139670
rect 161368 139612 161480 139618
rect 161368 139606 161532 139612
rect 161368 139590 161520 139606
rect 175016 139369 175044 151786
rect 175200 149802 175228 195298
rect 175292 149977 175320 199668
rect 175464 199640 175516 199646
rect 175464 199582 175516 199588
rect 175556 199640 175608 199646
rect 175556 199582 175608 199588
rect 175372 199572 175424 199578
rect 175372 199514 175424 199520
rect 175384 195362 175412 199514
rect 175372 195356 175424 195362
rect 175372 195298 175424 195304
rect 175476 194002 175504 199582
rect 175568 199073 175596 199582
rect 175554 199064 175610 199073
rect 175554 198999 175610 199008
rect 175464 193996 175516 194002
rect 175464 193938 175516 193944
rect 175660 191834 175688 199736
rect 175832 199718 175884 199724
rect 175924 199776 175976 199782
rect 175924 199718 175976 199724
rect 176016 199776 176068 199782
rect 176016 199718 176068 199724
rect 175740 199708 175792 199714
rect 175740 199650 175792 199656
rect 175752 194274 175780 199650
rect 175844 198937 175872 199718
rect 175830 198928 175886 198937
rect 175830 198863 175886 198872
rect 175740 194268 175792 194274
rect 175740 194210 175792 194216
rect 175936 191834 175964 199718
rect 176028 198801 176056 199718
rect 176108 199708 176160 199714
rect 176108 199650 176160 199656
rect 176292 199708 176344 199714
rect 176292 199650 176344 199656
rect 176014 198792 176070 198801
rect 176014 198727 176070 198736
rect 176016 194064 176068 194070
rect 176016 194006 176068 194012
rect 175384 191806 175688 191834
rect 175844 191806 175964 191834
rect 175384 150278 175412 191806
rect 175556 191276 175608 191282
rect 175556 191218 175608 191224
rect 175464 191072 175516 191078
rect 175464 191014 175516 191020
rect 175372 150272 175424 150278
rect 175372 150214 175424 150220
rect 175476 150113 175504 191014
rect 175568 152930 175596 191218
rect 175844 186314 175872 191806
rect 175660 186286 175872 186314
rect 175556 152924 175608 152930
rect 175556 152866 175608 152872
rect 175660 152833 175688 186286
rect 175646 152824 175702 152833
rect 175646 152759 175702 152768
rect 175462 150104 175518 150113
rect 175462 150039 175518 150048
rect 175278 149968 175334 149977
rect 175278 149903 175334 149912
rect 175188 149796 175240 149802
rect 175188 149738 175240 149744
rect 175924 144152 175976 144158
rect 175924 144094 175976 144100
rect 175096 141908 175148 141914
rect 175096 141850 175148 141856
rect 175108 139890 175136 141850
rect 175936 139890 175964 144094
rect 176028 142050 176056 194006
rect 176120 191078 176148 199650
rect 176200 199572 176252 199578
rect 176200 199514 176252 199520
rect 176212 198218 176240 199514
rect 176200 198212 176252 198218
rect 176200 198154 176252 198160
rect 176200 198008 176252 198014
rect 176200 197950 176252 197956
rect 176108 191072 176160 191078
rect 176108 191014 176160 191020
rect 176016 142044 176068 142050
rect 176016 141986 176068 141992
rect 176212 140214 176240 197950
rect 176304 195673 176332 199650
rect 176384 199640 176436 199646
rect 176534 199628 176562 200124
rect 176626 199918 176654 200124
rect 176614 199912 176666 199918
rect 176614 199854 176666 199860
rect 176718 199764 176746 200124
rect 176810 199918 176838 200124
rect 176902 199923 176930 200124
rect 176798 199912 176850 199918
rect 176798 199854 176850 199860
rect 176888 199914 176944 199923
rect 176888 199849 176944 199858
rect 176384 199582 176436 199588
rect 176488 199600 176562 199628
rect 176672 199736 176746 199764
rect 176290 195664 176346 195673
rect 176290 195599 176346 195608
rect 176396 191282 176424 199582
rect 176384 191276 176436 191282
rect 176384 191218 176436 191224
rect 176488 190262 176516 199600
rect 176672 197520 176700 199736
rect 176844 199708 176896 199714
rect 176844 199650 176896 199656
rect 176752 199640 176804 199646
rect 176752 199582 176804 199588
rect 176764 197742 176792 199582
rect 176856 198529 176884 199650
rect 176994 199628 177022 200124
rect 176948 199600 177022 199628
rect 177086 199628 177114 200124
rect 177178 199918 177206 200124
rect 177166 199912 177218 199918
rect 177166 199854 177218 199860
rect 177270 199764 177298 200124
rect 177224 199736 177298 199764
rect 177086 199600 177160 199628
rect 176842 198520 176898 198529
rect 176842 198455 176898 198464
rect 176752 197736 176804 197742
rect 176752 197678 176804 197684
rect 176672 197492 176792 197520
rect 176660 197396 176712 197402
rect 176660 197338 176712 197344
rect 176476 190256 176528 190262
rect 176476 190198 176528 190204
rect 176672 152794 176700 197338
rect 176764 152862 176792 197492
rect 176948 197402 176976 199600
rect 177132 198694 177160 199600
rect 177028 198688 177080 198694
rect 177028 198630 177080 198636
rect 177120 198688 177172 198694
rect 177120 198630 177172 198636
rect 177040 198286 177068 198630
rect 177028 198280 177080 198286
rect 177028 198222 177080 198228
rect 176936 197396 176988 197402
rect 176936 197338 176988 197344
rect 177224 196568 177252 199736
rect 177362 199696 177390 200124
rect 177454 199866 177482 200124
rect 177546 199968 177574 200124
rect 177652 200110 177804 200138
rect 177546 199940 177620 199968
rect 177454 199838 177528 199866
rect 176856 196540 177252 196568
rect 177316 199668 177390 199696
rect 176752 152856 176804 152862
rect 176752 152798 176804 152804
rect 176660 152788 176712 152794
rect 176660 152730 176712 152736
rect 176856 152425 176884 196540
rect 177120 196172 177172 196178
rect 177120 196114 177172 196120
rect 176936 196036 176988 196042
rect 176936 195978 176988 195984
rect 176948 155417 176976 195978
rect 177028 194064 177080 194070
rect 177028 194006 177080 194012
rect 177040 158001 177068 194006
rect 177132 158642 177160 196114
rect 177316 190194 177344 199668
rect 177396 198960 177448 198966
rect 177396 198902 177448 198908
rect 177408 190454 177436 198902
rect 177500 196042 177528 199838
rect 177488 196036 177540 196042
rect 177488 195978 177540 195984
rect 177592 194070 177620 199940
rect 177672 199844 177724 199850
rect 177672 199786 177724 199792
rect 177684 198665 177712 199786
rect 177670 198656 177726 198665
rect 177670 198591 177726 198600
rect 177776 196178 177804 200110
rect 177868 199481 177896 200330
rect 177960 199714 177988 200359
rect 178500 200048 178552 200054
rect 178500 199990 178552 199996
rect 177948 199708 178000 199714
rect 177948 199650 178000 199656
rect 177854 199472 177910 199481
rect 177854 199407 177910 199416
rect 178512 198218 178540 199990
rect 179510 199880 179566 199889
rect 179510 199815 179566 199824
rect 178408 198212 178460 198218
rect 178408 198154 178460 198160
rect 178500 198212 178552 198218
rect 178500 198154 178552 198160
rect 178420 197849 178448 198154
rect 178684 197872 178736 197878
rect 178406 197840 178462 197849
rect 178684 197814 178736 197820
rect 178406 197775 178462 197784
rect 177764 196172 177816 196178
rect 177764 196114 177816 196120
rect 177580 194064 177632 194070
rect 177580 194006 177632 194012
rect 177408 190426 177712 190454
rect 177304 190188 177356 190194
rect 177304 190130 177356 190136
rect 177120 158636 177172 158642
rect 177120 158578 177172 158584
rect 177026 157992 177082 158001
rect 177026 157927 177082 157936
rect 177212 157820 177264 157826
rect 177212 157762 177264 157768
rect 176934 155408 176990 155417
rect 176934 155343 176990 155352
rect 176842 152416 176898 152425
rect 176842 152351 176898 152360
rect 176660 147416 176712 147422
rect 176660 147358 176712 147364
rect 176568 143472 176620 143478
rect 176568 143414 176620 143420
rect 176200 140208 176252 140214
rect 176200 140150 176252 140156
rect 176580 139890 176608 143414
rect 176672 140690 176700 147358
rect 176660 140684 176712 140690
rect 176660 140626 176712 140632
rect 177224 139890 177252 157762
rect 177684 148306 177712 190426
rect 177672 148300 177724 148306
rect 177672 148242 177724 148248
rect 178592 147484 178644 147490
rect 178592 147426 178644 147432
rect 178132 146192 178184 146198
rect 178132 146134 178184 146140
rect 178040 146124 178092 146130
rect 178040 146066 178092 146072
rect 177488 143404 177540 143410
rect 177488 143346 177540 143352
rect 177500 139890 177528 143346
rect 178052 140690 178080 146066
rect 177580 140684 177632 140690
rect 177580 140626 177632 140632
rect 178040 140684 178092 140690
rect 178040 140626 178092 140632
rect 175108 139862 175168 139890
rect 175720 139862 175964 139890
rect 176272 139862 176608 139890
rect 176824 139862 177252 139890
rect 177376 139862 177528 139890
rect 177592 139890 177620 140626
rect 178144 139890 178172 146134
rect 178604 143478 178632 147426
rect 178592 143472 178644 143478
rect 178592 143414 178644 143420
rect 178696 142154 178724 197814
rect 179420 197736 179472 197742
rect 179420 197678 179472 197684
rect 178776 197668 178828 197674
rect 178776 197610 178828 197616
rect 178604 142126 178724 142154
rect 178604 140146 178632 142126
rect 178684 140684 178736 140690
rect 178684 140626 178736 140632
rect 178592 140140 178644 140146
rect 178592 140082 178644 140088
rect 178696 139890 178724 140626
rect 178788 140185 178816 197610
rect 179432 194070 179460 197678
rect 179524 195634 179552 199815
rect 179604 199776 179656 199782
rect 179604 199718 179656 199724
rect 179616 199345 179644 199718
rect 179602 199336 179658 199345
rect 179602 199271 179658 199280
rect 179880 197532 179932 197538
rect 179880 197474 179932 197480
rect 179512 195628 179564 195634
rect 179512 195570 179564 195576
rect 179892 194206 179920 197474
rect 179880 194200 179932 194206
rect 179880 194142 179932 194148
rect 179420 194064 179472 194070
rect 179420 194006 179472 194012
rect 179604 147620 179656 147626
rect 179604 147562 179656 147568
rect 179512 146872 179564 146878
rect 179512 146814 179564 146820
rect 179420 145580 179472 145586
rect 179420 145522 179472 145528
rect 179432 143410 179460 145522
rect 179524 143546 179552 146814
rect 179512 143540 179564 143546
rect 179512 143482 179564 143488
rect 179420 143404 179472 143410
rect 179420 143346 179472 143352
rect 179616 142154 179644 147562
rect 179788 147552 179840 147558
rect 179788 147494 179840 147500
rect 179696 145512 179748 145518
rect 179696 145454 179748 145460
rect 179432 142126 179644 142154
rect 178774 140176 178830 140185
rect 178774 140111 178830 140120
rect 179432 139890 179460 142126
rect 179512 141364 179564 141370
rect 179512 141306 179564 141312
rect 179524 140894 179552 141306
rect 179512 140888 179564 140894
rect 179512 140830 179564 140836
rect 179708 139890 179736 145454
rect 179800 143342 179828 147494
rect 179788 143336 179840 143342
rect 179788 143278 179840 143284
rect 180076 140350 180104 200670
rect 180156 200660 180208 200666
rect 180156 200602 180208 200608
rect 180168 146266 180196 200602
rect 180536 200161 180564 200670
rect 182824 200592 182876 200598
rect 182824 200534 182876 200540
rect 181444 200320 181496 200326
rect 181444 200262 181496 200268
rect 180522 200152 180578 200161
rect 181456 200122 181484 200262
rect 180522 200087 180578 200096
rect 181444 200116 181496 200122
rect 181444 200058 181496 200064
rect 181352 199912 181404 199918
rect 181352 199854 181404 199860
rect 180522 199608 180578 199617
rect 180522 199543 180578 199552
rect 180340 198824 180392 198830
rect 180340 198766 180392 198772
rect 180248 198280 180300 198286
rect 180248 198222 180300 198228
rect 180156 146260 180208 146266
rect 180156 146202 180208 146208
rect 180260 144090 180288 198222
rect 180352 146169 180380 198766
rect 180432 195900 180484 195906
rect 180432 195842 180484 195848
rect 180338 146160 180394 146169
rect 180338 146095 180394 146104
rect 180444 144809 180472 195842
rect 180536 195362 180564 199543
rect 181364 199481 181392 199854
rect 181350 199472 181406 199481
rect 180800 199436 180852 199442
rect 181350 199407 181406 199416
rect 180800 199378 180852 199384
rect 180616 196240 180668 196246
rect 180616 196182 180668 196188
rect 180524 195356 180576 195362
rect 180524 195298 180576 195304
rect 180628 194041 180656 196182
rect 180614 194032 180670 194041
rect 180614 193967 180670 193976
rect 180430 144800 180486 144809
rect 180430 144735 180486 144744
rect 180248 144084 180300 144090
rect 180248 144026 180300 144032
rect 180616 141364 180668 141370
rect 180616 141306 180668 141312
rect 180064 140344 180116 140350
rect 180064 140286 180116 140292
rect 180628 139890 180656 141306
rect 177592 139862 177928 139890
rect 178144 139862 178480 139890
rect 178696 139862 179032 139890
rect 179432 139862 179584 139890
rect 179708 139862 180136 139890
rect 180628 139862 180688 139890
rect 180812 139534 180840 199378
rect 181536 198756 181588 198762
rect 181536 198698 181588 198704
rect 181444 198484 181496 198490
rect 181444 198426 181496 198432
rect 181456 198286 181484 198426
rect 181444 198280 181496 198286
rect 181444 198222 181496 198228
rect 181444 195220 181496 195226
rect 181444 195162 181496 195168
rect 180892 149184 180944 149190
rect 180892 149126 180944 149132
rect 180904 139890 180932 149126
rect 181456 140457 181484 195162
rect 181548 146810 181576 198698
rect 181628 198688 181680 198694
rect 181628 198630 181680 198636
rect 181640 198490 181668 198630
rect 181628 198484 181680 198490
rect 181628 198426 181680 198432
rect 182088 150408 182140 150414
rect 182088 150350 182140 150356
rect 182100 149190 182128 150350
rect 182088 149184 182140 149190
rect 182088 149126 182140 149132
rect 182732 147212 182784 147218
rect 182732 147154 182784 147160
rect 182640 147076 182692 147082
rect 182640 147018 182692 147024
rect 181536 146804 181588 146810
rect 181536 146746 181588 146752
rect 182652 146674 182680 147018
rect 182744 146742 182772 147154
rect 182732 146736 182784 146742
rect 182732 146678 182784 146684
rect 182640 146668 182692 146674
rect 182640 146610 182692 146616
rect 182732 142112 182784 142118
rect 182732 142054 182784 142060
rect 181442 140448 181498 140457
rect 181442 140383 181498 140392
rect 180904 139862 181240 139890
rect 182744 139754 182772 142054
rect 182836 140321 182864 200534
rect 187160 200161 187188 200806
rect 187146 200152 187202 200161
rect 187146 200087 187202 200096
rect 182916 199504 182968 199510
rect 182916 199446 182968 199452
rect 182928 147218 182956 199446
rect 183008 198892 183060 198898
rect 183008 198834 183060 198840
rect 182916 147212 182968 147218
rect 182916 147154 182968 147160
rect 182822 140312 182878 140321
rect 182822 140247 182878 140256
rect 182744 139726 182896 139754
rect 182638 139632 182694 139641
rect 182180 139596 182232 139602
rect 182744 139618 182772 139726
rect 182694 139590 182772 139618
rect 182638 139567 182694 139576
rect 182180 139538 182232 139544
rect 180800 139528 180852 139534
rect 180800 139470 180852 139476
rect 181444 139528 181496 139534
rect 182192 139482 182220 139538
rect 182640 139528 182692 139534
rect 181496 139476 181792 139482
rect 181444 139470 181792 139476
rect 181456 139454 181792 139470
rect 182192 139476 182640 139482
rect 183020 139505 183048 198834
rect 186964 198552 187016 198558
rect 186964 198494 187016 198500
rect 185492 197328 185544 197334
rect 185492 197270 185544 197276
rect 183100 194948 183152 194954
rect 183100 194890 183152 194896
rect 183112 140282 183140 194890
rect 183192 192364 183244 192370
rect 183192 192306 183244 192312
rect 183204 147665 183232 192306
rect 184388 155916 184440 155922
rect 184388 155858 184440 155864
rect 184296 155848 184348 155854
rect 184296 155790 184348 155796
rect 184204 155168 184256 155174
rect 184204 155110 184256 155116
rect 183468 152380 183520 152386
rect 183468 152322 183520 152328
rect 183190 147656 183246 147665
rect 183190 147591 183246 147600
rect 183192 147212 183244 147218
rect 183192 147154 183244 147160
rect 183204 140826 183232 147154
rect 183480 142769 183508 152322
rect 183466 142760 183522 142769
rect 183466 142695 183468 142704
rect 183520 142695 183522 142704
rect 183468 142666 183520 142672
rect 183480 142635 183508 142666
rect 184216 142154 184244 155110
rect 184124 142126 184244 142154
rect 183650 141264 183706 141273
rect 183650 141199 183706 141208
rect 183192 140820 183244 140826
rect 183192 140762 183244 140768
rect 183100 140276 183152 140282
rect 183100 140218 183152 140224
rect 183204 139890 183232 140762
rect 183664 139890 183692 141199
rect 183204 139862 183448 139890
rect 183664 139862 184000 139890
rect 182192 139470 182692 139476
rect 183006 139496 183062 139505
rect 182192 139454 182680 139470
rect 183006 139431 183062 139440
rect 184124 139369 184152 142126
rect 184308 141302 184336 155790
rect 184296 141296 184348 141302
rect 184296 141238 184348 141244
rect 184400 139369 184428 155858
rect 184940 153264 184992 153270
rect 184940 153206 184992 153212
rect 184664 152992 184716 152998
rect 184664 152934 184716 152940
rect 184480 142724 184532 142730
rect 184480 142666 184532 142672
rect 184492 139890 184520 142666
rect 184492 139862 184552 139890
rect 184676 139398 184704 152934
rect 184848 142520 184900 142526
rect 184848 142462 184900 142468
rect 184860 141273 184888 142462
rect 184846 141264 184902 141273
rect 184846 141199 184902 141208
rect 184952 139890 184980 153206
rect 185504 139913 185532 197270
rect 185768 195968 185820 195974
rect 185768 195910 185820 195916
rect 185676 190460 185728 190466
rect 185676 190402 185728 190408
rect 185688 143546 185716 190402
rect 185676 143540 185728 143546
rect 185676 143482 185728 143488
rect 185584 143268 185636 143274
rect 185584 143210 185636 143216
rect 185490 139904 185546 139913
rect 184952 139862 185104 139890
rect 185490 139839 185546 139848
rect 185398 139632 185454 139641
rect 185596 139618 185624 143210
rect 185780 139777 185808 195910
rect 185860 189712 185912 189718
rect 185860 189654 185912 189660
rect 185872 143818 185900 189654
rect 185950 155816 186006 155825
rect 185950 155751 186006 155760
rect 186044 155780 186096 155786
rect 185860 143812 185912 143818
rect 185860 143754 185912 143760
rect 185766 139768 185822 139777
rect 185766 139703 185822 139712
rect 185454 139590 185656 139618
rect 185398 139567 185454 139576
rect 184664 139392 184716 139398
rect 126242 139360 126298 139369
rect 126242 139295 126298 139304
rect 130566 139360 130622 139369
rect 130566 139295 130622 139304
rect 149426 139360 149482 139369
rect 149426 139295 149482 139304
rect 175002 139360 175058 139369
rect 175002 139295 175058 139304
rect 184110 139360 184166 139369
rect 184110 139295 184166 139304
rect 184386 139360 184442 139369
rect 185964 139369 185992 155751
rect 186044 155722 186096 155728
rect 186056 141234 186084 155722
rect 186976 152998 187004 198494
rect 187054 155680 187110 155689
rect 187054 155615 187110 155624
rect 186964 152992 187016 152998
rect 186964 152934 187016 152940
rect 186228 143472 186280 143478
rect 186228 143414 186280 143420
rect 186240 142390 186268 143414
rect 186228 142384 186280 142390
rect 186228 142326 186280 142332
rect 186044 141228 186096 141234
rect 186044 141170 186096 141176
rect 186240 140162 186268 142326
rect 186194 140134 186268 140162
rect 186194 139876 186222 140134
rect 186504 139392 186556 139398
rect 184664 139334 184716 139340
rect 185950 139360 186006 139369
rect 184386 139295 184442 139304
rect 185950 139295 186006 139304
rect 186502 139360 186504 139369
rect 187068 139369 187096 155615
rect 187332 153196 187384 153202
rect 187332 153138 187384 153144
rect 187148 153128 187200 153134
rect 187148 153070 187200 153076
rect 187160 139874 187188 153070
rect 187240 152448 187292 152454
rect 187240 152390 187292 152396
rect 187148 139868 187200 139874
rect 187148 139810 187200 139816
rect 187252 139806 187280 152390
rect 187344 139942 187372 153138
rect 187712 144265 187740 274654
rect 187792 260364 187844 260370
rect 187792 260306 187844 260312
rect 187804 259418 187832 260306
rect 187792 259412 187844 259418
rect 187792 259354 187844 259360
rect 187790 212528 187846 212537
rect 187790 212463 187846 212472
rect 187698 144256 187754 144265
rect 187698 144191 187754 144200
rect 187804 143478 187832 212463
rect 188344 191344 188396 191350
rect 188344 191286 188396 191292
rect 187976 151836 188028 151842
rect 187976 151778 188028 151784
rect 187988 148374 188016 151778
rect 187976 148368 188028 148374
rect 187976 148310 188028 148316
rect 187792 143472 187844 143478
rect 187792 143414 187844 143420
rect 188356 142154 188384 191286
rect 188528 155712 188580 155718
rect 188528 155654 188580 155660
rect 188436 155576 188488 155582
rect 188436 155518 188488 155524
rect 188264 142126 188384 142154
rect 188160 140208 188212 140214
rect 188160 140150 188212 140156
rect 187332 139936 187384 139942
rect 187332 139878 187384 139884
rect 187240 139800 187292 139806
rect 187240 139742 187292 139748
rect 186556 139360 186558 139369
rect 186502 139295 186558 139304
rect 187054 139360 187110 139369
rect 187054 139295 187110 139304
rect 188172 138718 188200 140150
rect 188264 138922 188292 142126
rect 188448 139330 188476 155518
rect 188436 139324 188488 139330
rect 188436 139266 188488 139272
rect 188252 138916 188304 138922
rect 188252 138858 188304 138864
rect 188540 138786 188568 155654
rect 188620 155508 188672 155514
rect 188620 155450 188672 155456
rect 188528 138780 188580 138786
rect 188528 138722 188580 138728
rect 188160 138712 188212 138718
rect 188160 138654 188212 138660
rect 124034 138136 124090 138145
rect 124034 138071 124090 138080
rect 188632 138038 188660 155450
rect 188712 153060 188764 153066
rect 188712 153002 188764 153008
rect 188724 140214 188752 153002
rect 188804 148980 188856 148986
rect 188804 148922 188856 148928
rect 188712 140208 188764 140214
rect 188712 140150 188764 140156
rect 188816 138854 188844 148922
rect 189092 144498 189120 284310
rect 207020 283620 207072 283626
rect 207020 283562 207072 283568
rect 207032 282946 207060 283562
rect 207020 282940 207072 282946
rect 207020 282882 207072 282888
rect 207032 277394 207060 282882
rect 207032 277366 207152 277394
rect 189172 273964 189224 273970
rect 189172 273906 189224 273912
rect 189184 273290 189212 273906
rect 189172 273284 189224 273290
rect 189172 273226 189224 273232
rect 189080 144492 189132 144498
rect 189080 144434 189132 144440
rect 189184 142905 189212 273226
rect 194876 265668 194928 265674
rect 194876 265610 194928 265616
rect 194784 265192 194836 265198
rect 194784 265134 194836 265140
rect 192208 265056 192260 265062
rect 192208 264998 192260 265004
rect 190644 263900 190696 263906
rect 190644 263842 190696 263848
rect 189356 262880 189408 262886
rect 189356 262822 189408 262828
rect 189264 260024 189316 260030
rect 189264 259966 189316 259972
rect 189170 142896 189226 142905
rect 189170 142831 189226 142840
rect 189276 141846 189304 259966
rect 189368 144634 189396 262822
rect 190460 262608 190512 262614
rect 190460 262550 190512 262556
rect 189538 260128 189594 260137
rect 189538 260063 189594 260072
rect 189446 259992 189502 260001
rect 189446 259927 189502 259936
rect 189356 144628 189408 144634
rect 189356 144570 189408 144576
rect 189356 144084 189408 144090
rect 189356 144026 189408 144032
rect 189264 141840 189316 141846
rect 189264 141782 189316 141788
rect 189172 140344 189224 140350
rect 189172 140286 189224 140292
rect 188804 138848 188856 138854
rect 188804 138790 188856 138796
rect 188620 138032 188672 138038
rect 122746 138000 122802 138009
rect 188620 137974 188672 137980
rect 188894 138000 188950 138009
rect 122746 137935 122802 137944
rect 188894 137935 188950 137944
rect 188158 137864 188214 137873
rect 188158 137799 188160 137808
rect 188212 137799 188214 137808
rect 188160 137770 188212 137776
rect 188908 136746 188936 137935
rect 188896 136740 188948 136746
rect 188896 136682 188948 136688
rect 122746 128480 122802 128489
rect 122746 128415 122802 128424
rect 122760 122913 122788 128415
rect 122746 122904 122802 122913
rect 122746 122839 122802 122848
rect 122746 84144 122802 84153
rect 122746 84079 122802 84088
rect 122194 80608 122250 80617
rect 122194 80543 122250 80552
rect 121184 80504 121236 80510
rect 121184 80446 121236 80452
rect 121460 75948 121512 75954
rect 121460 75890 121512 75896
rect 120906 71224 120962 71233
rect 120906 71159 120962 71168
rect 120816 66836 120868 66842
rect 120816 66778 120868 66784
rect 121472 16574 121500 75890
rect 122104 73228 122156 73234
rect 122104 73170 122156 73176
rect 121472 16546 122052 16574
rect 122024 3482 122052 16546
rect 122116 4078 122144 73170
rect 122208 71398 122236 80543
rect 122378 80200 122434 80209
rect 122378 80135 122434 80144
rect 122392 74390 122420 80135
rect 122760 75857 122788 84079
rect 188896 82816 188948 82822
rect 188896 82758 188948 82764
rect 124034 81152 124090 81161
rect 124034 81087 124090 81096
rect 124048 80617 124076 81087
rect 178224 80640 178276 80646
rect 124034 80608 124090 80617
rect 124034 80543 124090 80552
rect 129002 80608 129058 80617
rect 178224 80582 178276 80588
rect 181626 80608 181682 80617
rect 129002 80543 129058 80552
rect 124864 80436 124916 80442
rect 124864 80378 124916 80384
rect 123760 79620 123812 79626
rect 123760 79562 123812 79568
rect 122840 79552 122892 79558
rect 122840 79494 122892 79500
rect 122746 75848 122802 75857
rect 122746 75783 122802 75792
rect 122380 74384 122432 74390
rect 122380 74326 122432 74332
rect 122852 73234 122880 79494
rect 123772 77722 123800 79562
rect 124128 79552 124180 79558
rect 124128 79494 124180 79500
rect 124140 78878 124168 79494
rect 124128 78872 124180 78878
rect 124128 78814 124180 78820
rect 124220 77920 124272 77926
rect 124220 77862 124272 77868
rect 123760 77716 123812 77722
rect 123760 77658 123812 77664
rect 123772 75954 123800 77658
rect 123760 75948 123812 75954
rect 123760 75890 123812 75896
rect 123114 75848 123170 75857
rect 123114 75783 123170 75792
rect 123128 75138 123156 75783
rect 123116 75132 123168 75138
rect 123116 75074 123168 75080
rect 122840 73228 122892 73234
rect 122840 73170 122892 73176
rect 122196 71392 122248 71398
rect 122196 71334 122248 71340
rect 122104 4072 122156 4078
rect 122104 4014 122156 4020
rect 124232 3670 124260 77862
rect 124876 67590 124904 80378
rect 128266 79928 128322 79937
rect 128266 79863 128322 79872
rect 127072 79620 127124 79626
rect 127072 79562 127124 79568
rect 126980 79416 127032 79422
rect 126980 79358 127032 79364
rect 125508 78668 125560 78674
rect 125508 78610 125560 78616
rect 125520 77926 125548 78610
rect 125508 77920 125560 77926
rect 125508 77862 125560 77868
rect 126992 77518 127020 79358
rect 127084 78033 127112 79562
rect 127806 79384 127862 79393
rect 127806 79319 127862 79328
rect 127820 78849 127848 79319
rect 127806 78840 127862 78849
rect 127806 78775 127862 78784
rect 128174 78840 128230 78849
rect 128174 78775 128230 78784
rect 127164 78260 127216 78266
rect 127164 78202 127216 78208
rect 127070 78024 127126 78033
rect 127070 77959 127126 77968
rect 126980 77512 127032 77518
rect 126980 77454 127032 77460
rect 125600 76628 125652 76634
rect 125600 76570 125652 76576
rect 125612 76362 125640 76570
rect 125600 76356 125652 76362
rect 125600 76298 125652 76304
rect 124864 67584 124916 67590
rect 124864 67526 124916 67532
rect 124220 3664 124272 3670
rect 124220 3606 124272 3612
rect 124680 3664 124732 3670
rect 124680 3606 124732 3612
rect 122024 3454 122328 3482
rect 120724 3052 120776 3058
rect 120724 2994 120776 3000
rect 122300 480 122328 3454
rect 123484 3052 123536 3058
rect 123484 2994 123536 3000
rect 123496 480 123524 2994
rect 124692 480 124720 3606
rect 125612 3058 125640 76298
rect 126992 3534 127020 77454
rect 127084 3602 127112 77959
rect 127176 77897 127204 78202
rect 127716 78124 127768 78130
rect 127716 78066 127768 78072
rect 127162 77888 127218 77897
rect 127162 77823 127218 77832
rect 127624 77852 127676 77858
rect 127176 3942 127204 77823
rect 127624 77794 127676 77800
rect 127636 71738 127664 77794
rect 127728 73166 127756 78066
rect 128188 74534 128216 78775
rect 128280 78577 128308 79863
rect 128636 79552 128688 79558
rect 128636 79494 128688 79500
rect 128266 78568 128322 78577
rect 128266 78503 128322 78512
rect 128268 78056 128320 78062
rect 128268 77998 128320 78004
rect 128280 76634 128308 77998
rect 128648 76945 128676 79494
rect 128634 76936 128690 76945
rect 128634 76871 128690 76880
rect 128268 76628 128320 76634
rect 128268 76570 128320 76576
rect 128188 74506 128308 74534
rect 127716 73160 127768 73166
rect 127716 73102 127768 73108
rect 127624 71732 127676 71738
rect 127624 71674 127676 71680
rect 127164 3936 127216 3942
rect 127164 3878 127216 3884
rect 128280 3602 128308 74506
rect 129016 73030 129044 80543
rect 177764 80504 177816 80510
rect 178236 80481 178264 80582
rect 181626 80543 181682 80552
rect 177764 80446 177816 80452
rect 178222 80472 178278 80481
rect 131948 80436 132000 80442
rect 131948 80378 132000 80384
rect 131764 80368 131816 80374
rect 131764 80310 131816 80316
rect 130290 80200 130346 80209
rect 130290 80135 130346 80144
rect 131672 80164 131724 80170
rect 130304 78606 130332 80135
rect 131672 80106 131724 80112
rect 130384 80096 130436 80102
rect 130384 80038 130436 80044
rect 130292 78600 130344 78606
rect 130292 78542 130344 78548
rect 129464 78396 129516 78402
rect 129464 78338 129516 78344
rect 129004 73024 129056 73030
rect 129004 72966 129056 72972
rect 129476 72350 129504 78338
rect 129648 78260 129700 78266
rect 129648 78202 129700 78208
rect 129556 77784 129608 77790
rect 129556 77726 129608 77732
rect 128360 72344 128412 72350
rect 128360 72286 128412 72292
rect 129464 72344 129516 72350
rect 129464 72286 129516 72292
rect 127072 3596 127124 3602
rect 127072 3538 127124 3544
rect 128268 3596 128320 3602
rect 128268 3538 128320 3544
rect 126980 3528 127032 3534
rect 126980 3470 127032 3476
rect 128176 3528 128228 3534
rect 128176 3470 128228 3476
rect 126980 3324 127032 3330
rect 126980 3266 127032 3272
rect 125876 3256 125928 3262
rect 125876 3198 125928 3204
rect 125600 3052 125652 3058
rect 125600 2994 125652 3000
rect 125888 480 125916 3198
rect 126992 480 127020 3266
rect 128188 480 128216 3470
rect 128372 490 128400 72286
rect 129568 70854 129596 77726
rect 129660 77518 129688 78202
rect 129832 78192 129884 78198
rect 129832 78134 129884 78140
rect 129648 77512 129700 77518
rect 129648 77454 129700 77460
rect 129738 75168 129794 75177
rect 129738 75103 129794 75112
rect 128452 70848 128504 70854
rect 128452 70790 128504 70796
rect 129556 70848 129608 70854
rect 129556 70790 129608 70796
rect 128464 3330 128492 70790
rect 129752 3482 129780 75103
rect 129844 4010 129872 78134
rect 129924 76424 129976 76430
rect 129924 76366 129976 76372
rect 129832 4004 129884 4010
rect 129832 3946 129884 3952
rect 129936 3670 129964 76366
rect 130016 75064 130068 75070
rect 130016 75006 130068 75012
rect 130028 3874 130056 75006
rect 130396 73817 130424 80038
rect 130476 80028 130528 80034
rect 130476 79970 130528 79976
rect 130382 73808 130438 73817
rect 130382 73743 130438 73752
rect 130488 73001 130516 79970
rect 130568 79688 130620 79694
rect 130568 79630 130620 79636
rect 131028 79688 131080 79694
rect 131028 79630 131080 79636
rect 130474 72992 130530 73001
rect 130474 72927 130530 72936
rect 130580 70394 130608 79630
rect 131040 79422 131068 79630
rect 130844 79416 130896 79422
rect 130844 79358 130896 79364
rect 131028 79416 131080 79422
rect 131028 79358 131080 79364
rect 130856 78742 130884 79358
rect 131212 79348 131264 79354
rect 131212 79290 131264 79296
rect 130844 78736 130896 78742
rect 130844 78678 130896 78684
rect 130856 78282 130884 78678
rect 130672 78254 130884 78282
rect 130672 75018 130700 78254
rect 130752 78192 130804 78198
rect 130752 78134 130804 78140
rect 130764 77761 130792 78134
rect 131028 78056 131080 78062
rect 131028 77998 131080 78004
rect 130844 77852 130896 77858
rect 130844 77794 130896 77800
rect 130750 77752 130806 77761
rect 130750 77687 130806 77696
rect 130856 76430 130884 77794
rect 130936 77512 130988 77518
rect 130936 77454 130988 77460
rect 130844 76424 130896 76430
rect 130844 76366 130896 76372
rect 130948 75177 130976 77454
rect 131040 76226 131068 77998
rect 131028 76220 131080 76226
rect 131028 76162 131080 76168
rect 131120 75336 131172 75342
rect 131120 75278 131172 75284
rect 130934 75168 130990 75177
rect 130934 75103 130990 75112
rect 130672 74990 131068 75018
rect 130580 70366 130976 70394
rect 130948 3874 130976 70366
rect 130016 3868 130068 3874
rect 130016 3810 130068 3816
rect 130936 3868 130988 3874
rect 130936 3810 130988 3816
rect 131040 3670 131068 74990
rect 129924 3664 129976 3670
rect 129924 3606 129976 3612
rect 131028 3664 131080 3670
rect 131028 3606 131080 3612
rect 129752 3454 130608 3482
rect 128452 3324 128504 3330
rect 128452 3266 128504 3272
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128372 462 128952 490
rect 130580 480 130608 3454
rect 131132 3194 131160 75278
rect 131120 3188 131172 3194
rect 131120 3130 131172 3136
rect 128924 354 128952 462
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131224 354 131252 79290
rect 131684 77994 131712 80106
rect 131304 77988 131356 77994
rect 131304 77930 131356 77936
rect 131672 77988 131724 77994
rect 131672 77930 131724 77936
rect 131316 3806 131344 77930
rect 131396 76628 131448 76634
rect 131396 76570 131448 76576
rect 131304 3800 131356 3806
rect 131304 3742 131356 3748
rect 131408 3738 131436 76570
rect 131488 73636 131540 73642
rect 131488 73578 131540 73584
rect 131396 3732 131448 3738
rect 131396 3674 131448 3680
rect 131500 3262 131528 73578
rect 131776 73137 131804 80310
rect 131960 78334 131988 80378
rect 177776 80374 177804 80446
rect 178222 80407 178278 80416
rect 178406 80472 178462 80481
rect 178406 80407 178462 80416
rect 177764 80368 177816 80374
rect 177764 80310 177816 80316
rect 178316 80368 178368 80374
rect 178316 80310 178368 80316
rect 178132 80232 178184 80238
rect 178132 80174 178184 80180
rect 178040 80164 178092 80170
rect 178040 80106 178092 80112
rect 132052 80022 132388 80050
rect 131948 78328 132000 78334
rect 131948 78270 132000 78276
rect 132052 75886 132080 80022
rect 132466 79914 132494 80036
rect 132558 79937 132586 80036
rect 132420 79886 132494 79914
rect 132544 79928 132600 79937
rect 132314 79792 132370 79801
rect 132314 79727 132316 79736
rect 132368 79727 132370 79736
rect 132316 79698 132368 79704
rect 132316 79348 132368 79354
rect 132316 79290 132368 79296
rect 132328 78606 132356 79290
rect 132316 78600 132368 78606
rect 132316 78542 132368 78548
rect 132224 78328 132276 78334
rect 132224 78270 132276 78276
rect 132236 76906 132264 78270
rect 132316 77988 132368 77994
rect 132316 77930 132368 77936
rect 132224 76900 132276 76906
rect 132224 76842 132276 76848
rect 132040 75880 132092 75886
rect 132040 75822 132092 75828
rect 132328 73642 132356 77930
rect 132316 73636 132368 73642
rect 132316 73578 132368 73584
rect 131762 73128 131818 73137
rect 131762 73063 131818 73072
rect 132420 71058 132448 79886
rect 132650 79898 132678 80036
rect 132544 79863 132600 79872
rect 132638 79892 132690 79898
rect 132638 79834 132690 79840
rect 132742 79778 132770 80036
rect 132592 79756 132644 79762
rect 132592 79698 132644 79704
rect 132696 79750 132770 79778
rect 132834 79778 132862 80036
rect 132926 79971 132954 80036
rect 132912 79962 132968 79971
rect 133018 79966 133046 80036
rect 132912 79897 132968 79906
rect 133006 79960 133058 79966
rect 133006 79902 133058 79908
rect 133110 79830 133138 80036
rect 133098 79824 133150 79830
rect 132958 79792 133014 79801
rect 132834 79750 132908 79778
rect 132500 79484 132552 79490
rect 132500 79426 132552 79432
rect 132408 71052 132460 71058
rect 132408 70994 132460 71000
rect 132512 69562 132540 79426
rect 132500 69556 132552 69562
rect 132500 69498 132552 69504
rect 131580 68536 131632 68542
rect 131580 68478 131632 68484
rect 131592 3398 131620 68478
rect 132604 64666 132632 79698
rect 132696 68542 132724 79750
rect 132776 79688 132828 79694
rect 132776 79630 132828 79636
rect 132788 79422 132816 79630
rect 132776 79416 132828 79422
rect 132776 79358 132828 79364
rect 132880 77625 132908 79750
rect 133098 79766 133150 79772
rect 132958 79727 133014 79736
rect 132972 79694 133000 79727
rect 132960 79688 133012 79694
rect 132960 79630 133012 79636
rect 133052 79688 133104 79694
rect 133202 79676 133230 80036
rect 133294 79898 133322 80036
rect 133386 79898 133414 80036
rect 133478 79898 133506 80036
rect 133570 79971 133598 80036
rect 133556 79962 133612 79971
rect 133662 79966 133690 80036
rect 133754 79971 133782 80036
rect 133282 79892 133334 79898
rect 133282 79834 133334 79840
rect 133374 79892 133426 79898
rect 133374 79834 133426 79840
rect 133466 79892 133518 79898
rect 133556 79897 133612 79906
rect 133650 79960 133702 79966
rect 133650 79902 133702 79908
rect 133740 79962 133796 79971
rect 133740 79897 133796 79906
rect 133846 79898 133874 80036
rect 133938 79898 133966 80036
rect 134030 79971 134058 80036
rect 134016 79962 134072 79971
rect 134122 79966 134150 80036
rect 134214 79971 134242 80036
rect 133466 79834 133518 79840
rect 133834 79892 133886 79898
rect 133834 79834 133886 79840
rect 133926 79892 133978 79898
rect 134016 79897 134072 79906
rect 134110 79960 134162 79966
rect 134110 79902 134162 79908
rect 134200 79962 134256 79971
rect 134200 79897 134256 79906
rect 133926 79834 133978 79840
rect 134306 79812 134334 80036
rect 133326 79792 133382 79801
rect 133740 79792 133796 79801
rect 133662 79750 133740 79778
rect 133662 79744 133690 79750
rect 133326 79727 133382 79736
rect 133052 79630 133104 79636
rect 133156 79648 133230 79676
rect 132866 77616 132922 77625
rect 132866 77551 132922 77560
rect 133064 77294 133092 79630
rect 133156 79558 133184 79648
rect 133144 79552 133196 79558
rect 133144 79494 133196 79500
rect 133144 78464 133196 78470
rect 133144 78406 133196 78412
rect 133156 77450 133184 78406
rect 133144 77444 133196 77450
rect 133144 77386 133196 77392
rect 132880 77266 133092 77294
rect 132776 76016 132828 76022
rect 132776 75958 132828 75964
rect 132788 70174 132816 75958
rect 132880 71641 132908 77266
rect 133340 74534 133368 79727
rect 133616 79716 133690 79744
rect 134154 79792 134210 79801
rect 133740 79727 133796 79736
rect 133880 79756 133932 79762
rect 133512 79688 133564 79694
rect 133512 79630 133564 79636
rect 133420 79620 133472 79626
rect 133420 79562 133472 79568
rect 133432 77489 133460 79562
rect 133418 77480 133474 77489
rect 133418 77415 133474 77424
rect 133524 76022 133552 79630
rect 133616 77353 133644 79716
rect 134154 79727 134210 79736
rect 134260 79784 134334 79812
rect 133880 79698 133932 79704
rect 133788 79688 133840 79694
rect 133788 79630 133840 79636
rect 133602 77344 133658 77353
rect 133602 77279 133658 77288
rect 133512 76016 133564 76022
rect 133512 75958 133564 75964
rect 133800 75342 133828 79630
rect 133788 75336 133840 75342
rect 133788 75278 133840 75284
rect 132972 74506 133368 74534
rect 132972 74322 133000 74506
rect 132960 74316 133012 74322
rect 132960 74258 133012 74264
rect 132866 71632 132922 71641
rect 132866 71567 132922 71576
rect 132972 71482 133000 74258
rect 133892 71774 133920 79698
rect 133972 79620 134024 79626
rect 134168 79608 134196 79727
rect 133972 79562 134024 79568
rect 134076 79580 134196 79608
rect 133984 78033 134012 79562
rect 134076 78674 134104 79580
rect 134260 79506 134288 79784
rect 134398 79744 134426 80036
rect 134490 79966 134518 80036
rect 134582 79971 134610 80036
rect 134478 79960 134530 79966
rect 134478 79902 134530 79908
rect 134568 79962 134624 79971
rect 134568 79897 134624 79906
rect 134674 79898 134702 80036
rect 134662 79892 134714 79898
rect 134662 79834 134714 79840
rect 134766 79778 134794 80036
rect 134858 79966 134886 80036
rect 134950 79966 134978 80036
rect 135042 79971 135070 80036
rect 134846 79960 134898 79966
rect 134846 79902 134898 79908
rect 134938 79960 134990 79966
rect 134938 79902 134990 79908
rect 135028 79962 135084 79971
rect 135028 79897 135084 79906
rect 135134 79778 135162 80036
rect 135226 79830 135254 80036
rect 135318 79937 135346 80036
rect 135304 79928 135360 79937
rect 135304 79863 135360 79872
rect 135410 79830 135438 80036
rect 135502 79830 135530 80036
rect 135594 79937 135622 80036
rect 135580 79928 135636 79937
rect 135686 79898 135714 80036
rect 135778 79898 135806 80036
rect 135580 79863 135636 79872
rect 135674 79892 135726 79898
rect 135674 79834 135726 79840
rect 135766 79892 135818 79898
rect 135766 79834 135818 79840
rect 135870 79830 135898 80036
rect 134168 79478 134288 79506
rect 134352 79716 134426 79744
rect 134720 79750 134794 79778
rect 134996 79750 135162 79778
rect 135214 79824 135266 79830
rect 135214 79766 135266 79772
rect 135398 79824 135450 79830
rect 135398 79766 135450 79772
rect 135490 79824 135542 79830
rect 135490 79766 135542 79772
rect 135858 79824 135910 79830
rect 135858 79766 135910 79772
rect 134064 78668 134116 78674
rect 134064 78610 134116 78616
rect 133970 78024 134026 78033
rect 133970 77959 134026 77968
rect 133972 77920 134024 77926
rect 133972 77862 134024 77868
rect 133984 72457 134012 77862
rect 133970 72448 134026 72457
rect 133970 72383 134026 72392
rect 132880 71454 133000 71482
rect 133800 71746 133920 71774
rect 132776 70168 132828 70174
rect 132776 70110 132828 70116
rect 132684 68536 132736 68542
rect 132684 68478 132736 68484
rect 132592 64660 132644 64666
rect 132592 64602 132644 64608
rect 132788 37942 132816 70110
rect 132776 37936 132828 37942
rect 132776 37878 132828 37884
rect 132880 31074 132908 71454
rect 133800 70394 133828 71746
rect 133984 70394 134012 72383
rect 132972 70366 133828 70394
rect 133892 70366 134012 70394
rect 132972 60722 133000 70366
rect 132960 60716 133012 60722
rect 132960 60658 133012 60664
rect 132868 31068 132920 31074
rect 132868 31010 132920 31016
rect 133892 14482 133920 70366
rect 133972 67380 134024 67386
rect 133972 67322 134024 67328
rect 133984 35222 134012 67322
rect 134064 67312 134116 67318
rect 134064 67254 134116 67260
rect 133972 35216 134024 35222
rect 133972 35158 134024 35164
rect 133880 14476 133932 14482
rect 133880 14418 133932 14424
rect 134076 6186 134104 67254
rect 134168 67250 134196 79478
rect 134248 79416 134300 79422
rect 134248 79358 134300 79364
rect 134260 78810 134288 79358
rect 134248 78804 134300 78810
rect 134248 78746 134300 78752
rect 134352 77330 134380 79716
rect 134524 79620 134576 79626
rect 134524 79562 134576 79568
rect 134616 79620 134668 79626
rect 134616 79562 134668 79568
rect 134260 77302 134380 77330
rect 134260 68474 134288 77302
rect 134536 77194 134564 79562
rect 134628 77926 134656 79562
rect 134616 77920 134668 77926
rect 134616 77862 134668 77868
rect 134614 77344 134670 77353
rect 134614 77279 134670 77288
rect 134352 77166 134564 77194
rect 134248 68468 134300 68474
rect 134248 68410 134300 68416
rect 134156 67244 134208 67250
rect 134156 67186 134208 67192
rect 134168 29646 134196 67186
rect 134352 63510 134380 77166
rect 134524 76900 134576 76906
rect 134524 76842 134576 76848
rect 134432 76560 134484 76566
rect 134432 76502 134484 76508
rect 134444 65890 134472 76502
rect 134536 67386 134564 76842
rect 134524 67380 134576 67386
rect 134524 67322 134576 67328
rect 134628 67318 134656 77279
rect 134720 76673 134748 79750
rect 134892 79688 134944 79694
rect 134892 79630 134944 79636
rect 134800 79552 134852 79558
rect 134800 79494 134852 79500
rect 134812 76906 134840 79494
rect 134800 76900 134852 76906
rect 134800 76842 134852 76848
rect 134706 76664 134762 76673
rect 134706 76599 134762 76608
rect 134904 76566 134932 79630
rect 134892 76560 134944 76566
rect 134892 76502 134944 76508
rect 134996 74118 135024 79750
rect 135962 79744 135990 80036
rect 136054 79966 136082 80036
rect 136042 79960 136094 79966
rect 136042 79902 136094 79908
rect 135962 79716 136036 79744
rect 135076 79688 135128 79694
rect 135076 79630 135128 79636
rect 135536 79688 135588 79694
rect 135588 79648 135668 79676
rect 135536 79630 135588 79636
rect 135088 77586 135116 79630
rect 135168 79620 135220 79626
rect 135168 79562 135220 79568
rect 135352 79620 135404 79626
rect 135352 79562 135404 79568
rect 135076 77580 135128 77586
rect 135076 77522 135128 77528
rect 134984 74112 135036 74118
rect 134984 74054 135036 74060
rect 135180 70394 135208 79562
rect 135364 76634 135392 79562
rect 135444 79416 135496 79422
rect 135444 79358 135496 79364
rect 135352 76628 135404 76634
rect 135352 76570 135404 76576
rect 135456 71534 135484 79358
rect 135536 75948 135588 75954
rect 135536 75890 135588 75896
rect 135444 71528 135496 71534
rect 135444 71470 135496 71476
rect 134996 70366 135208 70394
rect 134996 69766 135024 70366
rect 134984 69760 135036 69766
rect 134984 69702 135036 69708
rect 135352 67584 135404 67590
rect 135352 67526 135404 67532
rect 134616 67312 134668 67318
rect 134616 67254 134668 67260
rect 134432 65884 134484 65890
rect 134432 65826 134484 65832
rect 134340 63504 134392 63510
rect 134340 63446 134392 63452
rect 135260 46980 135312 46986
rect 135260 46922 135312 46928
rect 134156 29640 134208 29646
rect 134156 29582 134208 29588
rect 134064 6180 134116 6186
rect 134064 6122 134116 6128
rect 134156 3460 134208 3466
rect 134156 3402 134208 3408
rect 131580 3392 131632 3398
rect 131580 3334 131632 3340
rect 131488 3256 131540 3262
rect 131488 3198 131540 3204
rect 132960 2984 133012 2990
rect 132960 2926 133012 2932
rect 132972 480 133000 2926
rect 134168 480 134196 3402
rect 135272 480 135300 46922
rect 135364 33794 135392 67526
rect 135548 66978 135576 75890
rect 135640 68678 135668 79648
rect 135812 79620 135864 79626
rect 136008 79608 136036 79716
rect 136146 79676 136174 80036
rect 136238 79903 136266 80036
rect 136224 79894 136280 79903
rect 136224 79829 136280 79838
rect 136330 79676 136358 80036
rect 136422 79898 136450 80036
rect 136514 79898 136542 80036
rect 136606 79966 136634 80036
rect 136594 79960 136646 79966
rect 136594 79902 136646 79908
rect 136410 79892 136462 79898
rect 136410 79834 136462 79840
rect 136502 79892 136554 79898
rect 136502 79834 136554 79840
rect 136456 79756 136508 79762
rect 136698 79744 136726 80036
rect 136456 79698 136508 79704
rect 136652 79716 136726 79744
rect 135812 79562 135864 79568
rect 135916 79580 136036 79608
rect 136100 79648 136174 79676
rect 136284 79648 136358 79676
rect 135824 77489 135852 79562
rect 135810 77480 135866 77489
rect 135810 77415 135866 77424
rect 135720 77308 135772 77314
rect 135720 77250 135772 77256
rect 135628 68672 135680 68678
rect 135628 68614 135680 68620
rect 135536 66972 135588 66978
rect 135536 66914 135588 66920
rect 135352 33788 135404 33794
rect 135352 33730 135404 33736
rect 135548 7614 135576 66914
rect 135732 59362 135760 77250
rect 135812 73432 135864 73438
rect 135812 73374 135864 73380
rect 135824 66094 135852 73374
rect 135916 67590 135944 79580
rect 135996 79484 136048 79490
rect 135996 79426 136048 79432
rect 136008 75002 136036 79426
rect 136100 77314 136128 79648
rect 136180 79552 136232 79558
rect 136180 79494 136232 79500
rect 136088 77308 136140 77314
rect 136088 77250 136140 77256
rect 135996 74996 136048 75002
rect 135996 74938 136048 74944
rect 136192 73438 136220 79494
rect 136284 77294 136312 79648
rect 136468 79608 136496 79698
rect 136468 79580 136588 79608
rect 136456 79484 136508 79490
rect 136456 79426 136508 79432
rect 136284 77266 136404 77294
rect 136272 74996 136324 75002
rect 136272 74938 136324 74944
rect 136180 73432 136232 73438
rect 136180 73374 136232 73380
rect 136284 70394 136312 74938
rect 136376 73846 136404 77266
rect 136468 75954 136496 79426
rect 136456 75948 136508 75954
rect 136456 75890 136508 75896
rect 136560 75410 136588 79580
rect 136652 76634 136680 79716
rect 136790 79642 136818 80036
rect 136882 79966 136910 80036
rect 136974 79971 137002 80036
rect 136870 79960 136922 79966
rect 136870 79902 136922 79908
rect 136960 79962 137016 79971
rect 136960 79897 137016 79906
rect 137066 79898 137094 80036
rect 137158 79937 137186 80036
rect 137144 79928 137200 79937
rect 137054 79892 137106 79898
rect 137144 79863 137200 79872
rect 137054 79834 137106 79840
rect 136916 79824 136968 79830
rect 136914 79792 136916 79801
rect 136968 79792 136970 79801
rect 136914 79727 136970 79736
rect 137100 79756 137152 79762
rect 137250 79744 137278 80036
rect 137342 79966 137370 80036
rect 137330 79960 137382 79966
rect 137330 79902 137382 79908
rect 137434 79898 137462 80036
rect 137526 79937 137554 80036
rect 137618 79966 137646 80036
rect 137606 79960 137658 79966
rect 137512 79928 137568 79937
rect 137422 79892 137474 79898
rect 137606 79902 137658 79908
rect 137512 79863 137568 79872
rect 137422 79834 137474 79840
rect 137710 79812 137738 80036
rect 137466 79792 137522 79801
rect 137250 79716 137324 79744
rect 137466 79727 137522 79736
rect 137664 79784 137738 79812
rect 137100 79698 137152 79704
rect 137008 79688 137060 79694
rect 136914 79656 136970 79665
rect 136790 79614 136864 79642
rect 136836 78305 136864 79614
rect 137008 79630 137060 79636
rect 136914 79591 136970 79600
rect 136928 79422 136956 79591
rect 136916 79416 136968 79422
rect 137020 79393 137048 79630
rect 136916 79358 136968 79364
rect 137006 79384 137062 79393
rect 137006 79319 137062 79328
rect 137008 78736 137060 78742
rect 137008 78678 137060 78684
rect 136822 78296 136878 78305
rect 136822 78231 136878 78240
rect 136822 78160 136878 78169
rect 136822 78095 136878 78104
rect 136640 76628 136692 76634
rect 136640 76570 136692 76576
rect 136640 76084 136692 76090
rect 136640 76026 136692 76032
rect 136548 75404 136600 75410
rect 136548 75346 136600 75352
rect 136364 73840 136416 73846
rect 136364 73782 136416 73788
rect 136652 73166 136680 76026
rect 136836 74534 136864 78095
rect 137020 77858 137048 78678
rect 137008 77852 137060 77858
rect 137008 77794 137060 77800
rect 137008 77308 137060 77314
rect 137008 77250 137060 77256
rect 136836 74506 136956 74534
rect 136640 73160 136692 73166
rect 136640 73102 136692 73108
rect 136192 70366 136312 70394
rect 135904 67584 135956 67590
rect 135904 67526 135956 67532
rect 136192 67114 136220 70366
rect 136180 67108 136232 67114
rect 136180 67050 136232 67056
rect 135812 66088 135864 66094
rect 135812 66030 135864 66036
rect 135720 59356 135772 59362
rect 135720 59298 135772 59304
rect 136652 42090 136680 73102
rect 136928 66162 136956 74506
rect 136916 66156 136968 66162
rect 136916 66098 136968 66104
rect 137020 60586 137048 77250
rect 137112 68814 137140 79698
rect 137190 79656 137246 79665
rect 137190 79591 137246 79600
rect 137204 77654 137232 79591
rect 137192 77648 137244 77654
rect 137192 77590 137244 77596
rect 137296 77314 137324 79716
rect 137374 78704 137430 78713
rect 137374 78639 137430 78648
rect 137284 77308 137336 77314
rect 137284 77250 137336 77256
rect 137388 76090 137416 78639
rect 137480 76809 137508 79727
rect 137560 79688 137612 79694
rect 137560 79630 137612 79636
rect 137572 78334 137600 79630
rect 137560 78328 137612 78334
rect 137560 78270 137612 78276
rect 137466 76800 137522 76809
rect 137466 76735 137522 76744
rect 137468 76628 137520 76634
rect 137468 76570 137520 76576
rect 137376 76084 137428 76090
rect 137376 76026 137428 76032
rect 137376 75880 137428 75886
rect 137376 75822 137428 75828
rect 137388 70394 137416 75822
rect 137296 70366 137416 70394
rect 137100 68808 137152 68814
rect 137100 68750 137152 68756
rect 137296 64874 137324 70366
rect 137204 64846 137324 64874
rect 137204 63442 137232 64846
rect 137480 64734 137508 76570
rect 137664 71126 137692 79784
rect 137802 79744 137830 80036
rect 137894 79937 137922 80036
rect 137986 79966 138014 80036
rect 138078 79966 138106 80036
rect 137974 79960 138026 79966
rect 137880 79928 137936 79937
rect 137974 79902 138026 79908
rect 138066 79960 138118 79966
rect 138066 79902 138118 79908
rect 137880 79863 137936 79872
rect 138170 79812 138198 80036
rect 138262 79898 138290 80036
rect 138250 79892 138302 79898
rect 138250 79834 138302 79840
rect 138032 79784 138198 79812
rect 137756 79716 137830 79744
rect 137928 79756 137980 79762
rect 137756 75886 137784 79716
rect 137928 79698 137980 79704
rect 137836 79552 137888 79558
rect 137836 79494 137888 79500
rect 137744 75880 137796 75886
rect 137744 75822 137796 75828
rect 137848 75750 137876 79494
rect 137836 75744 137888 75750
rect 137836 75686 137888 75692
rect 137940 75070 137968 79698
rect 138032 76129 138060 79784
rect 138354 79778 138382 80036
rect 138308 79750 138382 79778
rect 138112 79688 138164 79694
rect 138112 79630 138164 79636
rect 138018 76120 138074 76129
rect 138018 76055 138074 76064
rect 138020 76016 138072 76022
rect 138020 75958 138072 75964
rect 137928 75064 137980 75070
rect 137928 75006 137980 75012
rect 138032 71738 138060 75958
rect 138124 75177 138152 79630
rect 138204 78192 138256 78198
rect 138204 78134 138256 78140
rect 138110 75168 138166 75177
rect 138110 75103 138166 75112
rect 138216 72418 138244 78134
rect 138308 75274 138336 79750
rect 138446 79744 138474 80036
rect 138538 79966 138566 80036
rect 138526 79960 138578 79966
rect 138630 79937 138658 80036
rect 138526 79902 138578 79908
rect 138616 79928 138672 79937
rect 138616 79863 138672 79872
rect 138722 79812 138750 80036
rect 138676 79784 138750 79812
rect 138446 79716 138520 79744
rect 138388 79484 138440 79490
rect 138388 79426 138440 79432
rect 138296 75268 138348 75274
rect 138296 75210 138348 75216
rect 138204 72412 138256 72418
rect 138204 72354 138256 72360
rect 138216 71774 138244 72354
rect 138124 71746 138244 71774
rect 138020 71732 138072 71738
rect 138020 71674 138072 71680
rect 137652 71120 137704 71126
rect 137652 71062 137704 71068
rect 137468 64728 137520 64734
rect 137468 64670 137520 64676
rect 137192 63436 137244 63442
rect 137192 63378 137244 63384
rect 137008 60580 137060 60586
rect 137008 60522 137060 60528
rect 136640 42084 136692 42090
rect 136640 42026 136692 42032
rect 138020 39024 138072 39030
rect 138020 38966 138072 38972
rect 135536 7608 135588 7614
rect 135536 7550 135588 7556
rect 138032 6914 138060 38966
rect 138124 10334 138152 71746
rect 138296 71732 138348 71738
rect 138296 71674 138348 71680
rect 138308 39370 138336 71674
rect 138400 55214 138428 79426
rect 138492 78674 138520 79716
rect 138572 79620 138624 79626
rect 138572 79562 138624 79568
rect 138480 78668 138532 78674
rect 138480 78610 138532 78616
rect 138584 77110 138612 79562
rect 138572 77104 138624 77110
rect 138572 77046 138624 77052
rect 138676 76129 138704 79784
rect 138814 79744 138842 80036
rect 138906 79966 138934 80036
rect 138998 79966 139026 80036
rect 139090 79971 139118 80036
rect 138894 79960 138946 79966
rect 138894 79902 138946 79908
rect 138986 79960 139038 79966
rect 138986 79902 139038 79908
rect 139076 79962 139132 79971
rect 139182 79966 139210 80036
rect 139274 79966 139302 80036
rect 139076 79897 139132 79906
rect 139170 79960 139222 79966
rect 139170 79902 139222 79908
rect 139262 79960 139314 79966
rect 139262 79902 139314 79908
rect 139366 79778 139394 80036
rect 139320 79750 139394 79778
rect 138814 79716 138888 79744
rect 138860 79676 138888 79716
rect 139124 79688 139176 79694
rect 138860 79648 138980 79676
rect 138846 79520 138902 79529
rect 138846 79455 138902 79464
rect 138756 78668 138808 78674
rect 138756 78610 138808 78616
rect 138662 76120 138718 76129
rect 138662 76055 138718 76064
rect 138768 76022 138796 78610
rect 138756 76016 138808 76022
rect 138756 75958 138808 75964
rect 138860 75954 138888 79455
rect 138952 77897 138980 79648
rect 139122 79656 139124 79665
rect 139176 79656 139178 79665
rect 139320 79608 139348 79750
rect 139458 79642 139486 80036
rect 139550 79937 139578 80036
rect 139536 79928 139592 79937
rect 139536 79863 139592 79872
rect 139642 79676 139670 80036
rect 139734 79966 139762 80036
rect 139826 79966 139854 80036
rect 139722 79960 139774 79966
rect 139722 79902 139774 79908
rect 139814 79960 139866 79966
rect 139918 79937 139946 80036
rect 140010 79966 140038 80036
rect 139998 79960 140050 79966
rect 139814 79902 139866 79908
rect 139904 79928 139960 79937
rect 139998 79902 140050 79908
rect 140102 79898 140130 80036
rect 139904 79863 139960 79872
rect 140090 79892 140142 79898
rect 140090 79834 140142 79840
rect 139768 79756 139820 79762
rect 139768 79698 139820 79704
rect 139412 79626 139486 79642
rect 139122 79591 139178 79600
rect 139228 79580 139348 79608
rect 139400 79620 139486 79626
rect 139032 79552 139084 79558
rect 139032 79494 139084 79500
rect 139044 78198 139072 79494
rect 139122 79384 139178 79393
rect 139122 79319 139178 79328
rect 139032 78192 139084 78198
rect 139032 78134 139084 78140
rect 138938 77888 138994 77897
rect 138938 77823 138994 77832
rect 138480 75948 138532 75954
rect 138480 75890 138532 75896
rect 138848 75948 138900 75954
rect 138848 75890 138900 75896
rect 138492 64802 138520 75890
rect 138754 75848 138810 75857
rect 138754 75783 138810 75792
rect 138768 69698 138796 75783
rect 138848 75268 138900 75274
rect 138848 75210 138900 75216
rect 138756 69692 138808 69698
rect 138756 69634 138808 69640
rect 138860 67182 138888 75210
rect 139136 72690 139164 79319
rect 139228 75614 139256 79580
rect 139452 79614 139486 79620
rect 139596 79648 139670 79676
rect 139400 79562 139452 79568
rect 139308 79484 139360 79490
rect 139308 79426 139360 79432
rect 139320 78169 139348 79426
rect 139306 78160 139362 78169
rect 139306 78095 139362 78104
rect 139596 75914 139624 79648
rect 139676 79552 139728 79558
rect 139676 79494 139728 79500
rect 139688 76362 139716 79494
rect 139780 78305 139808 79698
rect 139952 79688 140004 79694
rect 139952 79630 140004 79636
rect 140042 79656 140098 79665
rect 139860 79484 139912 79490
rect 139860 79426 139912 79432
rect 139766 78296 139822 78305
rect 139766 78231 139822 78240
rect 139676 76356 139728 76362
rect 139676 76298 139728 76304
rect 139674 76256 139730 76265
rect 139674 76191 139730 76200
rect 139412 75886 139624 75914
rect 139216 75608 139268 75614
rect 139216 75550 139268 75556
rect 139412 73982 139440 75886
rect 139400 73976 139452 73982
rect 139400 73918 139452 73924
rect 139124 72684 139176 72690
rect 139124 72626 139176 72632
rect 139688 68338 139716 76191
rect 139768 75268 139820 75274
rect 139768 75210 139820 75216
rect 139676 68332 139728 68338
rect 139676 68274 139728 68280
rect 138848 67176 138900 67182
rect 138848 67118 138900 67124
rect 138480 64796 138532 64802
rect 138480 64738 138532 64744
rect 138664 62824 138716 62830
rect 138664 62766 138716 62772
rect 138388 55208 138440 55214
rect 138388 55150 138440 55156
rect 138296 39364 138348 39370
rect 138296 39306 138348 39312
rect 138112 10328 138164 10334
rect 138112 10270 138164 10276
rect 138032 6886 138612 6914
rect 137652 3732 137704 3738
rect 137652 3674 137704 3680
rect 136456 3188 136508 3194
rect 136456 3130 136508 3136
rect 136468 480 136496 3130
rect 137664 480 137692 3674
rect 138584 3482 138612 6886
rect 138676 3738 138704 62766
rect 139780 60654 139808 75210
rect 139872 66026 139900 79426
rect 139964 75342 139992 79630
rect 140194 79642 140222 80036
rect 140286 79898 140314 80036
rect 140378 79937 140406 80036
rect 140470 79966 140498 80036
rect 140562 79966 140590 80036
rect 140654 79966 140682 80036
rect 140458 79960 140510 79966
rect 140364 79928 140420 79937
rect 140274 79892 140326 79898
rect 140458 79902 140510 79908
rect 140550 79960 140602 79966
rect 140550 79902 140602 79908
rect 140642 79960 140694 79966
rect 140642 79902 140694 79908
rect 140364 79863 140420 79872
rect 140274 79834 140326 79840
rect 140746 79812 140774 80036
rect 140838 79966 140866 80036
rect 140826 79960 140878 79966
rect 140930 79937 140958 80036
rect 140826 79902 140878 79908
rect 140916 79928 140972 79937
rect 141022 79898 141050 80036
rect 140916 79863 140972 79872
rect 141010 79892 141062 79898
rect 141010 79834 141062 79840
rect 140608 79784 140774 79812
rect 140320 79756 140372 79762
rect 140320 79698 140372 79704
rect 140412 79756 140464 79762
rect 140412 79698 140464 79704
rect 140042 79591 140098 79600
rect 140148 79614 140222 79642
rect 140056 77518 140084 79591
rect 140044 77512 140096 77518
rect 140044 77454 140096 77460
rect 139952 75336 140004 75342
rect 139952 75278 140004 75284
rect 140148 72282 140176 79614
rect 140228 79484 140280 79490
rect 140228 79426 140280 79432
rect 140240 78674 140268 79426
rect 140228 78668 140280 78674
rect 140228 78610 140280 78616
rect 140332 75274 140360 79698
rect 140320 75268 140372 75274
rect 140320 75210 140372 75216
rect 140136 72276 140188 72282
rect 140136 72218 140188 72224
rect 140424 70394 140452 79698
rect 140608 79608 140636 79784
rect 141114 79744 141142 80036
rect 140976 79716 141142 79744
rect 140688 79688 140740 79694
rect 140688 79630 140740 79636
rect 140516 79580 140636 79608
rect 140516 71330 140544 79580
rect 140700 79529 140728 79630
rect 140872 79620 140924 79626
rect 140872 79562 140924 79568
rect 140686 79520 140742 79529
rect 140596 79484 140648 79490
rect 140686 79455 140742 79464
rect 140596 79426 140648 79432
rect 140608 78878 140636 79426
rect 140596 78872 140648 78878
rect 140596 78814 140648 78820
rect 140778 78704 140834 78713
rect 140688 78668 140740 78674
rect 140778 78639 140834 78648
rect 140688 78610 140740 78616
rect 140700 76430 140728 78610
rect 140688 76424 140740 76430
rect 140688 76366 140740 76372
rect 140792 75342 140820 78639
rect 140884 77761 140912 79562
rect 140870 77752 140926 77761
rect 140870 77687 140926 77696
rect 140780 75336 140832 75342
rect 140780 75278 140832 75284
rect 140976 72486 141004 79716
rect 141206 79676 141234 80036
rect 141298 79898 141326 80036
rect 141286 79892 141338 79898
rect 141286 79834 141338 79840
rect 141390 79744 141418 80036
rect 141482 79971 141510 80036
rect 141468 79962 141524 79971
rect 141574 79966 141602 80036
rect 141468 79897 141524 79906
rect 141562 79960 141614 79966
rect 141562 79902 141614 79908
rect 141666 79812 141694 80036
rect 141758 79966 141786 80036
rect 141850 79966 141878 80036
rect 141942 79966 141970 80036
rect 141746 79960 141798 79966
rect 141746 79902 141798 79908
rect 141838 79960 141890 79966
rect 141838 79902 141890 79908
rect 141930 79960 141982 79966
rect 141930 79902 141982 79908
rect 142034 79812 142062 80036
rect 142126 79898 142154 80036
rect 142218 79966 142246 80036
rect 142310 79971 142338 80036
rect 142206 79960 142258 79966
rect 142206 79902 142258 79908
rect 142296 79962 142352 79971
rect 142114 79892 142166 79898
rect 142296 79897 142352 79906
rect 142114 79834 142166 79840
rect 141160 79648 141234 79676
rect 141344 79716 141418 79744
rect 141528 79784 141694 79812
rect 141896 79784 142062 79812
rect 141160 79642 141188 79648
rect 141068 79614 141188 79642
rect 140964 72480 141016 72486
rect 140964 72422 141016 72428
rect 140504 71324 140556 71330
rect 140504 71266 140556 71272
rect 140148 70366 140452 70394
rect 140044 68604 140096 68610
rect 140044 68546 140096 68552
rect 139860 66020 139912 66026
rect 139860 65962 139912 65968
rect 139768 60648 139820 60654
rect 139768 60590 139820 60596
rect 140056 6914 140084 68546
rect 140148 67046 140176 70366
rect 140136 67040 140188 67046
rect 140136 66982 140188 66988
rect 141068 66842 141096 79614
rect 141148 79552 141200 79558
rect 141148 79494 141200 79500
rect 141240 79552 141292 79558
rect 141240 79494 141292 79500
rect 141160 66910 141188 79494
rect 141252 79257 141280 79494
rect 141238 79248 141294 79257
rect 141238 79183 141294 79192
rect 141240 78668 141292 78674
rect 141240 78610 141292 78616
rect 141252 69358 141280 78610
rect 141344 75177 141372 79716
rect 141528 79608 141556 79784
rect 141608 79688 141660 79694
rect 141608 79630 141660 79636
rect 141436 79580 141556 79608
rect 141436 79490 141464 79580
rect 141424 79484 141476 79490
rect 141424 79426 141476 79432
rect 141516 79484 141568 79490
rect 141516 79426 141568 79432
rect 141422 79248 141478 79257
rect 141422 79183 141478 79192
rect 141436 77994 141464 79183
rect 141424 77988 141476 77994
rect 141424 77930 141476 77936
rect 141330 75168 141386 75177
rect 141330 75103 141386 75112
rect 141528 73778 141556 79426
rect 141620 78674 141648 79630
rect 141700 79620 141752 79626
rect 141700 79562 141752 79568
rect 141608 78668 141660 78674
rect 141608 78610 141660 78616
rect 141712 77722 141740 79562
rect 141792 79552 141844 79558
rect 141792 79494 141844 79500
rect 141804 78130 141832 79494
rect 141792 78124 141844 78130
rect 141792 78066 141844 78072
rect 141896 77926 141924 79784
rect 142402 79778 142430 80036
rect 142494 79898 142522 80036
rect 142586 79898 142614 80036
rect 142678 79971 142706 80036
rect 142664 79962 142720 79971
rect 142482 79892 142534 79898
rect 142482 79834 142534 79840
rect 142574 79892 142626 79898
rect 142664 79897 142720 79906
rect 142574 79834 142626 79840
rect 142770 79812 142798 80036
rect 142862 79971 142890 80036
rect 142848 79962 142904 79971
rect 142848 79897 142904 79906
rect 142356 79750 142430 79778
rect 142724 79784 142798 79812
rect 142620 79756 142672 79762
rect 142252 79688 142304 79694
rect 142252 79630 142304 79636
rect 142160 79620 142212 79626
rect 142160 79562 142212 79568
rect 141884 77920 141936 77926
rect 141884 77862 141936 77868
rect 142172 77790 142200 79562
rect 142264 79257 142292 79630
rect 142250 79248 142306 79257
rect 142250 79183 142306 79192
rect 142356 78402 142384 79750
rect 142620 79698 142672 79704
rect 142632 79642 142660 79698
rect 142448 79614 142660 79642
rect 142448 78742 142476 79614
rect 142526 79520 142582 79529
rect 142724 79506 142752 79784
rect 142802 79656 142858 79665
rect 142954 79642 142982 80036
rect 143046 79812 143074 80036
rect 143138 79966 143166 80036
rect 143230 79966 143258 80036
rect 143322 79971 143350 80036
rect 143126 79960 143178 79966
rect 143126 79902 143178 79908
rect 143218 79960 143270 79966
rect 143218 79902 143270 79908
rect 143308 79962 143364 79971
rect 143414 79966 143442 80036
rect 143506 79966 143534 80036
rect 143308 79897 143364 79906
rect 143402 79960 143454 79966
rect 143402 79902 143454 79908
rect 143494 79960 143546 79966
rect 143494 79902 143546 79908
rect 143046 79784 143212 79812
rect 143184 79665 143212 79784
rect 143264 79756 143316 79762
rect 143264 79698 143316 79704
rect 143170 79656 143226 79665
rect 142954 79614 143028 79642
rect 142802 79591 142858 79600
rect 142526 79455 142528 79464
rect 142580 79455 142582 79464
rect 142632 79478 142752 79506
rect 142528 79426 142580 79432
rect 142436 78736 142488 78742
rect 142436 78678 142488 78684
rect 142344 78396 142396 78402
rect 142344 78338 142396 78344
rect 142250 78296 142306 78305
rect 142250 78231 142252 78240
rect 142304 78231 142306 78240
rect 142252 78202 142304 78208
rect 142160 77784 142212 77790
rect 142160 77726 142212 77732
rect 141700 77716 141752 77722
rect 141700 77658 141752 77664
rect 142252 77580 142304 77586
rect 142252 77522 142304 77528
rect 141976 75336 142028 75342
rect 141976 75278 142028 75284
rect 141516 73772 141568 73778
rect 141516 73714 141568 73720
rect 141528 70394 141556 73714
rect 141436 70366 141556 70394
rect 141240 69352 141292 69358
rect 141240 69294 141292 69300
rect 141148 66904 141200 66910
rect 141148 66846 141200 66852
rect 141056 66836 141108 66842
rect 141056 66778 141108 66784
rect 140136 59832 140188 59838
rect 140136 59774 140188 59780
rect 139964 6886 140084 6914
rect 138664 3732 138716 3738
rect 138664 3674 138716 3680
rect 138584 3454 138888 3482
rect 138860 480 138888 3454
rect 139964 3194 139992 6886
rect 140044 3528 140096 3534
rect 140044 3470 140096 3476
rect 139952 3188 140004 3194
rect 139952 3130 140004 3136
rect 140056 480 140084 3470
rect 140148 3466 140176 59774
rect 140136 3460 140188 3466
rect 140136 3402 140188 3408
rect 141240 3052 141292 3058
rect 141240 2994 141292 3000
rect 141252 480 141280 2994
rect 141436 2990 141464 70366
rect 141988 68270 142016 75278
rect 142264 72758 142292 77522
rect 142632 77432 142660 79478
rect 142816 79422 142844 79591
rect 142712 79416 142764 79422
rect 142710 79384 142712 79393
rect 142804 79416 142856 79422
rect 142764 79384 142766 79393
rect 142804 79358 142856 79364
rect 142896 79416 142948 79422
rect 142896 79358 142948 79364
rect 142710 79319 142766 79328
rect 142908 77518 142936 79358
rect 143000 77586 143028 79614
rect 143080 79620 143132 79626
rect 143170 79591 143226 79600
rect 143080 79562 143132 79568
rect 142988 77580 143040 77586
rect 142988 77522 143040 77528
rect 142712 77512 142764 77518
rect 142712 77454 142764 77460
rect 142896 77512 142948 77518
rect 142896 77454 142948 77460
rect 142540 77404 142660 77432
rect 142434 77344 142490 77353
rect 142434 77279 142490 77288
rect 142342 73808 142398 73817
rect 142342 73743 142398 73752
rect 142252 72752 142304 72758
rect 142252 72694 142304 72700
rect 142160 69624 142212 69630
rect 142160 69566 142212 69572
rect 141976 68264 142028 68270
rect 141976 68206 142028 68212
rect 142172 66042 142200 69566
rect 142264 68610 142292 72694
rect 142356 71262 142384 73743
rect 142344 71256 142396 71262
rect 142344 71198 142396 71204
rect 142252 68604 142304 68610
rect 142252 68546 142304 68552
rect 142172 66014 142292 66042
rect 142160 65952 142212 65958
rect 142160 65894 142212 65900
rect 141516 64932 141568 64938
rect 141516 64874 141568 64880
rect 141528 3534 141556 64874
rect 141516 3528 141568 3534
rect 141516 3470 141568 3476
rect 141424 2984 141476 2990
rect 141424 2926 141476 2932
rect 131734 354 131846 480
rect 131224 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142172 354 142200 65894
rect 142264 64938 142292 66014
rect 142252 64932 142304 64938
rect 142252 64874 142304 64880
rect 142356 62830 142384 71198
rect 142448 70106 142476 77279
rect 142436 70100 142488 70106
rect 142436 70042 142488 70048
rect 142344 62824 142396 62830
rect 142344 62766 142396 62772
rect 142448 46986 142476 70042
rect 142540 70038 142568 77404
rect 142620 77308 142672 77314
rect 142620 77250 142672 77256
rect 142528 70032 142580 70038
rect 142528 69974 142580 69980
rect 142540 59838 142568 69974
rect 142632 65958 142660 77250
rect 142724 68746 142752 77454
rect 142986 77344 143042 77353
rect 142986 77279 143042 77288
rect 142896 75268 142948 75274
rect 142896 75210 142948 75216
rect 142908 70394 142936 75210
rect 142816 70366 142936 70394
rect 142816 69902 142844 70366
rect 142804 69896 142856 69902
rect 142804 69838 142856 69844
rect 142712 68740 142764 68746
rect 142712 68682 142764 68688
rect 142712 68400 142764 68406
rect 142712 68342 142764 68348
rect 142620 65952 142672 65958
rect 142620 65894 142672 65900
rect 142528 59832 142580 59838
rect 142528 59774 142580 59780
rect 142436 46980 142488 46986
rect 142436 46922 142488 46928
rect 142724 3058 142752 68342
rect 142816 5574 142844 69838
rect 142896 68740 142948 68746
rect 142896 68682 142948 68688
rect 142908 39030 142936 68682
rect 143000 68406 143028 77279
rect 143092 69630 143120 79562
rect 143170 79520 143226 79529
rect 143170 79455 143226 79464
rect 143184 79354 143212 79455
rect 143172 79348 143224 79354
rect 143172 79290 143224 79296
rect 143276 75274 143304 79698
rect 143356 79688 143408 79694
rect 143598 79676 143626 80036
rect 143690 79744 143718 80036
rect 143782 79971 143810 80036
rect 143768 79962 143824 79971
rect 143768 79897 143824 79906
rect 143874 79898 143902 80036
rect 143966 79898 143994 80036
rect 144058 79971 144086 80036
rect 144044 79962 144100 79971
rect 143862 79892 143914 79898
rect 143862 79834 143914 79840
rect 143954 79892 144006 79898
rect 144044 79897 144100 79906
rect 144150 79898 144178 80036
rect 144242 79971 144270 80036
rect 144228 79962 144284 79971
rect 143954 79834 144006 79840
rect 144138 79892 144190 79898
rect 144228 79897 144284 79906
rect 144334 79898 144362 80036
rect 144426 79966 144454 80036
rect 144518 79966 144546 80036
rect 144414 79960 144466 79966
rect 144414 79902 144466 79908
rect 144506 79960 144558 79966
rect 144506 79902 144558 79908
rect 144610 79898 144638 80036
rect 144702 79937 144730 80036
rect 144688 79928 144744 79937
rect 144138 79834 144190 79840
rect 144322 79892 144374 79898
rect 144322 79834 144374 79840
rect 144598 79892 144650 79898
rect 144688 79863 144690 79872
rect 144598 79834 144650 79840
rect 144742 79863 144744 79872
rect 144690 79834 144742 79840
rect 144414 79824 144466 79830
rect 144288 79772 144414 79778
rect 144702 79803 144730 79834
rect 144288 79766 144466 79772
rect 144092 79756 144144 79762
rect 143690 79716 144040 79744
rect 143356 79630 143408 79636
rect 143552 79648 143626 79676
rect 143368 77314 143396 79630
rect 143552 77450 143580 79648
rect 143816 79620 143868 79626
rect 143816 79562 143868 79568
rect 143632 79552 143684 79558
rect 143632 79494 143684 79500
rect 143722 79520 143778 79529
rect 143540 77444 143592 77450
rect 143540 77386 143592 77392
rect 143356 77308 143408 77314
rect 143356 77250 143408 77256
rect 143354 77072 143410 77081
rect 143354 77007 143410 77016
rect 143368 76974 143396 77007
rect 143356 76968 143408 76974
rect 143356 76910 143408 76916
rect 143368 76566 143396 76910
rect 143448 76764 143500 76770
rect 143448 76706 143500 76712
rect 143356 76560 143408 76566
rect 143356 76502 143408 76508
rect 143460 75954 143488 76706
rect 143448 75948 143500 75954
rect 143448 75890 143500 75896
rect 143264 75268 143316 75274
rect 143264 75210 143316 75216
rect 143080 69624 143132 69630
rect 143080 69566 143132 69572
rect 142988 68400 143040 68406
rect 142988 68342 143040 68348
rect 142896 39024 142948 39030
rect 142896 38966 142948 38972
rect 143552 5710 143580 77386
rect 143644 8974 143672 79494
rect 143722 79455 143778 79464
rect 143736 21418 143764 79455
rect 143828 49706 143856 79562
rect 143908 79552 143960 79558
rect 143908 79494 143960 79500
rect 143920 66230 143948 79494
rect 144012 77450 144040 79716
rect 144092 79698 144144 79704
rect 144288 79750 144454 79766
rect 144104 77489 144132 79698
rect 144184 79688 144236 79694
rect 144184 79630 144236 79636
rect 144090 77480 144146 77489
rect 144000 77444 144052 77450
rect 144090 77415 144146 77424
rect 144000 77386 144052 77392
rect 144092 77376 144144 77382
rect 143998 77344 144054 77353
rect 144092 77318 144144 77324
rect 143998 77279 144054 77288
rect 144012 69970 144040 77279
rect 144000 69964 144052 69970
rect 144000 69906 144052 69912
rect 143908 66224 143960 66230
rect 143908 66166 143960 66172
rect 144104 64870 144132 77318
rect 144196 76906 144224 79630
rect 144288 78441 144316 79750
rect 144794 79744 144822 80036
rect 144886 79966 144914 80036
rect 144874 79960 144926 79966
rect 144874 79902 144926 79908
rect 144978 79812 145006 80036
rect 145070 79971 145098 80036
rect 145056 79962 145112 79971
rect 145162 79966 145190 80036
rect 145254 79966 145282 80036
rect 145346 79966 145374 80036
rect 145056 79897 145112 79906
rect 145150 79960 145202 79966
rect 145150 79902 145202 79908
rect 145242 79960 145294 79966
rect 145242 79902 145294 79908
rect 145334 79960 145386 79966
rect 145438 79937 145466 80036
rect 145334 79902 145386 79908
rect 145424 79928 145480 79937
rect 145424 79863 145480 79872
rect 144932 79784 145006 79812
rect 144932 79778 144960 79784
rect 144748 79716 144822 79744
rect 144886 79750 144960 79778
rect 145196 79756 145248 79762
rect 144460 79688 144512 79694
rect 144460 79630 144512 79636
rect 144274 78432 144330 78441
rect 144274 78367 144330 78376
rect 144184 76900 144236 76906
rect 144184 76842 144236 76848
rect 144288 64874 144316 78367
rect 144472 77625 144500 79630
rect 144552 79416 144604 79422
rect 144552 79358 144604 79364
rect 144458 77616 144514 77625
rect 144458 77551 144514 77560
rect 144368 76900 144420 76906
rect 144368 76842 144420 76848
rect 144380 68542 144408 76842
rect 144564 75041 144592 79358
rect 144748 76945 144776 79716
rect 144886 79676 144914 79750
rect 145530 79744 145558 80036
rect 145622 79966 145650 80036
rect 145714 79971 145742 80036
rect 145610 79960 145662 79966
rect 145610 79902 145662 79908
rect 145700 79962 145756 79971
rect 145700 79897 145756 79906
rect 145806 79898 145834 80036
rect 145898 79966 145926 80036
rect 145990 79966 146018 80036
rect 145886 79960 145938 79966
rect 145886 79902 145938 79908
rect 145978 79960 146030 79966
rect 145978 79902 146030 79908
rect 146082 79898 146110 80036
rect 146174 79898 146202 80036
rect 145794 79892 145846 79898
rect 145794 79834 145846 79840
rect 146070 79892 146122 79898
rect 146070 79834 146122 79840
rect 146162 79892 146214 79898
rect 146162 79834 146214 79840
rect 146266 79778 146294 80036
rect 146358 79966 146386 80036
rect 146450 79966 146478 80036
rect 146346 79960 146398 79966
rect 146346 79902 146398 79908
rect 146438 79960 146490 79966
rect 146438 79902 146490 79908
rect 146542 79898 146570 80036
rect 146634 79966 146662 80036
rect 146726 79966 146754 80036
rect 146818 79966 146846 80036
rect 146622 79960 146674 79966
rect 146622 79902 146674 79908
rect 146714 79960 146766 79966
rect 146714 79902 146766 79908
rect 146806 79960 146858 79966
rect 146806 79902 146858 79908
rect 146530 79892 146582 79898
rect 146530 79834 146582 79840
rect 146910 79830 146938 80036
rect 147002 79966 147030 80036
rect 147094 79966 147122 80036
rect 147186 79966 147214 80036
rect 147278 79971 147306 80036
rect 146990 79960 147042 79966
rect 146990 79902 147042 79908
rect 147082 79960 147134 79966
rect 147082 79902 147134 79908
rect 147174 79960 147226 79966
rect 147174 79902 147226 79908
rect 147264 79962 147320 79971
rect 147264 79897 147320 79906
rect 146898 79824 146950 79830
rect 146358 79784 146478 79812
rect 146358 79778 146386 79784
rect 145840 79756 145892 79762
rect 145530 79716 145604 79744
rect 145196 79698 145248 79704
rect 144886 79648 144960 79676
rect 144932 77858 144960 79648
rect 145010 79520 145066 79529
rect 145010 79455 145066 79464
rect 145024 79286 145052 79455
rect 145012 79280 145064 79286
rect 145012 79222 145064 79228
rect 144920 77852 144972 77858
rect 144920 77794 144972 77800
rect 144734 76936 144790 76945
rect 144734 76871 144790 76880
rect 144920 76628 144972 76634
rect 144920 76570 144972 76576
rect 144550 75032 144606 75041
rect 144550 74967 144606 74976
rect 144368 68536 144420 68542
rect 144368 68478 144420 68484
rect 144092 64864 144144 64870
rect 144092 64806 144144 64812
rect 144196 64846 144316 64874
rect 144104 63578 144132 64806
rect 144092 63572 144144 63578
rect 144092 63514 144144 63520
rect 143816 49700 143868 49706
rect 143816 49642 143868 49648
rect 143724 21412 143776 21418
rect 143724 21354 143776 21360
rect 144196 13122 144224 64846
rect 144380 64054 144408 68478
rect 144368 64048 144420 64054
rect 144368 63990 144420 63996
rect 144276 63572 144328 63578
rect 144276 63514 144328 63520
rect 144288 33862 144316 63514
rect 144276 33856 144328 33862
rect 144276 33798 144328 33804
rect 144932 26926 144960 76570
rect 145024 70394 145052 79222
rect 145208 78849 145236 79698
rect 145380 79688 145432 79694
rect 145380 79630 145432 79636
rect 145194 78840 145250 78849
rect 145194 78775 145250 78784
rect 145392 78538 145420 79630
rect 145472 79484 145524 79490
rect 145472 79426 145524 79432
rect 145380 78532 145432 78538
rect 145380 78474 145432 78480
rect 145392 76362 145420 78474
rect 145380 76356 145432 76362
rect 145380 76298 145432 76304
rect 145378 76256 145434 76265
rect 145378 76191 145434 76200
rect 145392 75954 145420 76191
rect 145380 75948 145432 75954
rect 145380 75890 145432 75896
rect 145024 70366 145144 70394
rect 145116 68950 145144 70366
rect 145104 68944 145156 68950
rect 145104 68886 145156 68892
rect 145012 33856 145064 33862
rect 145012 33798 145064 33804
rect 144920 26920 144972 26926
rect 144920 26862 144972 26868
rect 145024 16574 145052 33798
rect 145484 33794 145512 79426
rect 145576 76498 145604 79716
rect 145840 79698 145892 79704
rect 146116 79756 146168 79762
rect 146266 79750 146386 79778
rect 146450 79778 146478 79784
rect 146450 79750 146524 79778
rect 146898 79766 146950 79772
rect 146116 79698 146168 79704
rect 145656 79552 145708 79558
rect 145656 79494 145708 79500
rect 145564 76492 145616 76498
rect 145564 76434 145616 76440
rect 145564 76356 145616 76362
rect 145564 76298 145616 76304
rect 145576 42090 145604 76298
rect 145668 72690 145696 79494
rect 145748 79416 145800 79422
rect 145748 79358 145800 79364
rect 145760 78792 145788 79358
rect 145852 78946 145880 79698
rect 145932 79688 145984 79694
rect 145932 79630 145984 79636
rect 145840 78940 145892 78946
rect 145840 78882 145892 78888
rect 145760 78764 145880 78792
rect 145746 78704 145802 78713
rect 145746 78639 145802 78648
rect 145760 75478 145788 78639
rect 145852 75818 145880 78764
rect 145840 75812 145892 75818
rect 145840 75754 145892 75760
rect 145748 75472 145800 75478
rect 145748 75414 145800 75420
rect 145656 72684 145708 72690
rect 145656 72626 145708 72632
rect 145656 67584 145708 67590
rect 145656 67526 145708 67532
rect 145564 42084 145616 42090
rect 145564 42026 145616 42032
rect 145668 37942 145696 67526
rect 145760 50386 145788 75414
rect 145852 60722 145880 75754
rect 145944 75206 145972 79630
rect 146128 79082 146156 79698
rect 146208 79688 146260 79694
rect 146208 79630 146260 79636
rect 146116 79076 146168 79082
rect 146116 79018 146168 79024
rect 146024 78940 146076 78946
rect 146024 78882 146076 78888
rect 146036 76634 146064 78882
rect 146024 76628 146076 76634
rect 146024 76570 146076 76576
rect 146024 76492 146076 76498
rect 146024 76434 146076 76440
rect 145932 75200 145984 75206
rect 145932 75142 145984 75148
rect 145944 62286 145972 75142
rect 146036 67590 146064 76434
rect 146220 75177 146248 79630
rect 146300 79620 146352 79626
rect 146300 79562 146352 79568
rect 146392 79620 146444 79626
rect 146392 79562 146444 79568
rect 146312 79014 146340 79562
rect 146300 79008 146352 79014
rect 146300 78950 146352 78956
rect 146404 77178 146432 79562
rect 146392 77172 146444 77178
rect 146392 77114 146444 77120
rect 146300 76560 146352 76566
rect 146300 76502 146352 76508
rect 146206 75168 146262 75177
rect 146206 75103 146262 75112
rect 146024 67584 146076 67590
rect 146024 67526 146076 67532
rect 145932 62280 145984 62286
rect 145932 62222 145984 62228
rect 145840 60716 145892 60722
rect 145840 60658 145892 60664
rect 145748 50380 145800 50386
rect 145748 50322 145800 50328
rect 145656 37936 145708 37942
rect 145656 37878 145708 37884
rect 145472 33788 145524 33794
rect 145472 33730 145524 33736
rect 146312 16574 146340 76502
rect 146404 74866 146432 77114
rect 146496 75313 146524 79750
rect 147370 79744 147398 80036
rect 147462 79971 147490 80036
rect 147448 79962 147504 79971
rect 147448 79897 147504 79906
rect 147554 79830 147582 80036
rect 147542 79824 147594 79830
rect 147646 79812 147674 80036
rect 147738 79971 147766 80036
rect 147724 79962 147780 79971
rect 147724 79897 147780 79906
rect 147646 79784 147720 79812
rect 147542 79766 147594 79772
rect 147324 79716 147398 79744
rect 146576 79688 146628 79694
rect 146668 79688 146720 79694
rect 146576 79630 146628 79636
rect 146666 79656 146668 79665
rect 146720 79656 146722 79665
rect 146588 77042 146616 79630
rect 146666 79591 146722 79600
rect 147220 79620 147272 79626
rect 146576 77036 146628 77042
rect 146576 76978 146628 76984
rect 146588 76566 146616 76978
rect 146576 76560 146628 76566
rect 146576 76502 146628 76508
rect 146482 75304 146538 75313
rect 146680 75274 146708 79591
rect 147220 79562 147272 79568
rect 146760 79552 146812 79558
rect 146760 79494 146812 79500
rect 146772 79257 146800 79494
rect 146852 79484 146904 79490
rect 146852 79426 146904 79432
rect 146758 79248 146814 79257
rect 146864 79218 146892 79426
rect 147036 79416 147088 79422
rect 147036 79358 147088 79364
rect 146758 79183 146814 79192
rect 146852 79212 146904 79218
rect 146852 79154 146904 79160
rect 146482 75239 146538 75248
rect 146668 75268 146720 75274
rect 146392 74860 146444 74866
rect 146392 74802 146444 74808
rect 146496 71097 146524 75239
rect 146668 75210 146720 75216
rect 146864 74534 146892 79154
rect 147048 78792 147076 79358
rect 147232 79150 147260 79562
rect 147220 79144 147272 79150
rect 147220 79086 147272 79092
rect 146772 74506 146892 74534
rect 146956 78764 147076 78792
rect 146482 71088 146538 71097
rect 146482 71023 146538 71032
rect 146772 70394 146800 74506
rect 146956 71534 146984 78764
rect 147036 78668 147088 78674
rect 147036 78610 147088 78616
rect 147048 76838 147076 78610
rect 147036 76832 147088 76838
rect 147036 76774 147088 76780
rect 146944 71528 146996 71534
rect 146944 71470 146996 71476
rect 146496 70366 146800 70394
rect 146956 70394 146984 71470
rect 147048 71126 147076 76774
rect 147232 76498 147260 79086
rect 147324 76702 147352 79716
rect 147496 79688 147548 79694
rect 147496 79630 147548 79636
rect 147588 79688 147640 79694
rect 147692 79665 147720 79784
rect 147830 79778 147858 80036
rect 147922 79971 147950 80036
rect 147908 79962 147964 79971
rect 147908 79897 147964 79906
rect 148014 79778 148042 80036
rect 148106 79966 148134 80036
rect 148094 79960 148146 79966
rect 148094 79902 148146 79908
rect 148198 79812 148226 80036
rect 148290 79830 148318 80036
rect 147830 79750 147904 79778
rect 147588 79630 147640 79636
rect 147678 79656 147734 79665
rect 147404 79552 147456 79558
rect 147404 79494 147456 79500
rect 147416 78674 147444 79494
rect 147404 78668 147456 78674
rect 147404 78610 147456 78616
rect 147508 78554 147536 79630
rect 147416 78526 147536 78554
rect 147312 76696 147364 76702
rect 147312 76638 147364 76644
rect 147220 76492 147272 76498
rect 147220 76434 147272 76440
rect 147036 71120 147088 71126
rect 147036 71062 147088 71068
rect 146956 70366 147260 70394
rect 146496 64874 146524 70366
rect 146944 69964 146996 69970
rect 146944 69906 146996 69912
rect 146404 64846 146524 64874
rect 146404 61402 146432 64846
rect 146392 61396 146444 61402
rect 146392 61338 146444 61344
rect 146956 16574 146984 69906
rect 147036 68944 147088 68950
rect 147036 68886 147088 68892
rect 145024 16546 145512 16574
rect 146312 16546 146800 16574
rect 144184 13116 144236 13122
rect 144184 13058 144236 13064
rect 143632 8968 143684 8974
rect 143632 8910 143684 8916
rect 143540 5704 143592 5710
rect 143540 5646 143592 5652
rect 144736 5704 144788 5710
rect 144736 5646 144788 5652
rect 142804 5568 142856 5574
rect 142804 5510 142856 5516
rect 143540 5568 143592 5574
rect 143540 5510 143592 5516
rect 142712 3052 142764 3058
rect 142712 2994 142764 3000
rect 143552 480 143580 5510
rect 144748 480 144776 5646
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 146772 3482 146800 16546
rect 146864 16546 146984 16574
rect 146864 4078 146892 16546
rect 147048 11778 147076 68886
rect 147128 66224 147180 66230
rect 147128 66166 147180 66172
rect 146956 11750 147076 11778
rect 146852 4072 146904 4078
rect 146852 4014 146904 4020
rect 146956 3806 146984 11750
rect 147140 6914 147168 66166
rect 147232 64874 147260 70366
rect 147324 68338 147352 76638
rect 147312 68332 147364 68338
rect 147312 68274 147364 68280
rect 147232 64846 147352 64874
rect 147220 64048 147272 64054
rect 147220 63990 147272 63996
rect 147048 6886 147168 6914
rect 146944 3800 146996 3806
rect 146944 3742 146996 3748
rect 147048 3738 147076 6886
rect 147036 3732 147088 3738
rect 147036 3674 147088 3680
rect 146772 3454 147168 3482
rect 147232 3466 147260 63990
rect 147324 60042 147352 64846
rect 147416 64190 147444 78526
rect 147494 76256 147550 76265
rect 147494 76191 147550 76200
rect 147508 75682 147536 76191
rect 147496 75676 147548 75682
rect 147496 75618 147548 75624
rect 147508 69698 147536 75618
rect 147600 75449 147628 79630
rect 147876 79626 147904 79750
rect 147968 79750 148042 79778
rect 148152 79784 148226 79812
rect 148278 79824 148330 79830
rect 147678 79591 147734 79600
rect 147864 79620 147916 79626
rect 147864 79562 147916 79568
rect 147968 79393 147996 79750
rect 148048 79688 148100 79694
rect 148046 79656 148048 79665
rect 148100 79656 148102 79665
rect 148046 79591 148102 79600
rect 147770 79384 147826 79393
rect 147770 79319 147826 79328
rect 147954 79384 148010 79393
rect 147954 79319 148010 79328
rect 147586 75440 147642 75449
rect 147586 75375 147642 75384
rect 147496 69692 147548 69698
rect 147496 69634 147548 69640
rect 147404 64184 147456 64190
rect 147404 64126 147456 64132
rect 147784 60734 147812 79319
rect 147864 79280 147916 79286
rect 147862 79248 147864 79257
rect 147916 79248 147918 79257
rect 147862 79183 147918 79192
rect 147876 78810 147904 79183
rect 147864 78804 147916 78810
rect 147864 78746 147916 78752
rect 147954 77480 148010 77489
rect 147954 77415 148010 77424
rect 147968 73154 147996 77415
rect 148060 75138 148088 79591
rect 148048 75132 148100 75138
rect 148048 75074 148100 75080
rect 147968 73126 148088 73154
rect 147864 72956 147916 72962
rect 147864 72898 147916 72904
rect 147876 65618 147904 72898
rect 147956 72616 148008 72622
rect 147956 72558 148008 72564
rect 147968 67114 147996 72558
rect 148060 72554 148088 73126
rect 148152 72826 148180 79784
rect 148278 79766 148330 79772
rect 148382 79676 148410 80036
rect 148474 79898 148502 80036
rect 148462 79892 148514 79898
rect 148462 79834 148514 79840
rect 148566 79744 148594 80036
rect 148336 79648 148410 79676
rect 148520 79716 148594 79744
rect 148232 79620 148284 79626
rect 148232 79562 148284 79568
rect 148140 72820 148192 72826
rect 148140 72762 148192 72768
rect 148048 72548 148100 72554
rect 148048 72490 148100 72496
rect 148244 71466 148272 79562
rect 148336 72214 148364 79648
rect 148520 79608 148548 79716
rect 148658 79676 148686 80036
rect 148750 79778 148778 80036
rect 148842 79898 148870 80036
rect 148830 79892 148882 79898
rect 148830 79834 148882 79840
rect 148750 79750 148824 79778
rect 148658 79648 148732 79676
rect 148428 79580 148548 79608
rect 148428 77489 148456 79580
rect 148508 79484 148560 79490
rect 148508 79426 148560 79432
rect 148414 77480 148470 77489
rect 148414 77415 148470 77424
rect 148416 72820 148468 72826
rect 148416 72762 148468 72768
rect 148324 72208 148376 72214
rect 148324 72150 148376 72156
rect 148232 71460 148284 71466
rect 148232 71402 148284 71408
rect 148428 69902 148456 72762
rect 148520 72622 148548 79426
rect 148704 77353 148732 79648
rect 148690 77344 148746 77353
rect 148690 77279 148746 77288
rect 148796 72962 148824 79750
rect 148934 79744 148962 80036
rect 149026 79971 149054 80036
rect 149012 79962 149068 79971
rect 149118 79966 149146 80036
rect 149012 79897 149068 79906
rect 149106 79960 149158 79966
rect 149106 79902 149158 79908
rect 149210 79830 149238 80036
rect 149302 79966 149330 80036
rect 149394 79971 149422 80036
rect 149290 79960 149342 79966
rect 149290 79902 149342 79908
rect 149380 79962 149436 79971
rect 149486 79966 149514 80036
rect 149578 79966 149606 80036
rect 149380 79897 149436 79906
rect 149474 79960 149526 79966
rect 149474 79902 149526 79908
rect 149566 79960 149618 79966
rect 149566 79902 149618 79908
rect 149198 79824 149250 79830
rect 149198 79766 149250 79772
rect 149520 79824 149572 79830
rect 149520 79766 149572 79772
rect 148888 79716 148962 79744
rect 148888 79529 148916 79716
rect 148966 79656 149022 79665
rect 148966 79591 148968 79600
rect 149020 79591 149022 79600
rect 149152 79620 149204 79626
rect 148968 79562 149020 79568
rect 149152 79562 149204 79568
rect 148874 79520 148930 79529
rect 148874 79455 148930 79464
rect 148876 79416 148928 79422
rect 148876 79358 148928 79364
rect 148784 72956 148836 72962
rect 148784 72898 148836 72904
rect 148508 72616 148560 72622
rect 148508 72558 148560 72564
rect 148508 72208 148560 72214
rect 148508 72150 148560 72156
rect 148416 69896 148468 69902
rect 148416 69838 148468 69844
rect 147956 67108 148008 67114
rect 147956 67050 148008 67056
rect 147864 65612 147916 65618
rect 147864 65554 147916 65560
rect 148324 62280 148376 62286
rect 148324 62222 148376 62228
rect 147692 60706 147812 60734
rect 147312 60036 147364 60042
rect 147312 59978 147364 59984
rect 147692 49162 147720 60706
rect 147680 49156 147732 49162
rect 147680 49098 147732 49104
rect 148336 5114 148364 62222
rect 148416 49700 148468 49706
rect 148416 49642 148468 49648
rect 148428 16574 148456 49642
rect 148520 36922 148548 72150
rect 148692 71460 148744 71466
rect 148692 71402 148744 71408
rect 148600 68876 148652 68882
rect 148600 68818 148652 68824
rect 148612 44878 148640 68818
rect 148704 47666 148732 71402
rect 148888 68882 148916 79358
rect 148980 76702 149008 79562
rect 148968 76696 149020 76702
rect 148968 76638 149020 76644
rect 149164 73250 149192 79562
rect 149244 79552 149296 79558
rect 149244 79494 149296 79500
rect 149256 76634 149284 79494
rect 149336 79484 149388 79490
rect 149336 79426 149388 79432
rect 149244 76628 149296 76634
rect 149244 76570 149296 76576
rect 149164 73222 149284 73250
rect 149152 73092 149204 73098
rect 149152 73034 149204 73040
rect 148968 72548 149020 72554
rect 148968 72490 149020 72496
rect 148980 71058 149008 72490
rect 148968 71052 149020 71058
rect 148968 70994 149020 71000
rect 148876 68876 148928 68882
rect 148876 68818 148928 68824
rect 149164 68610 149192 73034
rect 149256 70990 149284 73222
rect 149348 72894 149376 79426
rect 149428 79416 149480 79422
rect 149428 79358 149480 79364
rect 149440 78441 149468 79358
rect 149426 78432 149482 78441
rect 149426 78367 149482 78376
rect 149336 72888 149388 72894
rect 149336 72830 149388 72836
rect 149244 70984 149296 70990
rect 149244 70926 149296 70932
rect 149256 70786 149284 70926
rect 149244 70780 149296 70786
rect 149244 70722 149296 70728
rect 149532 68814 149560 79766
rect 149670 79608 149698 80036
rect 149762 79676 149790 80036
rect 149854 79966 149882 80036
rect 149842 79960 149894 79966
rect 149842 79902 149894 79908
rect 149946 79778 149974 80036
rect 150038 79966 150066 80036
rect 150130 79966 150158 80036
rect 150026 79960 150078 79966
rect 150026 79902 150078 79908
rect 150118 79960 150170 79966
rect 150222 79937 150250 80036
rect 150118 79902 150170 79908
rect 150208 79928 150264 79937
rect 150208 79863 150264 79872
rect 149946 79750 150020 79778
rect 149762 79648 149928 79676
rect 149670 79580 149744 79608
rect 149612 79484 149664 79490
rect 149612 79426 149664 79432
rect 149624 73098 149652 79426
rect 149716 74662 149744 79580
rect 149796 79552 149848 79558
rect 149796 79494 149848 79500
rect 149704 74656 149756 74662
rect 149704 74598 149756 74604
rect 149704 74520 149756 74526
rect 149704 74462 149756 74468
rect 149612 73092 149664 73098
rect 149612 73034 149664 73040
rect 149520 68808 149572 68814
rect 149520 68750 149572 68756
rect 149152 68604 149204 68610
rect 149152 68546 149204 68552
rect 149532 67658 149560 68750
rect 149520 67652 149572 67658
rect 149520 67594 149572 67600
rect 148692 47660 148744 47666
rect 148692 47602 148744 47608
rect 148600 44872 148652 44878
rect 148600 44814 148652 44820
rect 148508 36916 148560 36922
rect 148508 36858 148560 36864
rect 148428 16546 148548 16574
rect 148336 5086 148456 5114
rect 147140 480 147168 3454
rect 147220 3460 147272 3466
rect 147220 3402 147272 3408
rect 148324 3460 148376 3466
rect 148324 3402 148376 3408
rect 148336 480 148364 3402
rect 148428 3330 148456 5086
rect 148416 3324 148468 3330
rect 148416 3266 148468 3272
rect 148520 3194 148548 16546
rect 149716 16182 149744 74462
rect 149808 73574 149836 79494
rect 149900 73914 149928 79648
rect 149992 74458 150020 79750
rect 150072 79756 150124 79762
rect 150072 79698 150124 79704
rect 150084 74526 150112 79698
rect 150314 79608 150342 80036
rect 150406 79642 150434 80036
rect 150498 79778 150526 80036
rect 150590 79898 150618 80036
rect 150682 79966 150710 80036
rect 150774 79966 150802 80036
rect 150670 79960 150722 79966
rect 150670 79902 150722 79908
rect 150762 79960 150814 79966
rect 150866 79937 150894 80036
rect 150762 79902 150814 79908
rect 150852 79928 150908 79937
rect 150578 79892 150630 79898
rect 150852 79863 150908 79872
rect 150578 79834 150630 79840
rect 150958 79778 150986 80036
rect 150498 79750 150664 79778
rect 150532 79688 150584 79694
rect 150406 79614 150480 79642
rect 150532 79630 150584 79636
rect 150268 79580 150342 79608
rect 150268 78577 150296 79580
rect 150452 78713 150480 79614
rect 150544 79121 150572 79630
rect 150530 79112 150586 79121
rect 150530 79047 150586 79056
rect 150438 78704 150494 78713
rect 150636 78690 150664 79750
rect 150820 79750 150986 79778
rect 150820 79744 150848 79750
rect 150728 79716 150848 79744
rect 150728 78878 150756 79716
rect 151050 79676 151078 80036
rect 151004 79648 151078 79676
rect 151142 79676 151170 80036
rect 151234 79778 151262 80036
rect 151326 79971 151354 80036
rect 151312 79962 151368 79971
rect 151418 79966 151446 80036
rect 151312 79897 151368 79906
rect 151406 79960 151458 79966
rect 151406 79902 151458 79908
rect 151510 79801 151538 80036
rect 151602 79898 151630 80036
rect 151590 79892 151642 79898
rect 151590 79834 151642 79840
rect 151496 79792 151552 79801
rect 151234 79750 151308 79778
rect 151142 79648 151216 79676
rect 150808 79620 150860 79626
rect 150808 79562 150860 79568
rect 150716 78872 150768 78878
rect 150716 78814 150768 78820
rect 150636 78662 150756 78690
rect 150438 78639 150494 78648
rect 150254 78568 150310 78577
rect 150254 78503 150310 78512
rect 150348 76628 150400 76634
rect 150348 76570 150400 76576
rect 150360 75410 150388 76570
rect 150624 76220 150676 76226
rect 150624 76162 150676 76168
rect 150348 75404 150400 75410
rect 150348 75346 150400 75352
rect 150256 74656 150308 74662
rect 150256 74598 150308 74604
rect 150072 74520 150124 74526
rect 150072 74462 150124 74468
rect 149980 74452 150032 74458
rect 149980 74394 150032 74400
rect 149888 73908 149940 73914
rect 149888 73850 149940 73856
rect 149796 73568 149848 73574
rect 149796 73510 149848 73516
rect 149808 64462 149836 73510
rect 149888 67652 149940 67658
rect 149888 67594 149940 67600
rect 149796 64456 149848 64462
rect 149796 64398 149848 64404
rect 149794 56536 149850 56545
rect 149794 56471 149850 56480
rect 149704 16176 149756 16182
rect 149704 16118 149756 16124
rect 149808 3806 149836 56471
rect 149900 17474 149928 67594
rect 149992 32570 150020 74394
rect 150164 72888 150216 72894
rect 150164 72830 150216 72836
rect 150072 70780 150124 70786
rect 150072 70722 150124 70728
rect 150084 47598 150112 70722
rect 150176 51746 150204 72830
rect 150268 71194 150296 74598
rect 150256 71188 150308 71194
rect 150256 71130 150308 71136
rect 150268 56234 150296 71130
rect 150636 69737 150664 76162
rect 150728 70242 150756 78662
rect 150820 75342 150848 79562
rect 151004 76226 151032 79648
rect 151084 79552 151136 79558
rect 151084 79494 151136 79500
rect 150992 76220 151044 76226
rect 150992 76162 151044 76168
rect 150900 75472 150952 75478
rect 150900 75414 150952 75420
rect 150808 75336 150860 75342
rect 150808 75278 150860 75284
rect 150912 74186 150940 75414
rect 150900 74180 150952 74186
rect 150900 74122 150952 74128
rect 151096 70310 151124 79494
rect 151188 70922 151216 79648
rect 151280 75478 151308 79750
rect 151694 79778 151722 80036
rect 151786 79937 151814 80036
rect 151772 79928 151828 79937
rect 151772 79863 151828 79872
rect 151648 79762 151722 79778
rect 151496 79727 151552 79736
rect 151636 79756 151722 79762
rect 151688 79750 151722 79756
rect 151878 79778 151906 80036
rect 151970 79898 151998 80036
rect 151958 79892 152010 79898
rect 151958 79834 152010 79840
rect 151878 79750 151952 79778
rect 151636 79698 151688 79704
rect 151544 79620 151596 79626
rect 151544 79562 151596 79568
rect 151452 79552 151504 79558
rect 151450 79520 151452 79529
rect 151504 79520 151506 79529
rect 151360 79484 151412 79490
rect 151450 79455 151506 79464
rect 151360 79426 151412 79432
rect 151268 75472 151320 75478
rect 151268 75414 151320 75420
rect 151268 75336 151320 75342
rect 151268 75278 151320 75284
rect 151176 70916 151228 70922
rect 151176 70858 151228 70864
rect 151084 70304 151136 70310
rect 151084 70246 151136 70252
rect 150716 70236 150768 70242
rect 150716 70178 150768 70184
rect 150622 69728 150678 69737
rect 150622 69663 150678 69672
rect 150636 69057 150664 69663
rect 150728 69086 150756 70178
rect 150716 69080 150768 69086
rect 150622 69048 150678 69057
rect 150716 69022 150768 69028
rect 150622 68983 150678 68992
rect 150256 56228 150308 56234
rect 150256 56170 150308 56176
rect 150164 51740 150216 51746
rect 150164 51682 150216 51688
rect 150072 47592 150124 47598
rect 150072 47534 150124 47540
rect 149980 32564 150032 32570
rect 149980 32506 150032 32512
rect 149888 17468 149940 17474
rect 149888 17410 149940 17416
rect 151096 5098 151124 70246
rect 151188 12034 151216 70858
rect 151280 66774 151308 75278
rect 151372 71670 151400 79426
rect 151464 76634 151492 79455
rect 151452 76628 151504 76634
rect 151452 76570 151504 76576
rect 151556 74390 151584 79562
rect 151820 79484 151872 79490
rect 151820 79426 151872 79432
rect 151634 79384 151690 79393
rect 151634 79319 151690 79328
rect 151648 77228 151676 79319
rect 151726 79112 151782 79121
rect 151726 79047 151782 79056
rect 151740 78713 151768 79047
rect 151726 78704 151782 78713
rect 151726 78639 151782 78648
rect 151648 77200 151768 77228
rect 151544 74384 151596 74390
rect 151544 74326 151596 74332
rect 151556 73846 151584 74326
rect 151636 74180 151688 74186
rect 151636 74122 151688 74128
rect 151544 73840 151596 73846
rect 151544 73782 151596 73788
rect 151360 71664 151412 71670
rect 151360 71606 151412 71612
rect 151268 66768 151320 66774
rect 151268 66710 151320 66716
rect 151176 12028 151228 12034
rect 151176 11970 151228 11976
rect 151280 10606 151308 66710
rect 151372 39642 151400 71606
rect 151544 69080 151596 69086
rect 151450 69048 151506 69057
rect 151544 69022 151596 69028
rect 151450 68983 151506 68992
rect 151464 42362 151492 68983
rect 151556 46306 151584 69022
rect 151648 53242 151676 74122
rect 151636 53236 151688 53242
rect 151636 53178 151688 53184
rect 151544 46300 151596 46306
rect 151544 46242 151596 46248
rect 151452 42356 151504 42362
rect 151452 42298 151504 42304
rect 151360 39636 151412 39642
rect 151360 39578 151412 39584
rect 151740 32502 151768 77200
rect 151832 74254 151860 79426
rect 151820 74248 151872 74254
rect 151820 74190 151872 74196
rect 151832 73778 151860 74190
rect 151820 73772 151872 73778
rect 151820 73714 151872 73720
rect 151924 70378 151952 79750
rect 152062 79744 152090 80036
rect 152154 79966 152182 80036
rect 152142 79960 152194 79966
rect 152142 79902 152194 79908
rect 152246 79898 152274 80036
rect 152338 79937 152366 80036
rect 152430 79966 152458 80036
rect 152522 79966 152550 80036
rect 152418 79960 152470 79966
rect 152324 79928 152380 79937
rect 152234 79892 152286 79898
rect 152418 79902 152470 79908
rect 152510 79960 152562 79966
rect 152614 79937 152642 80036
rect 152510 79902 152562 79908
rect 152600 79928 152656 79937
rect 152324 79863 152380 79872
rect 152600 79863 152656 79872
rect 152234 79834 152286 79840
rect 152706 79830 152734 80036
rect 152798 79971 152826 80036
rect 152784 79962 152840 79971
rect 152784 79897 152840 79906
rect 152694 79824 152746 79830
rect 152278 79792 152334 79801
rect 152062 79716 152136 79744
rect 152554 79792 152610 79801
rect 152278 79727 152334 79736
rect 152372 79756 152424 79762
rect 152004 79620 152056 79626
rect 152004 79562 152056 79568
rect 152016 73137 152044 79562
rect 152108 78810 152136 79716
rect 152188 79688 152240 79694
rect 152188 79630 152240 79636
rect 152096 78804 152148 78810
rect 152096 78746 152148 78752
rect 152200 77217 152228 79630
rect 152186 77208 152242 77217
rect 152186 77143 152242 77152
rect 152292 75546 152320 79727
rect 152694 79766 152746 79772
rect 152554 79727 152610 79736
rect 152890 79744 152918 80036
rect 152982 79898 153010 80036
rect 153074 79937 153102 80036
rect 153060 79928 153116 79937
rect 152970 79892 153022 79898
rect 153166 79898 153194 80036
rect 153258 79898 153286 80036
rect 153350 79966 153378 80036
rect 153442 79966 153470 80036
rect 153534 79966 153562 80036
rect 153626 79971 153654 80036
rect 153338 79960 153390 79966
rect 153338 79902 153390 79908
rect 153430 79960 153482 79966
rect 153430 79902 153482 79908
rect 153522 79960 153574 79966
rect 153522 79902 153574 79908
rect 153612 79962 153668 79971
rect 153060 79863 153116 79872
rect 153154 79892 153206 79898
rect 152970 79834 153022 79840
rect 153154 79834 153206 79840
rect 153246 79892 153298 79898
rect 153612 79897 153668 79906
rect 153246 79834 153298 79840
rect 153290 79792 153346 79801
rect 152372 79698 152424 79704
rect 152384 76362 152412 79698
rect 152464 79688 152516 79694
rect 152464 79630 152516 79636
rect 152476 77761 152504 79630
rect 152462 77752 152518 77761
rect 152462 77687 152518 77696
rect 152464 77580 152516 77586
rect 152464 77522 152516 77528
rect 152476 77228 152504 77522
rect 152568 77353 152596 79727
rect 152890 79716 152964 79744
rect 153290 79727 153346 79736
rect 153384 79756 153436 79762
rect 152648 79688 152700 79694
rect 152648 79630 152700 79636
rect 152738 79656 152794 79665
rect 152554 77344 152610 77353
rect 152554 77279 152610 77288
rect 152476 77200 152596 77228
rect 152372 76356 152424 76362
rect 152372 76298 152424 76304
rect 152464 75948 152516 75954
rect 152464 75890 152516 75896
rect 152280 75540 152332 75546
rect 152280 75482 152332 75488
rect 152002 73128 152058 73137
rect 152002 73063 152058 73072
rect 151912 70372 151964 70378
rect 151912 70314 151964 70320
rect 151924 61606 151952 70314
rect 151912 61600 151964 61606
rect 151912 61542 151964 61548
rect 151910 46200 151966 46209
rect 151910 46135 151966 46144
rect 151728 32496 151780 32502
rect 151728 32438 151780 32444
rect 151268 10600 151320 10606
rect 151268 10542 151320 10548
rect 151924 6914 151952 46135
rect 151832 6886 151952 6914
rect 151084 5092 151136 5098
rect 151084 5034 151136 5040
rect 150624 3868 150676 3874
rect 150624 3810 150676 3816
rect 149796 3800 149848 3806
rect 149796 3742 149848 3748
rect 149520 3732 149572 3738
rect 149520 3674 149572 3680
rect 148508 3188 148560 3194
rect 148508 3130 148560 3136
rect 149532 480 149560 3674
rect 150636 480 150664 3810
rect 151832 480 151860 6886
rect 152476 3398 152504 75890
rect 152568 74089 152596 77200
rect 152660 76809 152688 79630
rect 152738 79591 152794 79600
rect 152832 79620 152884 79626
rect 152752 77586 152780 79591
rect 152832 79562 152884 79568
rect 152740 77580 152792 77586
rect 152740 77522 152792 77528
rect 152844 77432 152872 79562
rect 152752 77404 152872 77432
rect 152646 76800 152702 76809
rect 152646 76735 152702 76744
rect 152648 75540 152700 75546
rect 152648 75482 152700 75488
rect 152554 74080 152610 74089
rect 152554 74015 152610 74024
rect 152554 73128 152610 73137
rect 152554 73063 152610 73072
rect 152568 6594 152596 73063
rect 152660 64394 152688 75482
rect 152752 69834 152780 77404
rect 152832 76356 152884 76362
rect 152832 76298 152884 76304
rect 152844 73030 152872 76298
rect 152936 74769 152964 79716
rect 153106 77344 153162 77353
rect 153106 77279 153162 77288
rect 152922 74760 152978 74769
rect 152922 74695 152978 74704
rect 152936 74534 152964 74695
rect 152936 74506 153056 74534
rect 152924 73772 152976 73778
rect 152924 73714 152976 73720
rect 152832 73024 152884 73030
rect 152832 72966 152884 72972
rect 152740 69828 152792 69834
rect 152740 69770 152792 69776
rect 152648 64388 152700 64394
rect 152648 64330 152700 64336
rect 152648 60716 152700 60722
rect 152648 60658 152700 60664
rect 152556 6588 152608 6594
rect 152556 6530 152608 6536
rect 152660 3874 152688 60658
rect 152752 31210 152780 69770
rect 152844 38146 152872 72966
rect 152936 43586 152964 73714
rect 153028 57458 153056 74506
rect 153120 60178 153148 77279
rect 153200 76900 153252 76906
rect 153200 76842 153252 76848
rect 153212 64841 153240 76842
rect 153304 67454 153332 79727
rect 153384 79698 153436 79704
rect 153396 74526 153424 79698
rect 153476 79688 153528 79694
rect 153476 79630 153528 79636
rect 153568 79688 153620 79694
rect 153718 79676 153746 80036
rect 153810 79966 153838 80036
rect 153798 79960 153850 79966
rect 153902 79937 153930 80036
rect 153798 79902 153850 79908
rect 153888 79928 153944 79937
rect 153888 79863 153944 79872
rect 153994 79812 154022 80036
rect 154086 79966 154114 80036
rect 154178 79966 154206 80036
rect 154270 79971 154298 80036
rect 154074 79960 154126 79966
rect 154074 79902 154126 79908
rect 154166 79960 154218 79966
rect 154166 79902 154218 79908
rect 154256 79962 154312 79971
rect 154362 79966 154390 80036
rect 154256 79897 154312 79906
rect 154350 79960 154402 79966
rect 154350 79902 154402 79908
rect 154454 79812 154482 80036
rect 153994 79801 154068 79812
rect 154408 79801 154482 79812
rect 153994 79792 154082 79801
rect 153994 79784 154026 79792
rect 153844 79756 153896 79762
rect 154394 79792 154482 79801
rect 154026 79727 154082 79736
rect 154304 79756 154356 79762
rect 153844 79698 153896 79704
rect 154450 79784 154482 79792
rect 154546 79778 154574 80036
rect 154638 79966 154666 80036
rect 154626 79960 154678 79966
rect 154730 79937 154758 80036
rect 154626 79902 154678 79908
rect 154716 79928 154772 79937
rect 154716 79863 154772 79872
rect 154822 79778 154850 80036
rect 154914 79898 154942 80036
rect 155006 79966 155034 80036
rect 155098 79966 155126 80036
rect 155190 79966 155218 80036
rect 155282 79971 155310 80036
rect 154994 79960 155046 79966
rect 154994 79902 155046 79908
rect 155086 79960 155138 79966
rect 155086 79902 155138 79908
rect 155178 79960 155230 79966
rect 155178 79902 155230 79908
rect 155268 79962 155324 79971
rect 154902 79892 154954 79898
rect 155268 79897 155324 79906
rect 154902 79834 154954 79840
rect 155374 79812 155402 80036
rect 155466 79966 155494 80036
rect 155558 79966 155586 80036
rect 155454 79960 155506 79966
rect 155454 79902 155506 79908
rect 155546 79960 155598 79966
rect 155546 79902 155598 79908
rect 155650 79830 155678 80036
rect 155742 79966 155770 80036
rect 155834 79966 155862 80036
rect 155926 79966 155954 80036
rect 155730 79960 155782 79966
rect 155730 79902 155782 79908
rect 155822 79960 155874 79966
rect 155822 79902 155874 79908
rect 155914 79960 155966 79966
rect 155914 79902 155966 79908
rect 155328 79801 155402 79812
rect 155314 79792 155402 79801
rect 154546 79750 154620 79778
rect 154822 79750 154896 79778
rect 154394 79727 154450 79736
rect 154592 79744 154620 79750
rect 154592 79716 154712 79744
rect 154304 79698 154356 79704
rect 153568 79630 153620 79636
rect 153672 79648 153746 79676
rect 153488 77654 153516 79630
rect 153476 77648 153528 77654
rect 153476 77590 153528 77596
rect 153476 77308 153528 77314
rect 153476 77250 153528 77256
rect 153384 74520 153436 74526
rect 153384 74462 153436 74468
rect 153488 69018 153516 77250
rect 153476 69012 153528 69018
rect 153476 68954 153528 68960
rect 153488 67658 153516 68954
rect 153476 67652 153528 67658
rect 153476 67594 153528 67600
rect 153580 67561 153608 79630
rect 153672 71330 153700 79648
rect 153752 79552 153804 79558
rect 153752 79494 153804 79500
rect 153764 75002 153792 79494
rect 153856 77314 153884 79698
rect 153936 79620 153988 79626
rect 153936 79562 153988 79568
rect 153844 77308 153896 77314
rect 153844 77250 153896 77256
rect 153752 74996 153804 75002
rect 153752 74938 153804 74944
rect 153764 74534 153792 74938
rect 153764 74506 153884 74534
rect 153660 71324 153712 71330
rect 153660 71266 153712 71272
rect 153566 67552 153622 67561
rect 153566 67487 153622 67496
rect 153292 67448 153344 67454
rect 153292 67390 153344 67396
rect 153304 66298 153332 67390
rect 153580 66337 153608 67487
rect 153566 66328 153622 66337
rect 153292 66292 153344 66298
rect 153566 66263 153622 66272
rect 153292 66234 153344 66240
rect 153198 64832 153254 64841
rect 153198 64767 153254 64776
rect 153108 60172 153160 60178
rect 153108 60114 153160 60120
rect 153016 57452 153068 57458
rect 153016 57394 153068 57400
rect 152924 43580 152976 43586
rect 152924 43522 152976 43528
rect 152832 38140 152884 38146
rect 152832 38082 152884 38088
rect 152740 31204 152792 31210
rect 152740 31146 152792 31152
rect 153856 20194 153884 74506
rect 153948 70394 153976 79562
rect 154026 79520 154082 79529
rect 154026 79455 154082 79464
rect 154212 79484 154264 79490
rect 154040 74497 154068 79455
rect 154212 79426 154264 79432
rect 154026 74488 154082 74497
rect 154026 74423 154082 74432
rect 153948 70366 154160 70394
rect 154132 70145 154160 70366
rect 154118 70136 154174 70145
rect 154118 70071 154174 70080
rect 153934 66328 153990 66337
rect 153934 66263 153990 66272
rect 154028 66292 154080 66298
rect 153844 20188 153896 20194
rect 153844 20130 153896 20136
rect 153948 13394 153976 66263
rect 154028 66234 154080 66240
rect 154040 18834 154068 66234
rect 154132 25838 154160 70071
rect 154224 70009 154252 79426
rect 154316 76906 154344 79698
rect 154488 79688 154540 79694
rect 154488 79630 154540 79636
rect 154304 76900 154356 76906
rect 154304 76842 154356 76848
rect 154500 76401 154528 79630
rect 154580 79620 154632 79626
rect 154580 79562 154632 79568
rect 154486 76392 154542 76401
rect 154486 76327 154542 76336
rect 154486 74488 154542 74497
rect 154486 74423 154542 74432
rect 154304 71324 154356 71330
rect 154304 71266 154356 71272
rect 154210 70000 154266 70009
rect 154210 69935 154266 69944
rect 154224 69057 154252 69935
rect 154210 69048 154266 69057
rect 154210 68983 154266 68992
rect 154212 67652 154264 67658
rect 154212 67594 154264 67600
rect 154224 27198 154252 67594
rect 154316 67046 154344 71266
rect 154394 69048 154450 69057
rect 154394 68983 154450 68992
rect 154304 67040 154356 67046
rect 154304 66982 154356 66988
rect 154302 64832 154358 64841
rect 154302 64767 154358 64776
rect 154212 27192 154264 27198
rect 154212 27134 154264 27140
rect 154120 25832 154172 25838
rect 154120 25774 154172 25780
rect 154316 24342 154344 64767
rect 154408 36854 154436 68983
rect 154500 61538 154528 74423
rect 154488 61532 154540 61538
rect 154488 61474 154540 61480
rect 154592 49706 154620 79562
rect 154684 77217 154712 79716
rect 154762 79656 154818 79665
rect 154762 79591 154818 79600
rect 154670 77208 154726 77217
rect 154670 77143 154726 77152
rect 154776 76906 154804 79591
rect 154868 79506 154896 79750
rect 155370 79784 155402 79792
rect 155638 79824 155690 79830
rect 156018 79812 156046 80036
rect 155638 79766 155690 79772
rect 155972 79784 156046 79812
rect 155314 79727 155370 79736
rect 155408 79620 155460 79626
rect 155408 79562 155460 79568
rect 155040 79552 155092 79558
rect 154868 79478 154988 79506
rect 155040 79494 155092 79500
rect 155224 79552 155276 79558
rect 155224 79494 155276 79500
rect 154856 79416 154908 79422
rect 154856 79358 154908 79364
rect 154764 76900 154816 76906
rect 154764 76842 154816 76848
rect 154764 76764 154816 76770
rect 154764 76706 154816 76712
rect 154672 74724 154724 74730
rect 154672 74666 154724 74672
rect 154684 60722 154712 74666
rect 154776 63510 154804 76706
rect 154868 64569 154896 79358
rect 154960 78198 154988 79478
rect 154948 78192 155000 78198
rect 154948 78134 155000 78140
rect 154948 76900 155000 76906
rect 154948 76842 155000 76848
rect 154960 65958 154988 76842
rect 155052 76770 155080 79494
rect 155132 79416 155184 79422
rect 155132 79358 155184 79364
rect 155144 77042 155172 79358
rect 155132 77036 155184 77042
rect 155132 76978 155184 76984
rect 155040 76764 155092 76770
rect 155040 76706 155092 76712
rect 155236 72826 155264 79494
rect 155316 79484 155368 79490
rect 155316 79426 155368 79432
rect 155328 74730 155356 79426
rect 155420 77246 155448 79562
rect 155500 79552 155552 79558
rect 155500 79494 155552 79500
rect 155868 79552 155920 79558
rect 155868 79494 155920 79500
rect 155408 77240 155460 77246
rect 155408 77182 155460 77188
rect 155512 76242 155540 79494
rect 155776 79484 155828 79490
rect 155776 79426 155828 79432
rect 155512 76214 155724 76242
rect 155316 74724 155368 74730
rect 155316 74666 155368 74672
rect 155592 74180 155644 74186
rect 155592 74122 155644 74128
rect 155224 72820 155276 72826
rect 155224 72762 155276 72768
rect 154948 65952 155000 65958
rect 154948 65894 155000 65900
rect 154854 64560 154910 64569
rect 154854 64495 154910 64504
rect 154764 63504 154816 63510
rect 154764 63446 154816 63452
rect 154868 60734 154896 64495
rect 154672 60716 154724 60722
rect 154868 60706 155264 60734
rect 154672 60658 154724 60664
rect 154580 49700 154632 49706
rect 154580 49642 154632 49648
rect 154396 36848 154448 36854
rect 154396 36790 154448 36796
rect 154304 24336 154356 24342
rect 154304 24278 154356 24284
rect 155236 20126 155264 60706
rect 155604 29850 155632 74122
rect 155696 72622 155724 76214
rect 155788 72962 155816 79426
rect 155880 74390 155908 79494
rect 155972 78985 156000 79784
rect 156110 79744 156138 80036
rect 156064 79716 156138 79744
rect 155958 78976 156014 78985
rect 156064 78946 156092 79716
rect 156202 79676 156230 80036
rect 156294 79830 156322 80036
rect 156282 79824 156334 79830
rect 156386 79812 156414 80036
rect 156478 79937 156506 80036
rect 156464 79928 156520 79937
rect 156464 79863 156520 79872
rect 156386 79784 156460 79812
rect 156282 79766 156334 79772
rect 156202 79648 156276 79676
rect 156142 79520 156198 79529
rect 156142 79455 156198 79464
rect 155958 78911 156014 78920
rect 156052 78940 156104 78946
rect 156052 78882 156104 78888
rect 155960 78736 156012 78742
rect 155960 78678 156012 78684
rect 155868 74384 155920 74390
rect 155868 74326 155920 74332
rect 155880 74186 155908 74326
rect 155868 74180 155920 74186
rect 155868 74122 155920 74128
rect 155776 72956 155828 72962
rect 155776 72898 155828 72904
rect 155788 72842 155816 72898
rect 155788 72814 155908 72842
rect 155776 72752 155828 72758
rect 155776 72694 155828 72700
rect 155684 72616 155736 72622
rect 155684 72558 155736 72564
rect 155684 65952 155736 65958
rect 155684 65894 155736 65900
rect 155592 29844 155644 29850
rect 155592 29786 155644 29792
rect 155224 20120 155276 20126
rect 155224 20062 155276 20068
rect 155696 20058 155724 65894
rect 155684 20052 155736 20058
rect 155684 19994 155736 20000
rect 154028 18828 154080 18834
rect 154028 18770 154080 18776
rect 155788 14754 155816 72694
rect 155776 14748 155828 14754
rect 155776 14690 155828 14696
rect 153936 13388 153988 13394
rect 153936 13330 153988 13336
rect 155408 13116 155460 13122
rect 155408 13058 155460 13064
rect 153016 4072 153068 4078
rect 153016 4014 153068 4020
rect 152648 3868 152700 3874
rect 152648 3810 152700 3816
rect 152464 3392 152516 3398
rect 152464 3334 152516 3340
rect 153028 480 153056 4014
rect 154212 3188 154264 3194
rect 154212 3130 154264 3136
rect 154224 480 154252 3130
rect 155420 480 155448 13058
rect 155880 9178 155908 72814
rect 155972 52426 156000 78678
rect 156052 78668 156104 78674
rect 156052 78610 156104 78616
rect 156064 56302 156092 78610
rect 156156 57798 156184 79455
rect 156248 78606 156276 79648
rect 156432 78656 156460 79784
rect 156570 79744 156598 80036
rect 156340 78628 156460 78656
rect 156524 79716 156598 79744
rect 156236 78600 156288 78606
rect 156236 78542 156288 78548
rect 156340 70394 156368 78628
rect 156524 71534 156552 79716
rect 156662 79676 156690 80036
rect 156754 79744 156782 80036
rect 156846 79898 156874 80036
rect 156938 79898 156966 80036
rect 157030 79937 157058 80036
rect 157016 79928 157072 79937
rect 156834 79892 156886 79898
rect 156834 79834 156886 79840
rect 156926 79892 156978 79898
rect 157016 79863 157072 79872
rect 156926 79834 156978 79840
rect 156972 79756 157024 79762
rect 156754 79716 156920 79744
rect 156616 79648 156690 79676
rect 156616 72282 156644 79648
rect 156788 79620 156840 79626
rect 156788 79562 156840 79568
rect 156696 79552 156748 79558
rect 156696 79494 156748 79500
rect 156604 72276 156656 72282
rect 156604 72218 156656 72224
rect 156708 72214 156736 79494
rect 156696 72208 156748 72214
rect 156696 72150 156748 72156
rect 156800 71602 156828 79562
rect 156892 78674 156920 79716
rect 157122 79744 157150 80036
rect 157214 79937 157242 80036
rect 157200 79928 157256 79937
rect 157200 79863 157256 79872
rect 157306 79744 157334 80036
rect 157122 79716 157196 79744
rect 156972 79698 157024 79704
rect 156880 78668 156932 78674
rect 156880 78610 156932 78616
rect 156984 78577 157012 79698
rect 157064 78940 157116 78946
rect 157064 78882 157116 78888
rect 156970 78568 157026 78577
rect 156970 78503 157026 78512
rect 156880 72684 156932 72690
rect 156880 72626 156932 72632
rect 156788 71596 156840 71602
rect 156788 71538 156840 71544
rect 156512 71528 156564 71534
rect 156512 71470 156564 71476
rect 156340 70366 156644 70394
rect 156616 66065 156644 70366
rect 156602 66056 156658 66065
rect 156602 65991 156658 66000
rect 156144 57792 156196 57798
rect 156144 57734 156196 57740
rect 156052 56296 156104 56302
rect 156052 56238 156104 56244
rect 155960 52420 156012 52426
rect 155960 52362 156012 52368
rect 156616 40934 156644 65991
rect 156892 60734 156920 72626
rect 157076 72486 157104 78882
rect 157168 77586 157196 79716
rect 157260 79716 157334 79744
rect 157260 78742 157288 79716
rect 157398 79676 157426 80036
rect 157490 79898 157518 80036
rect 157582 79971 157610 80036
rect 157568 79962 157624 79971
rect 157478 79892 157530 79898
rect 157568 79897 157624 79906
rect 157478 79834 157530 79840
rect 157674 79744 157702 80036
rect 157766 79937 157794 80036
rect 157752 79928 157808 79937
rect 157858 79898 157886 80036
rect 157752 79863 157808 79872
rect 157846 79892 157898 79898
rect 157846 79834 157898 79840
rect 157950 79778 157978 80036
rect 158042 79966 158070 80036
rect 158030 79960 158082 79966
rect 158030 79902 158082 79908
rect 158134 79835 158162 80036
rect 158226 79966 158254 80036
rect 158318 79966 158346 80036
rect 158410 79971 158438 80036
rect 158214 79960 158266 79966
rect 158214 79902 158266 79908
rect 158306 79960 158358 79966
rect 158306 79902 158358 79908
rect 158396 79962 158452 79971
rect 158502 79966 158530 80036
rect 158594 79966 158622 80036
rect 158686 79966 158714 80036
rect 158396 79897 158452 79906
rect 158490 79960 158542 79966
rect 158490 79902 158542 79908
rect 158582 79960 158634 79966
rect 158582 79902 158634 79908
rect 158674 79960 158726 79966
rect 158674 79902 158726 79908
rect 158120 79826 158176 79835
rect 157950 79750 158024 79778
rect 158306 79824 158358 79830
rect 158120 79761 158176 79770
rect 158304 79792 158306 79801
rect 158628 79824 158680 79830
rect 158358 79792 158360 79801
rect 157352 79648 157426 79676
rect 157536 79716 157702 79744
rect 157248 78736 157300 78742
rect 157248 78678 157300 78684
rect 157156 77580 157208 77586
rect 157156 77522 157208 77528
rect 157352 76974 157380 79648
rect 157432 79552 157484 79558
rect 157432 79494 157484 79500
rect 157444 78130 157472 79494
rect 157536 78946 157564 79716
rect 157890 79656 157946 79665
rect 157616 79620 157668 79626
rect 157616 79562 157668 79568
rect 157720 79614 157890 79642
rect 157524 78940 157576 78946
rect 157524 78882 157576 78888
rect 157628 78656 157656 79562
rect 157536 78628 157656 78656
rect 157432 78124 157484 78130
rect 157432 78066 157484 78072
rect 157340 76968 157392 76974
rect 157340 76910 157392 76916
rect 157340 76832 157392 76838
rect 157340 76774 157392 76780
rect 157064 72480 157116 72486
rect 157064 72422 157116 72428
rect 157248 72208 157300 72214
rect 157248 72150 157300 72156
rect 157156 71596 157208 71602
rect 157156 71538 157208 71544
rect 157064 71528 157116 71534
rect 157064 71470 157116 71476
rect 156800 60706 156920 60734
rect 156604 40928 156656 40934
rect 156604 40870 156656 40876
rect 155868 9172 155920 9178
rect 155868 9114 155920 9120
rect 156800 3806 156828 60706
rect 157076 23050 157104 71470
rect 157064 23044 157116 23050
rect 157064 22986 157116 22992
rect 157168 14686 157196 71538
rect 157156 14680 157208 14686
rect 157156 14622 157208 14628
rect 157260 13326 157288 72150
rect 157248 13320 157300 13326
rect 157248 13262 157300 13268
rect 157352 11966 157380 76774
rect 157432 75132 157484 75138
rect 157432 75074 157484 75080
rect 157444 51066 157472 75074
rect 157536 59294 157564 78628
rect 157720 77294 157748 79614
rect 157890 79591 157946 79600
rect 157798 79520 157854 79529
rect 157798 79455 157854 79464
rect 157628 77266 157748 77294
rect 157628 63374 157656 77266
rect 157708 76968 157760 76974
rect 157708 76910 157760 76916
rect 157720 71738 157748 76910
rect 157812 73098 157840 79455
rect 157996 79257 158024 79750
rect 158778 79778 158806 80036
rect 158870 79801 158898 80036
rect 158962 79830 158990 80036
rect 159054 79830 159082 80036
rect 159146 79966 159174 80036
rect 159238 79966 159266 80036
rect 159330 79966 159358 80036
rect 159134 79960 159186 79966
rect 159134 79902 159186 79908
rect 159226 79960 159278 79966
rect 159226 79902 159278 79908
rect 159318 79960 159370 79966
rect 159318 79902 159370 79908
rect 158950 79824 159002 79830
rect 158628 79766 158680 79772
rect 158304 79727 158360 79736
rect 158260 79688 158312 79694
rect 158260 79630 158312 79636
rect 158168 79620 158220 79626
rect 158168 79562 158220 79568
rect 158076 79484 158128 79490
rect 158076 79426 158128 79432
rect 157982 79248 158038 79257
rect 157982 79183 158038 79192
rect 157892 78940 157944 78946
rect 157892 78882 157944 78888
rect 157904 75682 157932 78882
rect 157996 76838 158024 79183
rect 157984 76832 158036 76838
rect 157984 76774 158036 76780
rect 158088 75886 158116 79426
rect 158076 75880 158128 75886
rect 158076 75822 158128 75828
rect 157892 75676 157944 75682
rect 157892 75618 157944 75624
rect 157904 75002 157932 75618
rect 157892 74996 157944 75002
rect 157892 74938 157944 74944
rect 158088 73710 158116 75822
rect 158076 73704 158128 73710
rect 158076 73646 158128 73652
rect 157800 73092 157852 73098
rect 157800 73034 157852 73040
rect 157708 71732 157760 71738
rect 157708 71674 157760 71680
rect 158180 70394 158208 79562
rect 158272 73794 158300 79630
rect 158536 79620 158588 79626
rect 158536 79562 158588 79568
rect 158548 78577 158576 79562
rect 158534 78568 158590 78577
rect 158534 78503 158590 78512
rect 158640 75138 158668 79766
rect 158732 79750 158806 79778
rect 158856 79792 158912 79801
rect 158732 79694 158760 79750
rect 158950 79766 159002 79772
rect 159042 79824 159094 79830
rect 159042 79766 159094 79772
rect 159180 79824 159232 79830
rect 159180 79766 159232 79772
rect 158856 79727 158912 79736
rect 158720 79688 158772 79694
rect 158720 79630 158772 79636
rect 158812 79688 158864 79694
rect 158812 79630 158864 79636
rect 159086 79656 159142 79665
rect 158718 79520 158774 79529
rect 158718 79455 158774 79464
rect 158628 75132 158680 75138
rect 158628 75074 158680 75080
rect 158628 74996 158680 75002
rect 158628 74938 158680 74944
rect 158272 73766 158576 73794
rect 158444 73704 158496 73710
rect 158444 73646 158496 73652
rect 158352 71732 158404 71738
rect 158352 71674 158404 71680
rect 157720 70366 158208 70394
rect 157720 67454 157748 70366
rect 157708 67448 157760 67454
rect 157708 67390 157760 67396
rect 157616 63368 157668 63374
rect 157616 63310 157668 63316
rect 157524 59288 157576 59294
rect 157524 59230 157576 59236
rect 157432 51060 157484 51066
rect 157432 51002 157484 51008
rect 158364 28490 158392 71674
rect 158352 28484 158404 28490
rect 158352 28426 158404 28432
rect 158456 21418 158484 73646
rect 158548 70922 158576 73766
rect 158536 70916 158588 70922
rect 158536 70858 158588 70864
rect 157984 21412 158036 21418
rect 157984 21354 158036 21360
rect 158444 21412 158496 21418
rect 158444 21354 158496 21360
rect 157340 11960 157392 11966
rect 157340 11902 157392 11908
rect 157800 8968 157852 8974
rect 157800 8910 157852 8916
rect 156604 3800 156656 3806
rect 156604 3742 156656 3748
rect 156788 3800 156840 3806
rect 156788 3742 156840 3748
rect 156616 480 156644 3742
rect 157812 480 157840 8910
rect 157996 3534 158024 21354
rect 158548 10538 158576 70858
rect 158536 10532 158588 10538
rect 158536 10474 158588 10480
rect 158640 9110 158668 74938
rect 158628 9104 158680 9110
rect 158628 9046 158680 9052
rect 158732 6526 158760 79455
rect 158824 78577 158852 79630
rect 158904 79620 158956 79626
rect 158956 79580 159036 79608
rect 159086 79591 159142 79600
rect 158904 79562 158956 79568
rect 158904 79484 158956 79490
rect 158904 79426 158956 79432
rect 158810 78568 158866 78577
rect 158916 78538 158944 79426
rect 158810 78503 158866 78512
rect 158904 78532 158956 78538
rect 158904 78474 158956 78480
rect 158812 78260 158864 78266
rect 158812 78202 158864 78208
rect 158824 56370 158852 78202
rect 158904 75404 158956 75410
rect 158904 75346 158956 75352
rect 158916 60654 158944 75346
rect 159008 64802 159036 79580
rect 159100 78742 159128 79591
rect 159088 78736 159140 78742
rect 159088 78678 159140 78684
rect 159088 75132 159140 75138
rect 159088 75074 159140 75080
rect 159100 66978 159128 75074
rect 159192 69766 159220 79766
rect 159272 79756 159324 79762
rect 159422 79744 159450 80036
rect 159514 79966 159542 80036
rect 159606 79966 159634 80036
rect 159502 79960 159554 79966
rect 159594 79960 159646 79966
rect 159502 79902 159554 79908
rect 159592 79928 159594 79937
rect 159646 79928 159648 79937
rect 159592 79863 159648 79872
rect 159548 79756 159600 79762
rect 159422 79716 159496 79744
rect 159272 79698 159324 79704
rect 159284 74458 159312 79698
rect 159468 79665 159496 79716
rect 159698 79744 159726 80036
rect 159790 79830 159818 80036
rect 159778 79824 159830 79830
rect 159778 79766 159830 79772
rect 159882 79778 159910 80036
rect 159974 79966 160002 80036
rect 159962 79960 160014 79966
rect 160066 79937 160094 80036
rect 160158 79966 160186 80036
rect 160146 79960 160198 79966
rect 159962 79902 160014 79908
rect 160052 79928 160108 79937
rect 160146 79902 160198 79908
rect 160052 79863 160108 79872
rect 159882 79750 159956 79778
rect 159548 79698 159600 79704
rect 159652 79716 159726 79744
rect 159454 79656 159510 79665
rect 159454 79591 159510 79600
rect 159560 79506 159588 79698
rect 159468 79478 159588 79506
rect 159468 75410 159496 79478
rect 159548 79416 159600 79422
rect 159548 79358 159600 79364
rect 159456 75404 159508 75410
rect 159456 75346 159508 75352
rect 159272 74452 159324 74458
rect 159272 74394 159324 74400
rect 159560 71738 159588 79358
rect 159652 75138 159680 79716
rect 159824 79688 159876 79694
rect 159824 79630 159876 79636
rect 159732 78532 159784 78538
rect 159732 78474 159784 78480
rect 159640 75132 159692 75138
rect 159640 75074 159692 75080
rect 159744 72078 159772 78474
rect 159836 78266 159864 79630
rect 159824 78260 159876 78266
rect 159824 78202 159876 78208
rect 159928 76974 159956 79750
rect 160250 79744 160278 80036
rect 160342 79812 160370 80036
rect 160434 79937 160462 80036
rect 160526 79966 160554 80036
rect 160514 79960 160566 79966
rect 160420 79928 160476 79937
rect 160514 79902 160566 79908
rect 160618 79898 160646 80036
rect 160420 79863 160476 79872
rect 160606 79892 160658 79898
rect 160606 79834 160658 79840
rect 160468 79824 160520 79830
rect 160342 79784 160416 79812
rect 160250 79716 160324 79744
rect 160100 79688 160152 79694
rect 160100 79630 160152 79636
rect 160112 78826 160140 79630
rect 160112 78798 160232 78826
rect 160100 78736 160152 78742
rect 160100 78678 160152 78684
rect 159916 76968 159968 76974
rect 159916 76910 159968 76916
rect 159916 74452 159968 74458
rect 159916 74394 159968 74400
rect 159928 74050 159956 74394
rect 159916 74044 159968 74050
rect 159916 73986 159968 73992
rect 159732 72072 159784 72078
rect 159732 72014 159784 72020
rect 159548 71732 159600 71738
rect 159548 71674 159600 71680
rect 159744 70394 159772 72014
rect 159744 70366 159864 70394
rect 159180 69760 159232 69766
rect 159180 69702 159232 69708
rect 159088 66972 159140 66978
rect 159088 66914 159140 66920
rect 159732 66972 159784 66978
rect 159732 66914 159784 66920
rect 158996 64796 159048 64802
rect 158996 64738 159048 64744
rect 158904 60648 158956 60654
rect 158904 60590 158956 60596
rect 158812 56364 158864 56370
rect 158812 56306 158864 56312
rect 159744 42294 159772 66914
rect 159732 42288 159784 42294
rect 159732 42230 159784 42236
rect 159836 32434 159864 70366
rect 159928 34066 159956 73986
rect 160112 72418 160140 78678
rect 160204 75410 160232 78798
rect 160192 75404 160244 75410
rect 160192 75346 160244 75352
rect 160192 75132 160244 75138
rect 160192 75074 160244 75080
rect 160100 72412 160152 72418
rect 160100 72354 160152 72360
rect 160100 72140 160152 72146
rect 160100 72082 160152 72088
rect 160008 71732 160060 71738
rect 160008 71674 160060 71680
rect 160020 71466 160048 71674
rect 160008 71460 160060 71466
rect 160008 71402 160060 71408
rect 159916 34060 159968 34066
rect 159916 34002 159968 34008
rect 159824 32428 159876 32434
rect 159824 32370 159876 32376
rect 160020 7886 160048 71402
rect 160112 10470 160140 72082
rect 160204 57866 160232 75074
rect 160296 65822 160324 79716
rect 160388 69018 160416 79784
rect 160468 79766 160520 79772
rect 160480 77858 160508 79766
rect 160560 79756 160612 79762
rect 160560 79698 160612 79704
rect 160468 77852 160520 77858
rect 160468 77794 160520 77800
rect 160572 75138 160600 79698
rect 160710 79676 160738 80036
rect 160802 79898 160830 80036
rect 160894 79937 160922 80036
rect 160880 79928 160936 79937
rect 160790 79892 160842 79898
rect 160880 79863 160936 79872
rect 160790 79834 160842 79840
rect 160986 79801 161014 80036
rect 161078 79898 161106 80036
rect 161066 79892 161118 79898
rect 161066 79834 161118 79840
rect 160834 79792 160890 79801
rect 160834 79727 160890 79736
rect 160972 79792 161028 79801
rect 161170 79744 161198 80036
rect 160972 79727 161028 79736
rect 160664 79648 160738 79676
rect 160664 75138 160692 79648
rect 160848 79608 160876 79727
rect 161124 79716 161198 79744
rect 161262 79744 161290 80036
rect 161354 79898 161382 80036
rect 161342 79892 161394 79898
rect 161342 79834 161394 79840
rect 161446 79744 161474 80036
rect 161262 79716 161336 79744
rect 161020 79620 161072 79626
rect 160848 79580 160968 79608
rect 160834 79520 160890 79529
rect 160834 79455 160890 79464
rect 160744 79416 160796 79422
rect 160744 79358 160796 79364
rect 160756 76906 160784 79358
rect 160848 77081 160876 79455
rect 160834 77072 160890 77081
rect 160834 77007 160890 77016
rect 160744 76900 160796 76906
rect 160744 76842 160796 76848
rect 160756 75954 160784 76842
rect 160940 76616 160968 79580
rect 161020 79562 161072 79568
rect 161032 78402 161060 79562
rect 161020 78396 161072 78402
rect 161020 78338 161072 78344
rect 161124 77489 161152 79716
rect 161204 79620 161256 79626
rect 161204 79562 161256 79568
rect 161216 78946 161244 79562
rect 161204 78940 161256 78946
rect 161204 78882 161256 78888
rect 161110 77480 161166 77489
rect 161110 77415 161166 77424
rect 161216 77330 161244 78882
rect 161124 77302 161244 77330
rect 160940 76588 161060 76616
rect 160744 75948 160796 75954
rect 160744 75890 160796 75896
rect 160928 75404 160980 75410
rect 160928 75346 160980 75352
rect 160560 75132 160612 75138
rect 160560 75074 160612 75080
rect 160652 75132 160704 75138
rect 160652 75074 160704 75080
rect 160940 71194 160968 75346
rect 161032 71262 161060 76588
rect 161124 72146 161152 77302
rect 161204 75132 161256 75138
rect 161204 75074 161256 75080
rect 161216 74934 161244 75074
rect 161204 74928 161256 74934
rect 161204 74870 161256 74876
rect 161112 72140 161164 72146
rect 161112 72082 161164 72088
rect 161020 71256 161072 71262
rect 161020 71198 161072 71204
rect 160928 71188 160980 71194
rect 160928 71130 160980 71136
rect 160376 69012 160428 69018
rect 160376 68954 160428 68960
rect 160284 65816 160336 65822
rect 160284 65758 160336 65764
rect 160192 57860 160244 57866
rect 160192 57802 160244 57808
rect 160940 31142 160968 71130
rect 161032 70394 161060 71198
rect 161032 70366 161152 70394
rect 161020 65816 161072 65822
rect 161020 65758 161072 65764
rect 160928 31136 160980 31142
rect 160928 31078 160980 31084
rect 161032 19990 161060 65758
rect 161020 19984 161072 19990
rect 161020 19926 161072 19932
rect 161124 16114 161152 70366
rect 161112 16108 161164 16114
rect 161112 16050 161164 16056
rect 161216 16046 161244 74870
rect 161308 73030 161336 79716
rect 161400 79716 161474 79744
rect 161538 79744 161566 80036
rect 161630 79898 161658 80036
rect 161722 79898 161750 80036
rect 161618 79892 161670 79898
rect 161618 79834 161670 79840
rect 161710 79892 161762 79898
rect 161710 79834 161762 79840
rect 161814 79744 161842 80036
rect 161538 79716 161612 79744
rect 161400 78577 161428 79716
rect 161480 79620 161532 79626
rect 161480 79562 161532 79568
rect 161386 78568 161442 78577
rect 161386 78503 161442 78512
rect 161492 77382 161520 79562
rect 161480 77376 161532 77382
rect 161480 77318 161532 77324
rect 161388 75948 161440 75954
rect 161388 75890 161440 75896
rect 161296 73024 161348 73030
rect 161296 72966 161348 72972
rect 161204 16040 161256 16046
rect 161204 15982 161256 15988
rect 161110 15872 161166 15881
rect 161110 15807 161166 15816
rect 160100 10464 160152 10470
rect 160100 10406 160152 10412
rect 160008 7880 160060 7886
rect 160008 7822 160060 7828
rect 160098 7576 160154 7585
rect 160098 7511 160154 7520
rect 158720 6520 158772 6526
rect 158720 6462 158772 6468
rect 157984 3528 158036 3534
rect 157984 3470 158036 3476
rect 158904 3528 158956 3534
rect 158904 3470 158956 3476
rect 158916 480 158944 3470
rect 160112 480 160140 7511
rect 161124 3482 161152 15807
rect 161308 6914 161336 72966
rect 161400 7818 161428 75890
rect 161480 75540 161532 75546
rect 161480 75482 161532 75488
rect 161492 67561 161520 75482
rect 161584 69970 161612 79716
rect 161676 79716 161842 79744
rect 161572 69964 161624 69970
rect 161572 69906 161624 69912
rect 161676 69834 161704 79716
rect 161906 79676 161934 80036
rect 161998 79966 162026 80036
rect 162090 79966 162118 80036
rect 162182 79966 162210 80036
rect 162274 79971 162302 80036
rect 161986 79960 162038 79966
rect 161986 79902 162038 79908
rect 162078 79960 162130 79966
rect 162078 79902 162130 79908
rect 162170 79960 162222 79966
rect 162170 79902 162222 79908
rect 162260 79962 162316 79971
rect 162366 79966 162394 80036
rect 162458 79966 162486 80036
rect 162550 79966 162578 80036
rect 162642 79971 162670 80036
rect 162260 79897 162316 79906
rect 162354 79960 162406 79966
rect 162354 79902 162406 79908
rect 162446 79960 162498 79966
rect 162446 79902 162498 79908
rect 162538 79960 162590 79966
rect 162538 79902 162590 79908
rect 162628 79962 162684 79971
rect 162734 79966 162762 80036
rect 162628 79897 162684 79906
rect 162722 79960 162774 79966
rect 162722 79902 162774 79908
rect 162032 79824 162084 79830
rect 162032 79766 162084 79772
rect 162308 79824 162360 79830
rect 162446 79824 162498 79830
rect 162308 79766 162360 79772
rect 162412 79772 162446 79778
rect 162826 79812 162854 80036
rect 162412 79766 162498 79772
rect 162780 79784 162854 79812
rect 161768 79648 161934 79676
rect 161664 69828 161716 69834
rect 161664 69770 161716 69776
rect 161768 69494 161796 79648
rect 161848 79552 161900 79558
rect 161848 79494 161900 79500
rect 161860 77518 161888 79494
rect 161940 79484 161992 79490
rect 161940 79426 161992 79432
rect 161952 79150 161980 79426
rect 161940 79144 161992 79150
rect 161940 79086 161992 79092
rect 161848 77512 161900 77518
rect 161848 77454 161900 77460
rect 161848 77376 161900 77382
rect 161848 77318 161900 77324
rect 161860 74458 161888 77318
rect 161848 74452 161900 74458
rect 161848 74394 161900 74400
rect 162044 70394 162072 79766
rect 162124 79756 162176 79762
rect 162124 79698 162176 79704
rect 162136 77976 162164 79698
rect 162136 77948 162256 77976
rect 162124 77852 162176 77858
rect 162124 77794 162176 77800
rect 161860 70366 162072 70394
rect 161860 69630 161888 70366
rect 161848 69624 161900 69630
rect 161848 69566 161900 69572
rect 161756 69488 161808 69494
rect 161756 69430 161808 69436
rect 161478 67552 161534 67561
rect 161478 67487 161534 67496
rect 162136 66842 162164 77794
rect 162228 72350 162256 77948
rect 162320 74866 162348 79766
rect 162412 79750 162486 79766
rect 162412 75546 162440 79750
rect 162492 79688 162544 79694
rect 162490 79656 162492 79665
rect 162544 79656 162546 79665
rect 162490 79591 162546 79600
rect 162676 79620 162728 79626
rect 162676 79562 162728 79568
rect 162492 79552 162544 79558
rect 162492 79494 162544 79500
rect 162504 77722 162532 79494
rect 162582 79248 162638 79257
rect 162582 79183 162638 79192
rect 162596 78742 162624 79183
rect 162584 78736 162636 78742
rect 162584 78678 162636 78684
rect 162492 77716 162544 77722
rect 162492 77658 162544 77664
rect 162584 77580 162636 77586
rect 162584 77522 162636 77528
rect 162400 75540 162452 75546
rect 162400 75482 162452 75488
rect 162308 74860 162360 74866
rect 162308 74802 162360 74808
rect 162216 72344 162268 72350
rect 162216 72286 162268 72292
rect 162400 70236 162452 70242
rect 162400 70178 162452 70184
rect 162308 70168 162360 70174
rect 162308 70110 162360 70116
rect 162320 69970 162348 70110
rect 162308 69964 162360 69970
rect 162308 69906 162360 69912
rect 162124 66836 162176 66842
rect 162124 66778 162176 66784
rect 162136 64874 162164 66778
rect 162136 64846 162256 64874
rect 162228 36786 162256 64846
rect 162216 36780 162268 36786
rect 162216 36722 162268 36728
rect 162320 27130 162348 69906
rect 162412 69834 162440 70178
rect 162596 69834 162624 77522
rect 162688 76537 162716 79562
rect 162780 77217 162808 79784
rect 162918 79744 162946 80036
rect 163010 79830 163038 80036
rect 163102 79966 163130 80036
rect 163090 79960 163142 79966
rect 163090 79902 163142 79908
rect 162998 79824 163050 79830
rect 163194 79812 163222 80036
rect 163286 79966 163314 80036
rect 163378 79966 163406 80036
rect 163470 79966 163498 80036
rect 163274 79960 163326 79966
rect 163274 79902 163326 79908
rect 163366 79960 163418 79966
rect 163366 79902 163418 79908
rect 163458 79960 163510 79966
rect 163458 79902 163510 79908
rect 163194 79784 163268 79812
rect 162998 79766 163050 79772
rect 163240 79778 163268 79784
rect 163240 79750 163452 79778
rect 162872 79716 162946 79744
rect 162872 79665 162900 79716
rect 163136 79688 163188 79694
rect 162858 79656 162914 79665
rect 163136 79630 163188 79636
rect 163228 79688 163280 79694
rect 163228 79630 163280 79636
rect 163320 79688 163372 79694
rect 163320 79630 163372 79636
rect 162858 79591 162914 79600
rect 163044 79620 163096 79626
rect 163044 79562 163096 79568
rect 162860 79552 162912 79558
rect 162860 79494 162912 79500
rect 162872 79082 162900 79494
rect 162950 79248 163006 79257
rect 162950 79183 163006 79192
rect 162860 79076 162912 79082
rect 162860 79018 162912 79024
rect 162766 77208 162822 77217
rect 162766 77143 162822 77152
rect 162674 76528 162730 76537
rect 162674 76463 162730 76472
rect 162676 74860 162728 74866
rect 162676 74802 162728 74808
rect 162688 72690 162716 74802
rect 162676 72684 162728 72690
rect 162676 72626 162728 72632
rect 162400 69828 162452 69834
rect 162400 69770 162452 69776
rect 162584 69828 162636 69834
rect 162584 69770 162636 69776
rect 162308 27124 162360 27130
rect 162308 27066 162360 27072
rect 162412 25770 162440 69770
rect 162584 69624 162636 69630
rect 162584 69566 162636 69572
rect 162490 67552 162546 67561
rect 162490 67487 162546 67496
rect 162400 25764 162452 25770
rect 162400 25706 162452 25712
rect 162504 13190 162532 67487
rect 162596 13258 162624 69566
rect 162688 14618 162716 72626
rect 162768 69488 162820 69494
rect 162768 69430 162820 69436
rect 162676 14612 162728 14618
rect 162676 14554 162728 14560
rect 162584 13252 162636 13258
rect 162584 13194 162636 13200
rect 162492 13184 162544 13190
rect 162492 13126 162544 13132
rect 162780 11898 162808 69430
rect 162872 22982 162900 79018
rect 162964 29782 162992 79183
rect 163056 78470 163084 79562
rect 163044 78464 163096 78470
rect 163044 78406 163096 78412
rect 163044 78124 163096 78130
rect 163044 78066 163096 78072
rect 163056 73982 163084 78066
rect 163148 75936 163176 79630
rect 163240 76158 163268 79630
rect 163228 76152 163280 76158
rect 163228 76094 163280 76100
rect 163148 75908 163268 75936
rect 163136 75812 163188 75818
rect 163136 75754 163188 75760
rect 163044 73976 163096 73982
rect 163044 73918 163096 73924
rect 163044 73772 163096 73778
rect 163044 73714 163096 73720
rect 163056 43518 163084 73714
rect 163148 56438 163176 75754
rect 163240 62014 163268 75908
rect 163332 75818 163360 79630
rect 163424 79014 163452 79750
rect 163562 79744 163590 80036
rect 163654 79971 163682 80036
rect 163640 79962 163696 79971
rect 163640 79897 163696 79906
rect 163746 79898 163774 80036
rect 163734 79892 163786 79898
rect 163734 79834 163786 79840
rect 163838 79778 163866 80036
rect 163930 79812 163958 80036
rect 164022 79937 164050 80036
rect 164008 79928 164064 79937
rect 164008 79863 164064 79872
rect 164114 79830 164142 80036
rect 164102 79824 164154 79830
rect 163930 79784 164004 79812
rect 163746 79750 163866 79778
rect 163562 79716 163636 79744
rect 163502 79656 163558 79665
rect 163502 79591 163558 79600
rect 163412 79008 163464 79014
rect 163412 78950 163464 78956
rect 163412 76152 163464 76158
rect 163412 76094 163464 76100
rect 163320 75812 163372 75818
rect 163320 75754 163372 75760
rect 163320 75608 163372 75614
rect 163320 75550 163372 75556
rect 163332 66230 163360 75550
rect 163424 67590 163452 76094
rect 163516 69630 163544 79591
rect 163608 78130 163636 79716
rect 163746 79676 163774 79750
rect 163976 79676 164004 79784
rect 164102 79766 164154 79772
rect 164206 79744 164234 80036
rect 164298 79971 164326 80036
rect 164284 79962 164340 79971
rect 164390 79966 164418 80036
rect 164482 79971 164510 80036
rect 164284 79897 164340 79906
rect 164378 79960 164430 79966
rect 164378 79902 164430 79908
rect 164468 79962 164524 79971
rect 164574 79966 164602 80036
rect 164468 79897 164524 79906
rect 164562 79960 164614 79966
rect 164562 79902 164614 79908
rect 164666 79898 164694 80036
rect 164654 79892 164706 79898
rect 164654 79834 164706 79840
rect 164516 79756 164568 79762
rect 164206 79716 164280 79744
rect 164252 79676 164280 79716
rect 164516 79698 164568 79704
rect 164608 79756 164660 79762
rect 164758 79744 164786 80036
rect 164850 79812 164878 80036
rect 164942 79937 164970 80036
rect 165034 79966 165062 80036
rect 165022 79960 165074 79966
rect 164928 79928 164984 79937
rect 165022 79902 165074 79908
rect 164928 79863 164984 79872
rect 164850 79784 165016 79812
rect 164758 79716 164832 79744
rect 164608 79698 164660 79704
rect 163746 79648 163820 79676
rect 163686 79520 163742 79529
rect 163686 79455 163742 79464
rect 163596 78124 163648 78130
rect 163596 78066 163648 78072
rect 163700 76430 163728 79455
rect 163688 76424 163740 76430
rect 163688 76366 163740 76372
rect 163792 75614 163820 79648
rect 163884 79648 164004 79676
rect 164160 79648 164280 79676
rect 164332 79688 164384 79694
rect 163884 75993 163912 79648
rect 164056 79620 164108 79626
rect 164056 79562 164108 79568
rect 163870 75984 163926 75993
rect 163870 75919 163926 75928
rect 163780 75608 163832 75614
rect 163780 75550 163832 75556
rect 164068 73642 164096 79562
rect 164160 79121 164188 79648
rect 164332 79630 164384 79636
rect 164146 79112 164202 79121
rect 164146 79047 164202 79056
rect 164160 73778 164188 79047
rect 164344 77994 164372 79630
rect 164424 79416 164476 79422
rect 164424 79358 164476 79364
rect 164332 77988 164384 77994
rect 164332 77930 164384 77936
rect 164240 77308 164292 77314
rect 164240 77250 164292 77256
rect 164148 73772 164200 73778
rect 164148 73714 164200 73720
rect 164056 73636 164108 73642
rect 164056 73578 164108 73584
rect 163504 69624 163556 69630
rect 163504 69566 163556 69572
rect 163964 69624 164016 69630
rect 163964 69566 164016 69572
rect 163412 67584 163464 67590
rect 163412 67526 163464 67532
rect 163320 66224 163372 66230
rect 163320 66166 163372 66172
rect 163228 62008 163280 62014
rect 163228 61950 163280 61956
rect 163136 56432 163188 56438
rect 163136 56374 163188 56380
rect 163044 43512 163096 43518
rect 163044 43454 163096 43460
rect 162952 29776 163004 29782
rect 162952 29718 163004 29724
rect 163976 24274 164004 69566
rect 164148 67584 164200 67590
rect 164148 67526 164200 67532
rect 164056 66224 164108 66230
rect 164056 66166 164108 66172
rect 164068 65890 164096 66166
rect 164056 65884 164108 65890
rect 164056 65826 164108 65832
rect 163964 24268 164016 24274
rect 163964 24210 164016 24216
rect 162860 22976 162912 22982
rect 162860 22918 162912 22924
rect 164068 14550 164096 65826
rect 164056 14544 164108 14550
rect 164056 14486 164108 14492
rect 162768 11892 162820 11898
rect 162768 11834 162820 11840
rect 161388 7812 161440 7818
rect 161388 7754 161440 7760
rect 161216 6886 161336 6914
rect 161216 5030 161244 6886
rect 161204 5024 161256 5030
rect 161204 4966 161256 4972
rect 164160 4962 164188 67526
rect 164252 42226 164280 77250
rect 164332 77036 164384 77042
rect 164332 76978 164384 76984
rect 164344 55214 164372 76978
rect 164436 66094 164464 79358
rect 164528 67590 164556 79698
rect 164620 76974 164648 79698
rect 164698 78160 164754 78169
rect 164698 78095 164754 78104
rect 164608 76968 164660 76974
rect 164608 76910 164660 76916
rect 164712 76786 164740 78095
rect 164804 77042 164832 79716
rect 164884 79688 164936 79694
rect 164884 79630 164936 79636
rect 164896 79150 164924 79630
rect 164884 79144 164936 79150
rect 164884 79086 164936 79092
rect 164792 77036 164844 77042
rect 164792 76978 164844 76984
rect 164790 76936 164846 76945
rect 164790 76871 164846 76880
rect 164620 76758 164740 76786
rect 164620 70106 164648 76758
rect 164804 76616 164832 76871
rect 164712 76588 164832 76616
rect 164608 70100 164660 70106
rect 164608 70042 164660 70048
rect 164516 67584 164568 67590
rect 164516 67526 164568 67532
rect 164424 66088 164476 66094
rect 164424 66030 164476 66036
rect 164620 64874 164648 70042
rect 164712 70009 164740 76588
rect 164792 75948 164844 75954
rect 164792 75890 164844 75896
rect 164804 70038 164832 75890
rect 164988 73154 165016 79784
rect 165126 79744 165154 80036
rect 165218 79898 165246 80036
rect 165206 79892 165258 79898
rect 165206 79834 165258 79840
rect 165310 79830 165338 80036
rect 165402 79830 165430 80036
rect 165298 79824 165350 79830
rect 165298 79766 165350 79772
rect 165390 79824 165442 79830
rect 165494 79812 165522 80036
rect 165586 79966 165614 80036
rect 165574 79960 165626 79966
rect 165678 79937 165706 80036
rect 165770 79966 165798 80036
rect 165758 79960 165810 79966
rect 165574 79902 165626 79908
rect 165664 79928 165720 79937
rect 165862 79937 165890 80036
rect 165954 79966 165982 80036
rect 166046 79966 166074 80036
rect 166138 79971 166166 80036
rect 165942 79960 165994 79966
rect 165758 79902 165810 79908
rect 165848 79928 165904 79937
rect 165664 79863 165720 79872
rect 165942 79902 165994 79908
rect 166034 79960 166086 79966
rect 166034 79902 166086 79908
rect 166124 79962 166180 79971
rect 166124 79897 166180 79906
rect 165848 79863 165904 79872
rect 166034 79824 166086 79830
rect 165494 79784 165660 79812
rect 165390 79766 165442 79772
rect 165080 79716 165154 79744
rect 165080 75954 165108 79716
rect 165436 79688 165488 79694
rect 165436 79630 165488 79636
rect 165528 79688 165580 79694
rect 165528 79630 165580 79636
rect 165344 79620 165396 79626
rect 165344 79562 165396 79568
rect 165252 79008 165304 79014
rect 165252 78950 165304 78956
rect 165068 75948 165120 75954
rect 165068 75890 165120 75896
rect 164896 73126 165016 73154
rect 164792 70032 164844 70038
rect 164698 70000 164754 70009
rect 164792 69974 164844 69980
rect 164896 69970 164924 73126
rect 165264 70394 165292 78950
rect 165356 75993 165384 79562
rect 165448 78985 165476 79630
rect 165540 79257 165568 79630
rect 165526 79248 165582 79257
rect 165526 79183 165582 79192
rect 165434 78976 165490 78985
rect 165434 78911 165490 78920
rect 165436 78600 165488 78606
rect 165436 78542 165488 78548
rect 165448 78198 165476 78542
rect 165436 78192 165488 78198
rect 165436 78134 165488 78140
rect 165540 77314 165568 79183
rect 165632 78305 165660 79784
rect 165908 79784 166034 79812
rect 165804 79756 165856 79762
rect 165804 79698 165856 79704
rect 165618 78296 165674 78305
rect 165618 78231 165674 78240
rect 165816 77586 165844 79698
rect 165804 77580 165856 77586
rect 165804 77522 165856 77528
rect 165528 77308 165580 77314
rect 165908 77294 165936 79784
rect 166034 79766 166086 79772
rect 166230 79744 166258 80036
rect 166322 79966 166350 80036
rect 166414 79966 166442 80036
rect 166506 79966 166534 80036
rect 166310 79960 166362 79966
rect 166310 79902 166362 79908
rect 166402 79960 166454 79966
rect 166402 79902 166454 79908
rect 166494 79960 166546 79966
rect 166494 79902 166546 79908
rect 166598 79801 166626 80036
rect 166584 79792 166640 79801
rect 166230 79716 166304 79744
rect 166584 79727 166640 79736
rect 166690 79744 166718 80036
rect 166782 79812 166810 80036
rect 166874 79966 166902 80036
rect 166862 79960 166914 79966
rect 166862 79902 166914 79908
rect 166782 79784 166856 79812
rect 166966 79801 166994 80036
rect 167058 79966 167086 80036
rect 167046 79960 167098 79966
rect 167046 79902 167098 79908
rect 167150 79812 167178 80036
rect 167242 79903 167270 80036
rect 167228 79894 167284 79903
rect 167228 79829 167284 79838
rect 166690 79716 166764 79744
rect 166080 79620 166132 79626
rect 166080 79562 166132 79568
rect 166172 79620 166224 79626
rect 166172 79562 166224 79568
rect 165988 78668 166040 78674
rect 165988 78610 166040 78616
rect 165528 77250 165580 77256
rect 165724 77266 165936 77294
rect 165528 76968 165580 76974
rect 165528 76910 165580 76916
rect 165342 75984 165398 75993
rect 165342 75919 165398 75928
rect 165540 70854 165568 76910
rect 165724 76072 165752 77266
rect 166000 76106 166028 78610
rect 165632 76044 165752 76072
rect 165908 76078 166028 76106
rect 165528 70848 165580 70854
rect 165528 70790 165580 70796
rect 165264 70366 165384 70394
rect 165252 70304 165304 70310
rect 165252 70246 165304 70252
rect 165264 70038 165292 70246
rect 165252 70032 165304 70038
rect 165252 69974 165304 69980
rect 164698 69935 164754 69944
rect 164884 69964 164936 69970
rect 164712 68218 164740 69935
rect 164884 69906 164936 69912
rect 165264 68354 165292 69974
rect 165356 68474 165384 70366
rect 165436 69964 165488 69970
rect 165436 69906 165488 69912
rect 165344 68468 165396 68474
rect 165344 68410 165396 68416
rect 165264 68326 165384 68354
rect 164712 68190 165292 68218
rect 165160 67584 165212 67590
rect 165160 67526 165212 67532
rect 165172 67386 165200 67526
rect 165160 67380 165212 67386
rect 165160 67322 165212 67328
rect 164620 64846 165108 64874
rect 164332 55208 164384 55214
rect 164332 55150 164384 55156
rect 164240 42220 164292 42226
rect 164240 42162 164292 42168
rect 165080 39574 165108 64846
rect 165068 39568 165120 39574
rect 165068 39510 165120 39516
rect 165172 27062 165200 67322
rect 165160 27056 165212 27062
rect 165160 26998 165212 27004
rect 165264 25702 165292 68190
rect 165252 25696 165304 25702
rect 165252 25638 165304 25644
rect 165356 15978 165384 68326
rect 165344 15972 165396 15978
rect 165344 15914 165396 15920
rect 165448 11830 165476 69906
rect 165436 11824 165488 11830
rect 165436 11766 165488 11772
rect 165540 9042 165568 70790
rect 165632 67318 165660 76044
rect 165802 75984 165858 75993
rect 165802 75919 165858 75928
rect 165712 74588 165764 74594
rect 165712 74530 165764 74536
rect 165724 68746 165752 74530
rect 165816 68814 165844 75919
rect 165804 68808 165856 68814
rect 165804 68750 165856 68756
rect 165712 68740 165764 68746
rect 165712 68682 165764 68688
rect 165908 68406 165936 76078
rect 165988 76016 166040 76022
rect 165988 75958 166040 75964
rect 166000 68882 166028 75958
rect 166092 68950 166120 79562
rect 166184 74594 166212 79562
rect 166172 74588 166224 74594
rect 166172 74530 166224 74536
rect 166276 74322 166304 79716
rect 166448 79688 166500 79694
rect 166448 79630 166500 79636
rect 166538 79656 166594 79665
rect 166356 79552 166408 79558
rect 166356 79494 166408 79500
rect 166368 77790 166396 79494
rect 166460 78198 166488 79630
rect 166538 79591 166594 79600
rect 166632 79620 166684 79626
rect 166448 78192 166500 78198
rect 166448 78134 166500 78140
rect 166356 77784 166408 77790
rect 166356 77726 166408 77732
rect 166264 74316 166316 74322
rect 166264 74258 166316 74264
rect 166264 73636 166316 73642
rect 166264 73578 166316 73584
rect 166172 69964 166224 69970
rect 166172 69906 166224 69912
rect 166184 69562 166212 69906
rect 166172 69556 166224 69562
rect 166172 69498 166224 69504
rect 166080 68944 166132 68950
rect 166080 68886 166132 68892
rect 165988 68876 166040 68882
rect 165988 68818 166040 68824
rect 165896 68400 165948 68406
rect 165896 68342 165948 68348
rect 165620 67312 165672 67318
rect 165620 67254 165672 67260
rect 166000 66910 166028 68818
rect 166172 67516 166224 67522
rect 166172 67458 166224 67464
rect 166184 67318 166212 67458
rect 166172 67312 166224 67318
rect 166172 67254 166224 67260
rect 165988 66904 166040 66910
rect 165988 66846 166040 66852
rect 166184 18766 166212 67254
rect 166276 53718 166304 73578
rect 166552 72894 166580 79591
rect 166632 79562 166684 79568
rect 166644 78577 166672 79562
rect 166736 78674 166764 79716
rect 166724 78668 166776 78674
rect 166724 78610 166776 78616
rect 166630 78568 166686 78577
rect 166630 78503 166686 78512
rect 166828 77294 166856 79784
rect 166952 79792 167008 79801
rect 166952 79727 167008 79736
rect 167104 79784 167178 79812
rect 167000 79688 167052 79694
rect 167000 79630 167052 79636
rect 166908 79620 166960 79626
rect 166908 79562 166960 79568
rect 166920 77926 166948 79562
rect 167012 78577 167040 79630
rect 167104 79558 167132 79784
rect 167334 79778 167362 80036
rect 167426 79966 167454 80036
rect 167518 79966 167546 80036
rect 167414 79960 167466 79966
rect 167414 79902 167466 79908
rect 167506 79960 167558 79966
rect 167506 79902 167558 79908
rect 167610 79812 167638 80036
rect 167702 79971 167730 80036
rect 167688 79962 167744 79971
rect 167688 79897 167744 79906
rect 167610 79784 167684 79812
rect 167334 79750 167408 79778
rect 167274 79656 167330 79665
rect 167196 79614 167274 79642
rect 167092 79552 167144 79558
rect 167092 79494 167144 79500
rect 167092 79416 167144 79422
rect 167092 79358 167144 79364
rect 166998 78568 167054 78577
rect 166998 78503 167054 78512
rect 166908 77920 166960 77926
rect 166908 77862 166960 77868
rect 166908 77512 166960 77518
rect 166908 77454 166960 77460
rect 166736 77266 166856 77294
rect 166736 76022 166764 77266
rect 166920 77194 166948 77454
rect 166828 77166 166948 77194
rect 166724 76016 166776 76022
rect 166724 75958 166776 75964
rect 166724 75064 166776 75070
rect 166724 75006 166776 75012
rect 166736 74730 166764 75006
rect 166724 74724 166776 74730
rect 166724 74666 166776 74672
rect 166540 72888 166592 72894
rect 166540 72830 166592 72836
rect 166552 71774 166580 72830
rect 166552 71746 166672 71774
rect 166448 68808 166500 68814
rect 166448 68750 166500 68756
rect 166356 68740 166408 68746
rect 166356 68682 166408 68688
rect 166368 68066 166396 68682
rect 166460 68134 166488 68750
rect 166448 68128 166500 68134
rect 166448 68070 166500 68076
rect 166356 68060 166408 68066
rect 166356 68002 166408 68008
rect 166264 53712 166316 53718
rect 166264 53654 166316 53660
rect 166368 42158 166396 68002
rect 166356 42152 166408 42158
rect 166356 42094 166408 42100
rect 166460 28422 166488 68070
rect 166448 28416 166500 28422
rect 166448 28358 166500 28364
rect 166644 22914 166672 71746
rect 166828 70394 166856 77166
rect 166998 75984 167054 75993
rect 166998 75919 167054 75928
rect 166908 74316 166960 74322
rect 166908 74258 166960 74264
rect 166736 70366 166856 70394
rect 166736 67250 166764 70366
rect 166816 68944 166868 68950
rect 166816 68886 166868 68892
rect 166828 68678 166856 68886
rect 166816 68672 166868 68678
rect 166816 68614 166868 68620
rect 166724 67244 166776 67250
rect 166724 67186 166776 67192
rect 166828 67130 166856 68614
rect 166736 67102 166856 67130
rect 166632 22908 166684 22914
rect 166632 22850 166684 22856
rect 166172 18760 166224 18766
rect 166172 18702 166224 18708
rect 166736 10402 166764 67102
rect 166816 66904 166868 66910
rect 166816 66846 166868 66852
rect 166724 10396 166776 10402
rect 166724 10338 166776 10344
rect 165528 9036 165580 9042
rect 165528 8978 165580 8984
rect 166828 7682 166856 66846
rect 166920 7750 166948 74258
rect 167012 56506 167040 75919
rect 167000 56500 167052 56506
rect 167000 56442 167052 56448
rect 167000 42084 167052 42090
rect 167000 42026 167052 42032
rect 167012 16574 167040 42026
rect 167104 40866 167132 79358
rect 167196 59362 167224 79614
rect 167274 79591 167330 79600
rect 167274 79384 167330 79393
rect 167274 79319 167330 79328
rect 167184 59356 167236 59362
rect 167184 59298 167236 59304
rect 167288 43450 167316 79319
rect 167380 78441 167408 79750
rect 167552 79484 167604 79490
rect 167552 79426 167604 79432
rect 167460 78464 167512 78470
rect 167366 78432 167422 78441
rect 167460 78406 167512 78412
rect 167366 78367 167422 78376
rect 167472 77586 167500 78406
rect 167460 77580 167512 77586
rect 167460 77522 167512 77528
rect 167460 76968 167512 76974
rect 167460 76910 167512 76916
rect 167472 75936 167500 76910
rect 167380 75908 167500 75936
rect 167380 60586 167408 75908
rect 167564 71774 167592 79426
rect 167656 73166 167684 79784
rect 167794 79744 167822 80036
rect 167886 79801 167914 80036
rect 167978 79898 168006 80036
rect 168070 79937 168098 80036
rect 168056 79928 168112 79937
rect 167966 79892 168018 79898
rect 168162 79898 168190 80036
rect 168056 79863 168112 79872
rect 168150 79892 168202 79898
rect 167966 79834 168018 79840
rect 168150 79834 168202 79840
rect 168254 79812 168282 80036
rect 168346 79966 168374 80036
rect 168438 79966 168466 80036
rect 168334 79960 168386 79966
rect 168334 79902 168386 79908
rect 168426 79960 168478 79966
rect 168426 79902 168478 79908
rect 168530 79898 168558 80036
rect 168622 79937 168650 80036
rect 168714 79966 168742 80036
rect 168806 79971 168834 80036
rect 168702 79960 168754 79966
rect 168608 79928 168664 79937
rect 168518 79892 168570 79898
rect 168702 79902 168754 79908
rect 168792 79962 168848 79971
rect 168792 79897 168848 79906
rect 168898 79898 168926 80036
rect 168990 79966 169018 80036
rect 169082 79966 169110 80036
rect 169174 79966 169202 80036
rect 168978 79960 169030 79966
rect 168978 79902 169030 79908
rect 169070 79960 169122 79966
rect 169070 79902 169122 79908
rect 169162 79960 169214 79966
rect 169162 79902 169214 79908
rect 169266 79898 169294 80036
rect 168608 79863 168664 79872
rect 168886 79892 168938 79898
rect 168518 79834 168570 79840
rect 168886 79834 168938 79840
rect 169254 79892 169306 79898
rect 169254 79834 169306 79840
rect 168656 79824 168708 79830
rect 167748 79716 167822 79744
rect 167872 79792 167928 79801
rect 168254 79784 168328 79812
rect 167872 79727 167928 79736
rect 168104 79756 168156 79762
rect 167748 75993 167776 79716
rect 168104 79698 168156 79704
rect 168012 79688 168064 79694
rect 168012 79630 168064 79636
rect 167920 79552 167972 79558
rect 167920 79494 167972 79500
rect 167932 78266 167960 79494
rect 168024 78742 168052 79630
rect 168012 78736 168064 78742
rect 168012 78678 168064 78684
rect 168116 78470 168144 79698
rect 168196 79688 168248 79694
rect 168196 79630 168248 79636
rect 168104 78464 168156 78470
rect 168104 78406 168156 78412
rect 168012 78396 168064 78402
rect 168012 78338 168064 78344
rect 167920 78260 167972 78266
rect 167920 78202 167972 78208
rect 167734 75984 167790 75993
rect 167734 75919 167790 75928
rect 167644 73160 167696 73166
rect 167644 73102 167696 73108
rect 167472 71746 167592 71774
rect 167472 62966 167500 71746
rect 168024 70394 168052 78338
rect 168208 76974 168236 79630
rect 168196 76968 168248 76974
rect 168196 76910 168248 76916
rect 168196 76832 168248 76838
rect 168196 76774 168248 76780
rect 168024 70378 168144 70394
rect 168024 70372 168156 70378
rect 168024 70366 168104 70372
rect 168104 70314 168156 70320
rect 168104 63300 168156 63306
rect 168104 63242 168156 63248
rect 168116 62966 168144 63242
rect 167460 62960 167512 62966
rect 167460 62902 167512 62908
rect 168104 62960 168156 62966
rect 168104 62902 168156 62908
rect 167368 60580 167420 60586
rect 167368 60522 167420 60528
rect 167644 50380 167696 50386
rect 167644 50322 167696 50328
rect 167276 43444 167328 43450
rect 167276 43386 167328 43392
rect 167092 40860 167144 40866
rect 167092 40802 167144 40808
rect 167012 16546 167224 16574
rect 166908 7744 166960 7750
rect 166908 7686 166960 7692
rect 166816 7676 166868 7682
rect 166816 7618 166868 7624
rect 164148 4956 164200 4962
rect 164148 4898 164200 4904
rect 164884 3868 164936 3874
rect 164884 3810 164936 3816
rect 163688 3732 163740 3738
rect 163688 3674 163740 3680
rect 162492 3664 162544 3670
rect 162492 3606 162544 3612
rect 161124 3454 161336 3482
rect 161308 480 161336 3454
rect 162504 480 162532 3606
rect 163700 480 163728 3674
rect 164896 480 164924 3810
rect 166080 3596 166132 3602
rect 166080 3538 166132 3544
rect 166092 480 166120 3538
rect 167196 480 167224 16546
rect 167656 3466 167684 50322
rect 168116 33998 168144 62902
rect 168104 33992 168156 33998
rect 168104 33934 168156 33940
rect 168208 17406 168236 76774
rect 168300 73642 168328 79784
rect 168378 79792 168434 79801
rect 168378 79727 168434 79736
rect 168562 79792 168618 79801
rect 168656 79766 168708 79772
rect 168748 79824 168800 79830
rect 169358 79812 169386 80036
rect 169450 79937 169478 80036
rect 169542 79966 169570 80036
rect 169530 79960 169582 79966
rect 169436 79928 169492 79937
rect 169634 79937 169662 80036
rect 169530 79902 169582 79908
rect 169620 79928 169676 79937
rect 169436 79863 169492 79872
rect 169726 79898 169754 80036
rect 169818 79937 169846 80036
rect 169804 79928 169860 79937
rect 169620 79863 169676 79872
rect 169714 79892 169766 79898
rect 169804 79863 169860 79872
rect 169714 79834 169766 79840
rect 169910 79830 169938 80036
rect 170002 79830 170030 80036
rect 169898 79824 169950 79830
rect 169358 79801 169432 79812
rect 168748 79766 168800 79772
rect 169022 79792 169078 79801
rect 168562 79727 168618 79736
rect 168288 73636 168340 73642
rect 168288 73578 168340 73584
rect 168288 73160 168340 73166
rect 168288 73102 168340 73108
rect 168196 17400 168248 17406
rect 168196 17342 168248 17348
rect 168300 6254 168328 73102
rect 168392 55146 168420 79727
rect 168472 79620 168524 79626
rect 168472 79562 168524 79568
rect 168484 75954 168512 79562
rect 168472 75948 168524 75954
rect 168472 75890 168524 75896
rect 168472 74996 168524 75002
rect 168472 74938 168524 74944
rect 168484 57934 168512 74938
rect 168576 63442 168604 79727
rect 168668 78402 168696 79766
rect 168760 78985 168788 79766
rect 168840 79756 168892 79762
rect 169358 79792 169446 79801
rect 169358 79784 169390 79792
rect 169022 79727 169078 79736
rect 169116 79756 169168 79762
rect 168840 79698 168892 79704
rect 168746 78976 168802 78985
rect 168746 78911 168802 78920
rect 168852 78577 168880 79698
rect 168930 79520 168986 79529
rect 168930 79455 168932 79464
rect 168984 79455 168986 79464
rect 168932 79426 168984 79432
rect 168838 78568 168894 78577
rect 168838 78503 168894 78512
rect 168656 78396 168708 78402
rect 168656 78338 168708 78344
rect 168840 78396 168892 78402
rect 168840 78338 168892 78344
rect 168748 78328 168800 78334
rect 168748 78270 168800 78276
rect 168656 78056 168708 78062
rect 168656 77998 168708 78004
rect 168668 64734 168696 77998
rect 168760 75682 168788 78270
rect 168852 76906 168880 78338
rect 168930 78296 168986 78305
rect 168930 78231 168986 78240
rect 168840 76900 168892 76906
rect 168840 76842 168892 76848
rect 168840 75948 168892 75954
rect 168840 75890 168892 75896
rect 168748 75676 168800 75682
rect 168748 75618 168800 75624
rect 168748 75472 168800 75478
rect 168748 75414 168800 75420
rect 168760 67425 168788 75414
rect 168852 68746 168880 75890
rect 168944 75313 168972 78231
rect 169036 77294 169064 79727
rect 169116 79698 169168 79704
rect 169208 79756 169260 79762
rect 169758 79792 169814 79801
rect 169390 79727 169446 79736
rect 169484 79756 169536 79762
rect 169208 79698 169260 79704
rect 169898 79766 169950 79772
rect 169990 79824 170042 79830
rect 170094 79801 170122 80036
rect 170186 79830 170214 80036
rect 170278 79830 170306 80036
rect 170174 79824 170226 79830
rect 169990 79766 170042 79772
rect 170080 79792 170136 79801
rect 169758 79727 169814 79736
rect 170174 79766 170226 79772
rect 170266 79824 170318 79830
rect 170266 79766 170318 79772
rect 170080 79727 170136 79736
rect 169484 79698 169536 79704
rect 169128 77897 169156 79698
rect 169114 77888 169170 77897
rect 169114 77823 169170 77832
rect 169220 77294 169248 79698
rect 169392 79688 169444 79694
rect 169392 79630 169444 79636
rect 169300 79416 169352 79422
rect 169300 79358 169352 79364
rect 169312 78334 169340 79358
rect 169300 78328 169352 78334
rect 169300 78270 169352 78276
rect 169404 78062 169432 79630
rect 169392 78056 169444 78062
rect 169392 77998 169444 78004
rect 169036 77266 169156 77294
rect 169220 77266 169432 77294
rect 168930 75304 168986 75313
rect 168930 75239 168986 75248
rect 169024 75132 169076 75138
rect 169024 75074 169076 75080
rect 169036 74934 169064 75074
rect 169024 74928 169076 74934
rect 169024 74870 169076 74876
rect 169128 72457 169156 77266
rect 169208 76900 169260 76906
rect 169208 76842 169260 76848
rect 169220 73710 169248 76842
rect 169404 75002 169432 77266
rect 169496 75478 169524 79698
rect 169772 79608 169800 79727
rect 170036 79688 170088 79694
rect 170370 79676 170398 80036
rect 170462 79971 170490 80036
rect 170448 79962 170504 79971
rect 170448 79897 170504 79906
rect 170554 79812 170582 80036
rect 170646 79971 170674 80036
rect 170632 79962 170688 79971
rect 170632 79897 170688 79906
rect 170738 79898 170766 80036
rect 170830 79898 170858 80036
rect 170922 79966 170950 80036
rect 170910 79960 170962 79966
rect 171014 79937 171042 80036
rect 170910 79902 170962 79908
rect 171000 79928 171056 79937
rect 170726 79892 170778 79898
rect 170726 79834 170778 79840
rect 170818 79892 170870 79898
rect 171000 79863 171056 79872
rect 170818 79834 170870 79840
rect 171106 79812 171134 80036
rect 170554 79784 170628 79812
rect 170600 79744 170628 79784
rect 170954 79792 171010 79801
rect 170600 79716 170812 79744
rect 170954 79727 171010 79736
rect 171060 79784 171134 79812
rect 171198 79812 171226 80036
rect 171290 79966 171318 80036
rect 171382 79966 171410 80036
rect 171278 79960 171330 79966
rect 171278 79902 171330 79908
rect 171370 79960 171422 79966
rect 171474 79937 171502 80036
rect 171566 79966 171594 80036
rect 171658 79966 171686 80036
rect 171554 79960 171606 79966
rect 171370 79902 171422 79908
rect 171460 79928 171516 79937
rect 171554 79902 171606 79908
rect 171646 79960 171698 79966
rect 171646 79902 171698 79908
rect 171750 79898 171778 80036
rect 171842 79966 171870 80036
rect 171934 79966 171962 80036
rect 171830 79960 171882 79966
rect 171830 79902 171882 79908
rect 171922 79960 171974 79966
rect 171922 79902 171974 79908
rect 171460 79863 171516 79872
rect 171738 79892 171790 79898
rect 171738 79834 171790 79840
rect 171198 79801 171272 79812
rect 171198 79792 171286 79801
rect 171198 79784 171230 79792
rect 170036 79630 170088 79636
rect 170218 79656 170274 79665
rect 169680 79580 169800 79608
rect 169852 79620 169904 79626
rect 169576 79552 169628 79558
rect 169576 79494 169628 79500
rect 169588 78033 169616 79494
rect 169680 78402 169708 79580
rect 169852 79562 169904 79568
rect 169944 79620 169996 79626
rect 169944 79562 169996 79568
rect 169760 79484 169812 79490
rect 169760 79426 169812 79432
rect 169668 78396 169720 78402
rect 169668 78338 169720 78344
rect 169668 78260 169720 78266
rect 169668 78202 169720 78208
rect 169574 78024 169630 78033
rect 169574 77959 169630 77968
rect 169680 76838 169708 78202
rect 169668 76832 169720 76838
rect 169668 76774 169720 76780
rect 169576 75676 169628 75682
rect 169576 75618 169628 75624
rect 169484 75472 169536 75478
rect 169484 75414 169536 75420
rect 169482 75304 169538 75313
rect 169482 75239 169538 75248
rect 169392 74996 169444 75002
rect 169392 74938 169444 74944
rect 169208 73704 169260 73710
rect 169208 73646 169260 73652
rect 169114 72448 169170 72457
rect 169114 72383 169170 72392
rect 168840 68740 168892 68746
rect 168840 68682 168892 68688
rect 169392 68740 169444 68746
rect 169392 68682 169444 68688
rect 168746 67416 168802 67425
rect 168746 67351 168802 67360
rect 168656 64728 168708 64734
rect 168656 64670 168708 64676
rect 168564 63436 168616 63442
rect 168564 63378 168616 63384
rect 169300 63436 169352 63442
rect 169300 63378 169352 63384
rect 168472 57928 168524 57934
rect 168472 57870 168524 57876
rect 168380 55140 168432 55146
rect 168380 55082 168432 55088
rect 168472 37936 168524 37942
rect 168472 37878 168524 37884
rect 168484 16574 168512 37878
rect 169312 35290 169340 63378
rect 169404 38078 169432 68682
rect 169392 38072 169444 38078
rect 169392 38014 169444 38020
rect 169496 38010 169524 75239
rect 169588 71330 169616 75618
rect 169576 71324 169628 71330
rect 169576 71266 169628 71272
rect 169484 38004 169536 38010
rect 169484 37946 169536 37952
rect 169300 35284 169352 35290
rect 169300 35226 169352 35232
rect 169588 31074 169616 71266
rect 169666 67416 169722 67425
rect 169666 67351 169722 67360
rect 169576 31068 169628 31074
rect 169576 31010 169628 31016
rect 169680 17338 169708 67351
rect 169772 42090 169800 79426
rect 169864 75478 169892 79562
rect 169852 75472 169904 75478
rect 169852 75414 169904 75420
rect 169956 71738 169984 79562
rect 169944 71732 169996 71738
rect 169944 71674 169996 71680
rect 170048 71398 170076 79630
rect 170128 79620 170180 79626
rect 170370 79648 170444 79676
rect 170218 79591 170274 79600
rect 170128 79562 170180 79568
rect 170140 78441 170168 79562
rect 170126 78432 170182 78441
rect 170126 78367 170182 78376
rect 170232 76770 170260 79591
rect 170220 76764 170272 76770
rect 170220 76706 170272 76712
rect 170416 76673 170444 79648
rect 170680 79620 170732 79626
rect 170680 79562 170732 79568
rect 170496 79008 170548 79014
rect 170496 78950 170548 78956
rect 170402 76664 170458 76673
rect 170402 76599 170458 76608
rect 170126 76528 170182 76537
rect 170126 76463 170182 76472
rect 170140 76294 170168 76463
rect 170128 76288 170180 76294
rect 170128 76230 170180 76236
rect 170036 71392 170088 71398
rect 170036 71334 170088 71340
rect 170140 70394 170168 76230
rect 170416 73154 170444 76599
rect 170508 76537 170536 78950
rect 170586 78568 170642 78577
rect 170586 78503 170642 78512
rect 170494 76528 170550 76537
rect 170494 76463 170550 76472
rect 170600 76362 170628 78503
rect 170588 76356 170640 76362
rect 170588 76298 170640 76304
rect 170416 73126 170628 73154
rect 170600 70394 170628 73126
rect 170692 71777 170720 79562
rect 170784 79014 170812 79716
rect 170864 79688 170916 79694
rect 170864 79630 170916 79636
rect 170772 79008 170824 79014
rect 170772 78950 170824 78956
rect 170772 76356 170824 76362
rect 170772 76298 170824 76304
rect 170784 76158 170812 76298
rect 170772 76152 170824 76158
rect 170772 76094 170824 76100
rect 170678 71768 170734 71777
rect 170678 71703 170734 71712
rect 170140 70366 170536 70394
rect 170600 70366 170720 70394
rect 169760 42084 169812 42090
rect 169760 42026 169812 42032
rect 170508 36718 170536 70366
rect 170496 36712 170548 36718
rect 170496 36654 170548 36660
rect 170692 33930 170720 70366
rect 170680 33924 170732 33930
rect 170680 33866 170732 33872
rect 170784 29714 170812 76094
rect 170876 75546 170904 79630
rect 170968 75818 170996 79727
rect 171060 76129 171088 79784
rect 172026 79778 172054 80036
rect 172118 79966 172146 80036
rect 172106 79960 172158 79966
rect 172106 79902 172158 79908
rect 172210 79898 172238 80036
rect 172302 79966 172330 80036
rect 172290 79960 172342 79966
rect 172290 79902 172342 79908
rect 172198 79892 172250 79898
rect 172198 79834 172250 79840
rect 172394 79830 172422 80036
rect 172382 79824 172434 79830
rect 172150 79792 172206 79801
rect 171230 79727 171286 79736
rect 171416 79756 171468 79762
rect 171416 79698 171468 79704
rect 171508 79756 171560 79762
rect 171508 79698 171560 79704
rect 171796 79750 172150 79778
rect 171322 79656 171378 79665
rect 171232 79620 171284 79626
rect 171322 79591 171378 79600
rect 171232 79562 171284 79568
rect 171140 79416 171192 79422
rect 171140 79358 171192 79364
rect 171046 76120 171102 76129
rect 171046 76055 171102 76064
rect 170956 75812 171008 75818
rect 170956 75754 171008 75760
rect 170864 75540 170916 75546
rect 170864 75482 170916 75488
rect 170876 73154 170904 75482
rect 171048 75472 171100 75478
rect 171048 75414 171100 75420
rect 171060 74186 171088 75414
rect 171048 74180 171100 74186
rect 171048 74122 171100 74128
rect 170876 73126 170996 73154
rect 170864 71392 170916 71398
rect 170864 71334 170916 71340
rect 170876 70990 170904 71334
rect 170864 70984 170916 70990
rect 170864 70926 170916 70932
rect 170772 29708 170824 29714
rect 170772 29650 170824 29656
rect 169668 17332 169720 17338
rect 169668 17274 169720 17280
rect 168484 16546 169616 16574
rect 168288 6248 168340 6254
rect 168288 6190 168340 6196
rect 167644 3460 167696 3466
rect 167644 3402 167696 3408
rect 168380 3460 168432 3466
rect 168380 3402 168432 3408
rect 168392 480 168420 3402
rect 169588 480 169616 16546
rect 170876 13122 170904 70926
rect 170968 14482 170996 73126
rect 170956 14476 171008 14482
rect 170956 14418 171008 14424
rect 170864 13116 170916 13122
rect 170864 13058 170916 13064
rect 171060 4894 171088 74122
rect 171152 25634 171180 79358
rect 171244 26994 171272 79562
rect 171336 28354 171364 79591
rect 171428 78577 171456 79698
rect 171414 78568 171470 78577
rect 171414 78503 171470 78512
rect 171416 75472 171468 75478
rect 171416 75414 171468 75420
rect 171428 68814 171456 75414
rect 171520 68882 171548 79698
rect 171600 79688 171652 79694
rect 171600 79630 171652 79636
rect 171612 76537 171640 79630
rect 171796 79422 171824 79750
rect 172382 79766 172434 79772
rect 172150 79727 172206 79736
rect 172244 79756 172296 79762
rect 172244 79698 172296 79704
rect 171968 79688 172020 79694
rect 171968 79630 172020 79636
rect 171876 79620 171928 79626
rect 171876 79562 171928 79568
rect 171784 79416 171836 79422
rect 171784 79358 171836 79364
rect 171888 79098 171916 79562
rect 171796 79070 171916 79098
rect 171796 77058 171824 79070
rect 171876 78668 171928 78674
rect 171876 78610 171928 78616
rect 171888 78169 171916 78610
rect 171874 78160 171930 78169
rect 171874 78095 171930 78104
rect 171980 77761 172008 79630
rect 172060 79620 172112 79626
rect 172060 79562 172112 79568
rect 172152 79620 172204 79626
rect 172152 79562 172204 79568
rect 171966 77752 172022 77761
rect 171966 77687 172022 77696
rect 171796 77030 171916 77058
rect 171784 76968 171836 76974
rect 171784 76910 171836 76916
rect 171598 76528 171654 76537
rect 171598 76463 171654 76472
rect 171796 76430 171824 76910
rect 171784 76424 171836 76430
rect 171784 76366 171836 76372
rect 171888 75682 171916 77030
rect 171968 76764 172020 76770
rect 171968 76706 172020 76712
rect 171876 75676 171928 75682
rect 171876 75618 171928 75624
rect 171784 71392 171836 71398
rect 171784 71334 171836 71340
rect 171796 70854 171824 71334
rect 171784 70848 171836 70854
rect 171784 70790 171836 70796
rect 171980 70394 172008 76706
rect 172072 75478 172100 79562
rect 172164 76537 172192 79562
rect 172150 76528 172206 76537
rect 172150 76463 172206 76472
rect 172256 75954 172284 79698
rect 172486 79676 172514 80036
rect 172578 79830 172606 80036
rect 172670 79966 172698 80036
rect 172658 79960 172710 79966
rect 172658 79902 172710 79908
rect 172762 79898 172790 80036
rect 172854 79937 172882 80036
rect 172840 79928 172896 79937
rect 172750 79892 172802 79898
rect 172840 79863 172896 79872
rect 172750 79834 172802 79840
rect 172566 79824 172618 79830
rect 172566 79766 172618 79772
rect 172702 79792 172758 79801
rect 172702 79727 172758 79736
rect 172946 79744 172974 80036
rect 173038 79898 173066 80036
rect 173026 79892 173078 79898
rect 173026 79834 173078 79840
rect 173130 79801 173158 80036
rect 173116 79792 173172 79801
rect 172348 79648 172514 79676
rect 172612 79688 172664 79694
rect 172348 76537 172376 79648
rect 172612 79630 172664 79636
rect 172428 79552 172480 79558
rect 172428 79494 172480 79500
rect 172334 76528 172390 76537
rect 172334 76463 172390 76472
rect 172440 76106 172468 79494
rect 172520 79144 172572 79150
rect 172520 79086 172572 79092
rect 172532 78266 172560 79086
rect 172520 78260 172572 78266
rect 172520 78202 172572 78208
rect 172520 77852 172572 77858
rect 172520 77794 172572 77800
rect 172348 76078 172468 76106
rect 172244 75948 172296 75954
rect 172244 75890 172296 75896
rect 172242 75848 172298 75857
rect 172242 75783 172298 75792
rect 172060 75472 172112 75478
rect 172060 75414 172112 75420
rect 172256 75313 172284 75783
rect 172348 75750 172376 76078
rect 172428 75948 172480 75954
rect 172428 75890 172480 75896
rect 172336 75744 172388 75750
rect 172336 75686 172388 75692
rect 172242 75304 172298 75313
rect 172242 75239 172298 75248
rect 171980 70366 172100 70394
rect 171508 68876 171560 68882
rect 171508 68818 171560 68824
rect 171416 68808 171468 68814
rect 171416 68750 171468 68756
rect 172072 53786 172100 70366
rect 172152 68876 172204 68882
rect 172152 68818 172204 68824
rect 172164 68202 172192 68818
rect 172152 68196 172204 68202
rect 172152 68138 172204 68144
rect 172060 53780 172112 53786
rect 172060 53722 172112 53728
rect 172164 36650 172192 68138
rect 172256 40798 172284 75239
rect 172440 74254 172468 75890
rect 172428 74248 172480 74254
rect 172428 74190 172480 74196
rect 172336 68808 172388 68814
rect 172336 68750 172388 68756
rect 172348 68542 172376 68750
rect 172336 68536 172388 68542
rect 172336 68478 172388 68484
rect 172244 40792 172296 40798
rect 172244 40734 172296 40740
rect 172152 36644 172204 36650
rect 172152 36586 172204 36592
rect 171784 33788 171836 33794
rect 171784 33730 171836 33736
rect 171324 28348 171376 28354
rect 171324 28290 171376 28296
rect 171232 26988 171284 26994
rect 171232 26930 171284 26936
rect 171140 25628 171192 25634
rect 171140 25570 171192 25576
rect 171048 4888 171100 4894
rect 171048 4830 171100 4836
rect 170772 3800 170824 3806
rect 170772 3742 170824 3748
rect 170784 480 170812 3742
rect 171796 3466 171824 33730
rect 172348 26926 172376 68478
rect 171876 26920 171928 26926
rect 171876 26862 171928 26868
rect 172336 26920 172388 26926
rect 172336 26862 172388 26868
rect 171784 3460 171836 3466
rect 171784 3402 171836 3408
rect 171888 2990 171916 26862
rect 172440 24206 172468 74190
rect 172532 37942 172560 77794
rect 172624 76770 172652 79630
rect 172716 78674 172744 79727
rect 172946 79716 173020 79744
rect 173116 79727 173172 79736
rect 172794 79656 172850 79665
rect 172794 79591 172850 79600
rect 172704 78668 172756 78674
rect 172704 78610 172756 78616
rect 172702 78432 172758 78441
rect 172702 78367 172758 78376
rect 172612 76764 172664 76770
rect 172612 76706 172664 76712
rect 172716 76650 172744 78367
rect 172808 77858 172836 79591
rect 172992 79422 173020 79716
rect 173222 79540 173250 80036
rect 173314 79830 173342 80036
rect 173302 79824 173354 79830
rect 173406 79801 173434 80036
rect 173302 79766 173354 79772
rect 173392 79792 173448 79801
rect 173392 79727 173448 79736
rect 173348 79688 173400 79694
rect 173498 79676 173526 80036
rect 173590 79744 173618 80036
rect 173682 79937 173710 80036
rect 173668 79928 173724 79937
rect 173668 79863 173724 79872
rect 173590 79716 173664 79744
rect 173348 79630 173400 79636
rect 173452 79648 173526 79676
rect 173636 79676 173664 79716
rect 173774 79676 173802 80036
rect 173866 79801 173894 80036
rect 173958 79830 173986 80036
rect 174050 79966 174078 80036
rect 174142 79971 174170 80036
rect 174038 79960 174090 79966
rect 174038 79902 174090 79908
rect 174128 79962 174184 79971
rect 174128 79897 174184 79906
rect 174234 79898 174262 80036
rect 174222 79892 174274 79898
rect 173946 79824 173998 79830
rect 173852 79792 173908 79801
rect 173946 79766 173998 79772
rect 174128 79826 174184 79835
rect 174222 79834 174274 79840
rect 174326 79812 174354 80036
rect 174418 79937 174446 80036
rect 174510 79966 174538 80036
rect 174602 79966 174630 80036
rect 174694 79966 174722 80036
rect 174498 79960 174550 79966
rect 174404 79928 174460 79937
rect 174498 79902 174550 79908
rect 174590 79960 174642 79966
rect 174590 79902 174642 79908
rect 174682 79960 174734 79966
rect 174786 79937 174814 80036
rect 174682 79902 174734 79908
rect 174772 79928 174828 79937
rect 174404 79863 174460 79872
rect 174772 79863 174828 79872
rect 174544 79824 174596 79830
rect 174326 79784 174446 79812
rect 174184 79770 174216 79778
rect 174128 79761 174216 79770
rect 174142 79750 174216 79761
rect 173852 79727 173908 79736
rect 173900 79688 173952 79694
rect 173636 79648 173710 79676
rect 173774 79648 173848 79676
rect 173176 79512 173250 79540
rect 172888 79416 172940 79422
rect 172888 79358 172940 79364
rect 172980 79416 173032 79422
rect 172980 79358 173032 79364
rect 172900 78985 172928 79358
rect 173072 79348 173124 79354
rect 173072 79290 173124 79296
rect 172980 79280 173032 79286
rect 172980 79222 173032 79228
rect 172886 78976 172942 78985
rect 172886 78911 172942 78920
rect 172992 78674 173020 79222
rect 173084 79218 173112 79290
rect 173072 79212 173124 79218
rect 173072 79154 173124 79160
rect 172888 78668 172940 78674
rect 172888 78610 172940 78616
rect 172980 78668 173032 78674
rect 172980 78610 173032 78616
rect 172796 77852 172848 77858
rect 172796 77794 172848 77800
rect 172624 76622 172744 76650
rect 172624 45558 172652 76622
rect 172704 76220 172756 76226
rect 172704 76162 172756 76168
rect 172716 62082 172744 76162
rect 172796 75472 172848 75478
rect 172796 75414 172848 75420
rect 172808 66230 172836 75414
rect 172900 75070 172928 78610
rect 172888 75064 172940 75070
rect 172888 75006 172940 75012
rect 173176 70394 173204 79512
rect 173256 79416 173308 79422
rect 173256 79358 173308 79364
rect 173268 75721 173296 79358
rect 173360 79014 173388 79630
rect 173348 79008 173400 79014
rect 173348 78950 173400 78956
rect 173452 77761 173480 79648
rect 173532 79552 173584 79558
rect 173682 79540 173710 79648
rect 173532 79494 173584 79500
rect 173636 79512 173710 79540
rect 173438 77752 173494 77761
rect 173438 77687 173494 77696
rect 173544 76906 173572 79494
rect 173532 76900 173584 76906
rect 173532 76842 173584 76848
rect 173532 76764 173584 76770
rect 173532 76706 173584 76712
rect 173440 76424 173492 76430
rect 173440 76366 173492 76372
rect 173254 75712 173310 75721
rect 173254 75647 173310 75656
rect 173452 71641 173480 76366
rect 173438 71632 173494 71641
rect 173438 71567 173494 71576
rect 172900 70366 173204 70394
rect 172900 68882 172928 70366
rect 172888 68876 172940 68882
rect 172888 68818 172940 68824
rect 172796 66224 172848 66230
rect 172796 66166 172848 66172
rect 172704 62076 172756 62082
rect 172704 62018 172756 62024
rect 172612 45552 172664 45558
rect 172612 45494 172664 45500
rect 173544 39438 173572 76706
rect 173636 76226 173664 79512
rect 173714 78432 173770 78441
rect 173714 78367 173770 78376
rect 173728 76430 173756 78367
rect 173716 76424 173768 76430
rect 173716 76366 173768 76372
rect 173624 76220 173676 76226
rect 173624 76162 173676 76168
rect 173820 75478 173848 79648
rect 173900 79630 173952 79636
rect 173912 78334 173940 79630
rect 173992 79484 174044 79490
rect 173992 79426 174044 79432
rect 174004 79218 174032 79426
rect 173992 79212 174044 79218
rect 173992 79154 174044 79160
rect 174084 79212 174136 79218
rect 174084 79154 174136 79160
rect 173990 78432 174046 78441
rect 173990 78367 174046 78376
rect 173900 78328 173952 78334
rect 173900 78270 173952 78276
rect 173900 77988 173952 77994
rect 173900 77930 173952 77936
rect 173808 75472 173860 75478
rect 173808 75414 173860 75420
rect 173808 75064 173860 75070
rect 173808 75006 173860 75012
rect 173820 74118 173848 75006
rect 173808 74112 173860 74118
rect 173808 74054 173860 74060
rect 173716 68876 173768 68882
rect 173716 68818 173768 68824
rect 173728 68270 173756 68818
rect 173716 68264 173768 68270
rect 173716 68206 173768 68212
rect 173624 66224 173676 66230
rect 173624 66166 173676 66172
rect 173636 66026 173664 66166
rect 173624 66020 173676 66026
rect 173624 65962 173676 65968
rect 173532 39432 173584 39438
rect 173532 39374 173584 39380
rect 172520 37936 172572 37942
rect 172520 37878 172572 37884
rect 172428 24200 172480 24206
rect 172428 24142 172480 24148
rect 173636 24138 173664 65962
rect 173728 25566 173756 68206
rect 173716 25560 173768 25566
rect 173716 25502 173768 25508
rect 173624 24132 173676 24138
rect 173624 24074 173676 24080
rect 173820 22846 173848 74054
rect 173808 22840 173860 22846
rect 173808 22782 173860 22788
rect 173162 22672 173218 22681
rect 173162 22607 173218 22616
rect 173176 16574 173204 22607
rect 173176 16546 173296 16574
rect 173268 3534 173296 16546
rect 173912 7614 173940 77930
rect 174004 10334 174032 78367
rect 174096 11762 174124 79154
rect 174188 76430 174216 79750
rect 174268 79688 174320 79694
rect 174418 79642 174446 79784
rect 174544 79766 174596 79772
rect 174268 79630 174320 79636
rect 174280 78985 174308 79630
rect 174372 79614 174446 79642
rect 174266 78976 174322 78985
rect 174266 78911 174322 78920
rect 174280 77994 174308 78911
rect 174268 77988 174320 77994
rect 174268 77930 174320 77936
rect 174268 76900 174320 76906
rect 174268 76842 174320 76848
rect 174176 76424 174228 76430
rect 174176 76366 174228 76372
rect 174176 76220 174228 76226
rect 174176 76162 174228 76168
rect 174188 64870 174216 76162
rect 174280 72865 174308 76842
rect 174266 72856 174322 72865
rect 174266 72791 174322 72800
rect 174372 70394 174400 79614
rect 174452 79348 174504 79354
rect 174452 79290 174504 79296
rect 174464 79150 174492 79290
rect 174556 79218 174584 79766
rect 174878 79744 174906 80036
rect 174832 79716 174906 79744
rect 174970 79744 174998 80036
rect 175062 79937 175090 80036
rect 175048 79928 175104 79937
rect 175048 79863 175104 79872
rect 175154 79778 175182 80036
rect 175246 79801 175274 80036
rect 175338 79966 175366 80036
rect 175326 79960 175378 79966
rect 175326 79902 175378 79908
rect 175430 79812 175458 80036
rect 175522 79830 175550 80036
rect 175614 79971 175642 80036
rect 175600 79962 175656 79971
rect 175600 79897 175656 79906
rect 175706 79898 175734 80036
rect 175798 79903 175826 80036
rect 175890 79966 175918 80036
rect 175982 79966 176010 80036
rect 176074 79971 176102 80036
rect 175878 79960 175930 79966
rect 175694 79892 175746 79898
rect 175694 79834 175746 79840
rect 175784 79894 175840 79903
rect 175878 79902 175930 79908
rect 175970 79960 176022 79966
rect 175970 79902 176022 79908
rect 176060 79962 176116 79971
rect 176166 79966 176194 80036
rect 176060 79897 176116 79906
rect 176154 79960 176206 79966
rect 176258 79937 176286 80036
rect 176350 79966 176378 80036
rect 176442 79966 176470 80036
rect 176338 79960 176390 79966
rect 176154 79902 176206 79908
rect 176244 79928 176300 79937
rect 176338 79902 176390 79908
rect 176430 79960 176482 79966
rect 176430 79902 176482 79908
rect 176244 79863 176300 79872
rect 175108 79750 175182 79778
rect 175232 79792 175288 79801
rect 174970 79716 175044 79744
rect 174728 79688 174780 79694
rect 174634 79656 174690 79665
rect 174728 79630 174780 79636
rect 174634 79591 174690 79600
rect 174544 79212 174596 79218
rect 174544 79154 174596 79160
rect 174648 79150 174676 79591
rect 174452 79144 174504 79150
rect 174452 79086 174504 79092
rect 174636 79144 174688 79150
rect 174636 79086 174688 79092
rect 174636 78328 174688 78334
rect 174636 78270 174688 78276
rect 174648 75478 174676 78270
rect 174740 76537 174768 79630
rect 174832 76945 174860 79716
rect 174912 79416 174964 79422
rect 174912 79358 174964 79364
rect 174924 78674 174952 79358
rect 174912 78668 174964 78674
rect 174912 78610 174964 78616
rect 174818 76936 174874 76945
rect 174818 76871 174874 76880
rect 174726 76528 174782 76537
rect 174726 76463 174782 76472
rect 174636 75472 174688 75478
rect 174636 75414 174688 75420
rect 174450 72856 174506 72865
rect 174450 72791 174506 72800
rect 174280 70366 174400 70394
rect 174280 69630 174308 70366
rect 174268 69624 174320 69630
rect 174268 69566 174320 69572
rect 174464 64874 174492 72791
rect 174648 67634 174676 75414
rect 175016 71369 175044 79716
rect 175108 76537 175136 79750
rect 175232 79727 175288 79736
rect 175384 79784 175458 79812
rect 175510 79824 175562 79830
rect 175784 79829 175840 79838
rect 175188 79688 175240 79694
rect 175188 79630 175240 79636
rect 175280 79688 175332 79694
rect 175280 79630 175332 79636
rect 175094 76528 175150 76537
rect 175094 76463 175150 76472
rect 175200 76226 175228 79630
rect 175188 76220 175240 76226
rect 175188 76162 175240 76168
rect 175186 75576 175242 75585
rect 175186 75511 175242 75520
rect 175200 73778 175228 75511
rect 175188 73772 175240 73778
rect 175188 73714 175240 73720
rect 175002 71360 175058 71369
rect 175002 71295 175058 71304
rect 175096 69624 175148 69630
rect 175096 69566 175148 69572
rect 174648 67606 175044 67634
rect 174176 64864 174228 64870
rect 174464 64846 174952 64874
rect 174176 64806 174228 64812
rect 174924 40730 174952 64846
rect 174912 40724 174964 40730
rect 174912 40666 174964 40672
rect 175016 36582 175044 67606
rect 175004 36576 175056 36582
rect 175004 36518 175056 36524
rect 175108 22778 175136 69566
rect 175096 22772 175148 22778
rect 175096 22714 175148 22720
rect 174084 11756 174136 11762
rect 174084 11698 174136 11704
rect 173992 10328 174044 10334
rect 173992 10270 174044 10276
rect 173900 7608 173952 7614
rect 173900 7550 173952 7556
rect 175200 4826 175228 73714
rect 175292 35222 175320 79630
rect 175384 78334 175412 79784
rect 175510 79766 175562 79772
rect 175832 79756 175884 79762
rect 175832 79698 175884 79704
rect 176016 79756 176068 79762
rect 176016 79698 176068 79704
rect 176200 79756 176252 79762
rect 176200 79698 176252 79704
rect 176384 79756 176436 79762
rect 176534 79744 176562 80036
rect 176626 79898 176654 80036
rect 176614 79892 176666 79898
rect 176614 79834 176666 79840
rect 176718 79744 176746 80036
rect 176810 79898 176838 80036
rect 176902 79966 176930 80036
rect 176890 79960 176942 79966
rect 176890 79902 176942 79908
rect 176798 79892 176850 79898
rect 176798 79834 176850 79840
rect 176994 79744 177022 80036
rect 177086 79966 177114 80036
rect 177074 79960 177126 79966
rect 177074 79902 177126 79908
rect 177178 79898 177206 80036
rect 177166 79892 177218 79898
rect 177166 79834 177218 79840
rect 177270 79778 177298 80036
rect 177362 79812 177390 80036
rect 177454 79937 177482 80036
rect 177546 79948 177574 80036
rect 177652 80022 177988 80050
rect 177764 79960 177816 79966
rect 177440 79928 177496 79937
rect 177546 79920 177620 79948
rect 177440 79863 177496 79872
rect 177362 79784 177436 79812
rect 176534 79716 176608 79744
rect 176384 79698 176436 79704
rect 175464 79688 175516 79694
rect 175464 79630 175516 79636
rect 175554 79656 175610 79665
rect 175372 78328 175424 78334
rect 175372 78270 175424 78276
rect 175372 76900 175424 76906
rect 175372 76842 175424 76848
rect 175384 66230 175412 76842
rect 175476 67182 175504 79630
rect 175554 79591 175610 79600
rect 175738 79656 175794 79665
rect 175738 79591 175794 79600
rect 175568 74934 175596 79591
rect 175556 74928 175608 74934
rect 175556 74870 175608 74876
rect 175752 70394 175780 79591
rect 175844 76158 175872 79698
rect 175924 79620 175976 79626
rect 175924 79562 175976 79568
rect 175936 77858 175964 79562
rect 175924 77852 175976 77858
rect 175924 77794 175976 77800
rect 176028 76650 176056 79698
rect 176108 79620 176160 79626
rect 176108 79562 176160 79568
rect 176120 76945 176148 79562
rect 176106 76936 176162 76945
rect 176106 76871 176162 76880
rect 175936 76622 176056 76650
rect 175832 76152 175884 76158
rect 175832 76094 175884 76100
rect 175936 72865 175964 76622
rect 176212 76537 176240 79698
rect 176292 79688 176344 79694
rect 176292 79630 176344 79636
rect 176198 76528 176254 76537
rect 176198 76463 176254 76472
rect 176304 76265 176332 79630
rect 176396 76650 176424 79698
rect 176580 76906 176608 79716
rect 176672 79716 176746 79744
rect 176856 79716 177022 79744
rect 177120 79756 177172 79762
rect 176672 79558 176700 79716
rect 176856 79642 176884 79716
rect 177120 79698 177172 79704
rect 177224 79750 177298 79778
rect 176764 79614 176884 79642
rect 176936 79620 176988 79626
rect 176660 79552 176712 79558
rect 176660 79494 176712 79500
rect 176660 78668 176712 78674
rect 176660 78610 176712 78616
rect 176568 76900 176620 76906
rect 176568 76842 176620 76848
rect 176396 76622 176516 76650
rect 176384 76356 176436 76362
rect 176384 76298 176436 76304
rect 176290 76256 176346 76265
rect 176290 76191 176346 76200
rect 176108 76152 176160 76158
rect 176108 76094 176160 76100
rect 176120 75585 176148 76094
rect 176106 75576 176162 75585
rect 176106 75511 176162 75520
rect 175922 72856 175978 72865
rect 175922 72791 175978 72800
rect 175568 70366 175780 70394
rect 175568 70145 175596 70366
rect 175554 70136 175610 70145
rect 175554 70071 175610 70080
rect 175924 68808 175976 68814
rect 175924 68750 175976 68756
rect 175936 68134 175964 68750
rect 175924 68128 175976 68134
rect 175924 68070 175976 68076
rect 175464 67176 175516 67182
rect 175464 67118 175516 67124
rect 175372 66224 175424 66230
rect 175372 66166 175424 66172
rect 176120 39370 176148 75511
rect 176292 75268 176344 75274
rect 176292 75210 176344 75216
rect 176200 75200 176252 75206
rect 176200 75142 176252 75148
rect 176212 74905 176240 75142
rect 176304 75070 176332 75210
rect 176396 75138 176424 76298
rect 176384 75132 176436 75138
rect 176384 75074 176436 75080
rect 176292 75064 176344 75070
rect 176292 75006 176344 75012
rect 176292 74928 176344 74934
rect 176198 74896 176254 74905
rect 176292 74870 176344 74876
rect 176198 74831 176254 74840
rect 176304 74089 176332 74870
rect 176290 74080 176346 74089
rect 176290 74015 176346 74024
rect 176198 72584 176254 72593
rect 176198 72519 176254 72528
rect 176108 39364 176160 39370
rect 176108 39306 176160 39312
rect 175280 35216 175332 35222
rect 175280 35158 175332 35164
rect 176212 33862 176240 72519
rect 176304 72078 176332 74015
rect 176382 72856 176438 72865
rect 176382 72791 176438 72800
rect 176292 72072 176344 72078
rect 176292 72014 176344 72020
rect 176292 66224 176344 66230
rect 176292 66166 176344 66172
rect 176200 33856 176252 33862
rect 176200 33798 176252 33804
rect 176304 18698 176332 66166
rect 176292 18692 176344 18698
rect 176292 18634 176344 18640
rect 176396 15910 176424 72791
rect 176488 72593 176516 76622
rect 176566 76528 176622 76537
rect 176566 76463 176622 76472
rect 176474 72584 176530 72593
rect 176474 72519 176530 72528
rect 176476 72072 176528 72078
rect 176476 72014 176528 72020
rect 176384 15904 176436 15910
rect 176384 15846 176436 15852
rect 176488 8974 176516 72014
rect 176476 8968 176528 8974
rect 176476 8910 176528 8916
rect 176580 6186 176608 76463
rect 176672 44130 176700 78610
rect 176764 46918 176792 79614
rect 176936 79562 176988 79568
rect 177028 79620 177080 79626
rect 177028 79562 177080 79568
rect 176844 79552 176896 79558
rect 176844 79494 176896 79500
rect 176856 50998 176884 79494
rect 176948 75954 176976 79562
rect 176936 75948 176988 75954
rect 176936 75890 176988 75896
rect 176936 72616 176988 72622
rect 176936 72558 176988 72564
rect 176948 66230 176976 72558
rect 177040 67318 177068 79562
rect 177132 68921 177160 79698
rect 177224 78674 177252 79750
rect 177212 78668 177264 78674
rect 177212 78610 177264 78616
rect 177212 77852 177264 77858
rect 177212 77794 177264 77800
rect 177224 70394 177252 77794
rect 177304 75200 177356 75206
rect 177304 75142 177356 75148
rect 177316 74905 177344 75142
rect 177302 74896 177358 74905
rect 177302 74831 177358 74840
rect 177408 72622 177436 79784
rect 177592 78305 177620 79920
rect 177764 79902 177816 79908
rect 177578 78296 177634 78305
rect 177578 78231 177634 78240
rect 177672 76424 177724 76430
rect 177672 76366 177724 76372
rect 177396 72616 177448 72622
rect 177396 72558 177448 72564
rect 177224 70366 177528 70394
rect 177118 68912 177174 68921
rect 177118 68847 177174 68856
rect 177028 67312 177080 67318
rect 177028 67254 177080 67260
rect 176936 66224 176988 66230
rect 176936 66166 176988 66172
rect 176844 50992 176896 50998
rect 176844 50934 176896 50940
rect 176752 46912 176804 46918
rect 176752 46854 176804 46860
rect 176660 44124 176712 44130
rect 176660 44066 176712 44072
rect 177500 40050 177528 70366
rect 177684 68882 177712 76366
rect 177776 71505 177804 79902
rect 177960 77489 177988 80022
rect 177946 77480 178002 77489
rect 177946 77415 178002 77424
rect 177948 76900 178000 76906
rect 177948 76842 178000 76848
rect 177856 76424 177908 76430
rect 177856 76366 177908 76372
rect 177868 76294 177896 76366
rect 177856 76288 177908 76294
rect 177856 76230 177908 76236
rect 177960 75954 177988 76842
rect 177948 75948 178000 75954
rect 177948 75890 178000 75896
rect 177762 71496 177818 71505
rect 177762 71431 177818 71440
rect 177672 68876 177724 68882
rect 177672 68818 177724 68824
rect 177672 66224 177724 66230
rect 177672 66166 177724 66172
rect 177488 40044 177540 40050
rect 177488 39986 177540 39992
rect 177684 33794 177712 66166
rect 177672 33788 177724 33794
rect 177672 33730 177724 33736
rect 177776 29646 177804 71431
rect 177856 67312 177908 67318
rect 177856 67254 177908 67260
rect 177764 29640 177816 29646
rect 177764 29582 177816 29588
rect 177868 17270 177896 67254
rect 177960 18630 177988 75890
rect 178052 75041 178080 80106
rect 178144 75410 178172 80174
rect 178224 80096 178276 80102
rect 178224 80038 178276 80044
rect 178236 78985 178264 80038
rect 178222 78976 178278 78985
rect 178222 78911 178278 78920
rect 178224 78328 178276 78334
rect 178224 78270 178276 78276
rect 178236 76945 178264 78270
rect 178328 78169 178356 80310
rect 178420 80306 178448 80407
rect 181640 80345 181668 80543
rect 188344 80504 188396 80510
rect 188344 80446 188396 80452
rect 187056 80368 187108 80374
rect 181626 80336 181682 80345
rect 178408 80300 178460 80306
rect 187056 80310 187108 80316
rect 181626 80271 181682 80280
rect 178408 80242 178460 80248
rect 186964 80096 187016 80102
rect 186964 80038 187016 80044
rect 178776 80028 178828 80034
rect 178776 79970 178828 79976
rect 178314 78160 178370 78169
rect 178314 78095 178370 78104
rect 178222 76936 178278 76945
rect 178222 76871 178278 76880
rect 178684 76492 178736 76498
rect 178684 76434 178736 76440
rect 178132 75404 178184 75410
rect 178132 75346 178184 75352
rect 178038 75032 178094 75041
rect 178038 74967 178094 74976
rect 178038 71088 178094 71097
rect 178038 71023 178094 71032
rect 177948 18624 178000 18630
rect 177948 18566 178000 18572
rect 177856 17264 177908 17270
rect 177856 17206 177908 17212
rect 178052 16574 178080 71023
rect 178052 16546 178632 16574
rect 176568 6180 176620 6186
rect 176568 6122 176620 6128
rect 175188 4820 175240 4826
rect 175188 4762 175240 4768
rect 176660 3596 176712 3602
rect 176660 3538 176712 3544
rect 171968 3528 172020 3534
rect 171968 3470 172020 3476
rect 173256 3528 173308 3534
rect 173256 3470 173308 3476
rect 171876 2984 171928 2990
rect 171876 2926 171928 2932
rect 171980 480 172008 3470
rect 173164 3460 173216 3466
rect 173164 3402 173216 3408
rect 173176 480 173204 3402
rect 175464 3392 175516 3398
rect 175464 3334 175516 3340
rect 174268 2984 174320 2990
rect 174268 2926 174320 2932
rect 174280 480 174308 2926
rect 175476 480 175504 3334
rect 176672 480 176700 3538
rect 177856 3528 177908 3534
rect 177856 3470 177908 3476
rect 177868 480 177896 3470
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 178696 3534 178724 76434
rect 178788 56574 178816 79970
rect 180522 79928 180578 79937
rect 180522 79863 180578 79872
rect 180432 79688 180484 79694
rect 180432 79630 180484 79636
rect 178960 79620 179012 79626
rect 178960 79562 179012 79568
rect 178868 78056 178920 78062
rect 178868 77998 178920 78004
rect 178880 70854 178908 77998
rect 178972 77722 179000 79562
rect 179420 79484 179472 79490
rect 179420 79426 179472 79432
rect 179328 78736 179380 78742
rect 179328 78678 179380 78684
rect 179340 78334 179368 78678
rect 179328 78328 179380 78334
rect 179156 78276 179328 78282
rect 179156 78270 179380 78276
rect 179156 78254 179368 78270
rect 178960 77716 179012 77722
rect 178960 77658 179012 77664
rect 179052 73704 179104 73710
rect 179052 73646 179104 73652
rect 178868 70848 178920 70854
rect 178868 70790 178920 70796
rect 178880 70394 178908 70790
rect 178880 70366 179000 70394
rect 178776 56568 178828 56574
rect 178776 56510 178828 56516
rect 178972 3874 179000 70366
rect 178960 3868 179012 3874
rect 178960 3810 179012 3816
rect 178684 3528 178736 3534
rect 178684 3470 178736 3476
rect 179064 3466 179092 73646
rect 179156 6322 179184 78254
rect 179236 78124 179288 78130
rect 179236 78066 179288 78072
rect 179144 6316 179196 6322
rect 179144 6258 179196 6264
rect 179248 3942 179276 78066
rect 179328 77920 179380 77926
rect 179328 77862 179380 77868
rect 179340 77586 179368 77862
rect 179328 77580 179380 77586
rect 179328 77522 179380 77528
rect 179340 4010 179368 77522
rect 179328 4004 179380 4010
rect 179328 3946 179380 3952
rect 179236 3936 179288 3942
rect 179236 3878 179288 3884
rect 179432 3482 179460 79426
rect 179512 79348 179564 79354
rect 179512 79290 179564 79296
rect 179524 3602 179552 79290
rect 180444 78198 180472 79630
rect 180536 78441 180564 79863
rect 183744 79756 183796 79762
rect 183744 79698 183796 79704
rect 181442 78568 181498 78577
rect 181442 78503 181498 78512
rect 181626 78568 181682 78577
rect 181626 78503 181682 78512
rect 180522 78432 180578 78441
rect 180522 78367 180578 78376
rect 180156 78192 180208 78198
rect 180156 78134 180208 78140
rect 180432 78192 180484 78198
rect 180432 78134 180484 78140
rect 180616 78192 180668 78198
rect 181456 78169 181484 78503
rect 180616 78134 180668 78140
rect 181442 78160 181498 78169
rect 180064 77716 180116 77722
rect 180064 77658 180116 77664
rect 180076 74050 180104 77658
rect 180064 74044 180116 74050
rect 180064 73986 180116 73992
rect 180168 70394 180196 78134
rect 180432 77852 180484 77858
rect 180432 77794 180484 77800
rect 180340 77784 180392 77790
rect 180340 77726 180392 77732
rect 180352 75138 180380 77726
rect 180444 76362 180472 77794
rect 180628 77518 180656 78134
rect 180708 78124 180760 78130
rect 181442 78095 181498 78104
rect 180708 78066 180760 78072
rect 180616 77512 180668 77518
rect 180616 77454 180668 77460
rect 180432 76356 180484 76362
rect 180432 76298 180484 76304
rect 180340 75132 180392 75138
rect 180340 75074 180392 75080
rect 180076 70366 180196 70394
rect 180352 70394 180380 75074
rect 180628 72706 180656 77454
rect 180720 73166 180748 78066
rect 181640 77994 181668 78503
rect 183756 78266 183784 79698
rect 183744 78260 183796 78266
rect 183744 78202 183796 78208
rect 184204 78260 184256 78266
rect 184204 78202 184256 78208
rect 181628 77988 181680 77994
rect 181628 77930 181680 77936
rect 182088 77988 182140 77994
rect 182088 77930 182140 77936
rect 180800 74724 180852 74730
rect 180800 74666 180852 74672
rect 180708 73160 180760 73166
rect 180708 73102 180760 73108
rect 180628 72678 180748 72706
rect 180352 70366 180656 70394
rect 180076 6458 180104 70366
rect 180064 6452 180116 6458
rect 180064 6394 180116 6400
rect 180628 3738 180656 70366
rect 180616 3732 180668 3738
rect 180616 3674 180668 3680
rect 180720 3670 180748 72678
rect 180812 16574 180840 74666
rect 181996 74044 182048 74050
rect 181996 73986 182048 73992
rect 182008 73642 182036 73986
rect 181996 73636 182048 73642
rect 181996 73578 182048 73584
rect 180812 16546 181024 16574
rect 180708 3664 180760 3670
rect 180708 3606 180760 3612
rect 179512 3596 179564 3602
rect 179512 3538 179564 3544
rect 179052 3460 179104 3466
rect 179432 3454 180288 3482
rect 179052 3402 179104 3408
rect 180260 480 180288 3454
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 182008 4146 182036 73578
rect 182100 6390 182128 77930
rect 183558 77480 183614 77489
rect 183558 77415 183614 77424
rect 182824 76696 182876 76702
rect 182824 76638 182876 76644
rect 182180 76560 182232 76566
rect 182180 76502 182232 76508
rect 182088 6384 182140 6390
rect 182088 6326 182140 6332
rect 181996 4140 182048 4146
rect 181996 4082 182048 4088
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 76502
rect 182836 4078 182864 76638
rect 183572 75070 183600 77415
rect 183560 75064 183612 75070
rect 183560 75006 183612 75012
rect 182916 69692 182968 69698
rect 182916 69634 182968 69640
rect 182824 4072 182876 4078
rect 182824 4014 182876 4020
rect 182928 3058 182956 69634
rect 183560 64184 183612 64190
rect 183560 64126 183612 64132
rect 183572 16574 183600 64126
rect 183572 16546 183784 16574
rect 182916 3052 182968 3058
rect 182916 2994 182968 3000
rect 183756 480 183784 16546
rect 184216 6914 184244 78202
rect 184848 75064 184900 75070
rect 184848 75006 184900 75012
rect 184296 71120 184348 71126
rect 184296 71062 184348 71068
rect 184124 6886 184244 6914
rect 184124 3806 184152 6886
rect 184112 3800 184164 3806
rect 184112 3742 184164 3748
rect 184308 3398 184336 71062
rect 184860 28286 184888 75006
rect 185032 74996 185084 75002
rect 185032 74938 185084 74944
rect 184848 28280 184900 28286
rect 184848 28222 184900 28228
rect 185044 6914 185072 74938
rect 186976 65958 187004 80038
rect 186964 65952 187016 65958
rect 186964 65894 187016 65900
rect 187068 65822 187096 80310
rect 188356 66978 188384 80446
rect 188436 80436 188488 80442
rect 188436 80378 188488 80384
rect 188344 66972 188396 66978
rect 188344 66914 188396 66920
rect 188448 66910 188476 80378
rect 188908 80345 188936 82758
rect 188988 82136 189040 82142
rect 188988 82078 189040 82084
rect 188894 80336 188950 80345
rect 188894 80271 188950 80280
rect 189000 78577 189028 82078
rect 188986 78568 189042 78577
rect 188986 78503 189042 78512
rect 189080 72752 189132 72758
rect 189080 72694 189132 72700
rect 189092 72554 189120 72694
rect 189080 72548 189132 72554
rect 189080 72490 189132 72496
rect 188436 66904 188488 66910
rect 188436 66846 188488 66852
rect 187056 65816 187108 65822
rect 187056 65758 187108 65764
rect 188342 65512 188398 65521
rect 188342 65447 188398 65456
rect 185584 61396 185636 61402
rect 185584 61338 185636 61344
rect 184952 6886 185072 6914
rect 184296 3392 184348 3398
rect 184296 3334 184348 3340
rect 184952 480 184980 6886
rect 185596 3602 185624 61338
rect 187700 60036 187752 60042
rect 187700 59978 187752 59984
rect 187712 16574 187740 59978
rect 187712 16546 188292 16574
rect 187424 4140 187476 4146
rect 187424 4082 187476 4088
rect 187436 3602 187464 4082
rect 185584 3596 185636 3602
rect 185584 3538 185636 3544
rect 187332 3596 187384 3602
rect 187332 3538 187384 3544
rect 187424 3596 187476 3602
rect 187424 3538 187476 3544
rect 186136 3052 186188 3058
rect 186136 2994 186188 3000
rect 186148 480 186176 2994
rect 187344 480 187372 3538
rect 188264 3482 188292 16546
rect 188356 4146 188384 65447
rect 189080 60716 189132 60722
rect 189080 60658 189132 60664
rect 189092 60110 189120 60658
rect 189080 60104 189132 60110
rect 189080 60046 189132 60052
rect 189184 59106 189212 140286
rect 189368 60722 189396 144026
rect 189460 143177 189488 259927
rect 189552 143206 189580 260063
rect 189724 259752 189776 259758
rect 189724 259694 189776 259700
rect 189632 259616 189684 259622
rect 189632 259558 189684 259564
rect 189644 145518 189672 259558
rect 189736 146742 189764 259694
rect 190472 199510 190500 262550
rect 190552 262268 190604 262274
rect 190552 262210 190604 262216
rect 190460 199504 190512 199510
rect 190460 199446 190512 199452
rect 190564 199442 190592 262210
rect 190552 199436 190604 199442
rect 190552 199378 190604 199384
rect 190460 199300 190512 199306
rect 190460 199242 190512 199248
rect 189816 165640 189868 165646
rect 189816 165582 189868 165588
rect 189724 146736 189776 146742
rect 189724 146678 189776 146684
rect 189632 145512 189684 145518
rect 189632 145454 189684 145460
rect 189828 144294 189856 165582
rect 190092 146804 190144 146810
rect 190092 146746 190144 146752
rect 190000 146668 190052 146674
rect 190000 146610 190052 146616
rect 189816 144288 189868 144294
rect 189816 144230 189868 144236
rect 189632 143540 189684 143546
rect 189632 143482 189684 143488
rect 189540 143200 189592 143206
rect 189446 143168 189502 143177
rect 189540 143142 189592 143148
rect 189446 143103 189502 143112
rect 189448 139868 189500 139874
rect 189448 139810 189500 139816
rect 189460 69834 189488 139810
rect 189538 110664 189594 110673
rect 189538 110599 189594 110608
rect 189552 107137 189580 110599
rect 189538 107128 189594 107137
rect 189538 107063 189594 107072
rect 189644 72758 189672 143482
rect 189908 141704 189960 141710
rect 189908 141646 189960 141652
rect 189724 114572 189776 114578
rect 189724 114514 189776 114520
rect 189736 72826 189764 114514
rect 189920 113898 189948 141646
rect 190012 140078 190040 146610
rect 190000 140072 190052 140078
rect 190000 140014 190052 140020
rect 190000 138032 190052 138038
rect 190000 137974 190052 137980
rect 190012 114442 190040 137974
rect 190000 114436 190052 114442
rect 190000 114378 190052 114384
rect 189908 113892 189960 113898
rect 189908 113834 189960 113840
rect 189816 113756 189868 113762
rect 189816 113698 189868 113704
rect 189828 74390 189856 113698
rect 190104 80102 190132 146746
rect 190184 145648 190236 145654
rect 190184 145590 190236 145596
rect 190092 80096 190144 80102
rect 190092 80038 190144 80044
rect 189816 74384 189868 74390
rect 189816 74326 189868 74332
rect 189724 72820 189776 72826
rect 189724 72762 189776 72768
rect 189632 72752 189684 72758
rect 189632 72694 189684 72700
rect 189448 69828 189500 69834
rect 189448 69770 189500 69776
rect 189724 68332 189776 68338
rect 189724 68274 189776 68280
rect 189356 60716 189408 60722
rect 189356 60658 189408 60664
rect 189092 59078 189212 59106
rect 189092 56302 189120 59078
rect 189080 56296 189132 56302
rect 189080 56238 189132 56244
rect 189092 56166 189120 56238
rect 189080 56160 189132 56166
rect 189080 56102 189132 56108
rect 189632 52420 189684 52426
rect 189632 52362 189684 52368
rect 189644 52057 189672 52362
rect 189630 52048 189686 52057
rect 189630 51983 189686 51992
rect 189644 51134 189672 51983
rect 189632 51128 189684 51134
rect 189632 51070 189684 51076
rect 189448 49700 189500 49706
rect 189448 49642 189500 49648
rect 189460 49026 189488 49642
rect 189448 49020 189500 49026
rect 189448 48962 189500 48968
rect 189736 16574 189764 68274
rect 190196 49026 190224 145590
rect 190472 57798 190500 199242
rect 190656 141982 190684 263842
rect 190736 263764 190788 263770
rect 190736 263706 190788 263712
rect 190748 143138 190776 263706
rect 190828 262336 190880 262342
rect 190828 262278 190880 262284
rect 190736 143132 190788 143138
rect 190736 143074 190788 143080
rect 190840 142526 190868 262278
rect 192116 260976 192168 260982
rect 192116 260918 192168 260924
rect 190920 259956 190972 259962
rect 190920 259898 190972 259904
rect 190828 142520 190880 142526
rect 190828 142462 190880 142468
rect 190644 141976 190696 141982
rect 190644 141918 190696 141924
rect 190932 141778 190960 259898
rect 191010 259856 191066 259865
rect 191010 259791 191066 259800
rect 191024 143041 191052 259791
rect 191564 200320 191616 200326
rect 191564 200262 191616 200268
rect 191380 152720 191432 152726
rect 191380 152662 191432 152668
rect 191288 150340 191340 150346
rect 191288 150282 191340 150288
rect 191010 143032 191066 143041
rect 191010 142967 191066 142976
rect 191104 142996 191156 143002
rect 191104 142938 191156 142944
rect 190920 141772 190972 141778
rect 190920 141714 190972 141720
rect 190828 141568 190880 141574
rect 190828 141510 190880 141516
rect 190840 72962 190868 141510
rect 191012 140208 191064 140214
rect 191012 140150 191064 140156
rect 190920 140072 190972 140078
rect 190920 140014 190972 140020
rect 190828 72956 190880 72962
rect 190828 72898 190880 72904
rect 190932 72214 190960 140014
rect 191024 80578 191052 140150
rect 191116 114578 191144 142938
rect 191196 140004 191248 140010
rect 191196 139946 191248 139952
rect 191208 118726 191236 139946
rect 191300 138174 191328 150282
rect 191288 138168 191340 138174
rect 191288 138110 191340 138116
rect 191196 118720 191248 118726
rect 191196 118662 191248 118668
rect 191104 114572 191156 114578
rect 191104 114514 191156 114520
rect 191196 113892 191248 113898
rect 191196 113834 191248 113840
rect 191012 80572 191064 80578
rect 191012 80514 191064 80520
rect 190920 72208 190972 72214
rect 190920 72150 190972 72156
rect 191208 71602 191236 113834
rect 191286 109168 191342 109177
rect 191286 109103 191342 109112
rect 191300 80238 191328 109103
rect 191288 80232 191340 80238
rect 191288 80174 191340 80180
rect 191288 79348 191340 79354
rect 191288 79290 191340 79296
rect 191196 71596 191248 71602
rect 191196 71538 191248 71544
rect 191300 65890 191328 79290
rect 191392 70922 191420 152662
rect 191472 144424 191524 144430
rect 191472 144366 191524 144372
rect 191484 72622 191512 144366
rect 191576 78538 191604 200262
rect 192024 197124 192076 197130
rect 192024 197066 192076 197072
rect 191840 143064 191892 143070
rect 191840 143006 191892 143012
rect 191852 114594 191880 143006
rect 191932 118720 191984 118726
rect 191932 118662 191984 118668
rect 191668 114566 191880 114594
rect 191564 78532 191616 78538
rect 191564 78474 191616 78480
rect 191472 72616 191524 72622
rect 191472 72558 191524 72564
rect 191668 71534 191696 114566
rect 191944 113762 191972 118662
rect 191932 113756 191984 113762
rect 191932 113698 191984 113704
rect 191932 80232 191984 80238
rect 191932 80174 191984 80180
rect 191748 78532 191800 78538
rect 191748 78474 191800 78480
rect 191760 77994 191788 78474
rect 191748 77988 191800 77994
rect 191748 77930 191800 77936
rect 191656 71528 191708 71534
rect 191656 71470 191708 71476
rect 191380 70916 191432 70922
rect 191380 70858 191432 70864
rect 191288 65884 191340 65890
rect 191288 65826 191340 65832
rect 190460 57792 190512 57798
rect 190460 57734 190512 57740
rect 191748 57792 191800 57798
rect 191748 57734 191800 57740
rect 191760 57390 191788 57734
rect 191748 57384 191800 57390
rect 191748 57326 191800 57332
rect 190184 49020 190236 49026
rect 190184 48962 190236 48968
rect 191838 43480 191894 43489
rect 191838 43415 191894 43424
rect 191852 16574 191880 43415
rect 191944 39953 191972 80174
rect 192036 63374 192064 197066
rect 192128 139534 192156 260918
rect 192220 145858 192248 264998
rect 193772 263696 193824 263702
rect 193772 263638 193824 263644
rect 192392 262948 192444 262954
rect 192392 262890 192444 262896
rect 192298 260264 192354 260273
rect 192298 260199 192354 260208
rect 192208 145852 192260 145858
rect 192208 145794 192260 145800
rect 192208 145716 192260 145722
rect 192208 145658 192260 145664
rect 192116 139528 192168 139534
rect 192116 139470 192168 139476
rect 192220 73982 192248 145658
rect 192312 141642 192340 260199
rect 192404 144702 192432 262890
rect 193680 261248 193732 261254
rect 193680 261190 193732 261196
rect 192484 260228 192536 260234
rect 192484 260170 192536 260176
rect 192392 144696 192444 144702
rect 192392 144638 192444 144644
rect 192496 144566 192524 260170
rect 192576 259684 192628 259690
rect 192576 259626 192628 259632
rect 192588 153270 192616 259626
rect 193404 200252 193456 200258
rect 193404 200194 193456 200200
rect 192760 199368 192812 199374
rect 192760 199310 192812 199316
rect 192668 195764 192720 195770
rect 192668 195706 192720 195712
rect 192576 153264 192628 153270
rect 192576 153206 192628 153212
rect 192576 145988 192628 145994
rect 192576 145930 192628 145936
rect 192484 144560 192536 144566
rect 192484 144502 192536 144508
rect 192392 143812 192444 143818
rect 192392 143754 192444 143760
rect 192300 141636 192352 141642
rect 192300 141578 192352 141584
rect 192300 139936 192352 139942
rect 192300 139878 192352 139884
rect 192312 75614 192340 139878
rect 192404 80510 192432 143754
rect 192484 139324 192536 139330
rect 192484 139266 192536 139272
rect 192496 80646 192524 139266
rect 192588 122126 192616 145930
rect 192576 122120 192628 122126
rect 192576 122062 192628 122068
rect 192576 114436 192628 114442
rect 192576 114378 192628 114384
rect 192484 80640 192536 80646
rect 192484 80582 192536 80588
rect 192392 80504 192444 80510
rect 192392 80446 192444 80452
rect 192300 75608 192352 75614
rect 192300 75550 192352 75556
rect 192208 73976 192260 73982
rect 192208 73918 192260 73924
rect 192482 72448 192538 72457
rect 192482 72383 192538 72392
rect 192496 71602 192524 72383
rect 192484 71596 192536 71602
rect 192484 71538 192536 71544
rect 192588 67454 192616 114378
rect 192576 67448 192628 67454
rect 192576 67390 192628 67396
rect 192024 63368 192076 63374
rect 192024 63310 192076 63316
rect 192680 51066 192708 195706
rect 192772 59294 192800 199310
rect 193312 196988 193364 196994
rect 193312 196930 193364 196936
rect 193220 195560 193272 195566
rect 193220 195502 193272 195508
rect 192852 139868 192904 139874
rect 192852 139810 192904 139816
rect 192864 71670 192892 139810
rect 192852 71664 192904 71670
rect 192852 71606 192904 71612
rect 193128 71596 193180 71602
rect 193128 71538 193180 71544
rect 193036 67448 193088 67454
rect 193036 67390 193088 67396
rect 193048 66978 193076 67390
rect 193036 66972 193088 66978
rect 193036 66914 193088 66920
rect 193036 63368 193088 63374
rect 193036 63310 193088 63316
rect 193048 62830 193076 63310
rect 193036 62824 193088 62830
rect 193036 62766 193088 62772
rect 192760 59288 192812 59294
rect 192760 59230 192812 59236
rect 193036 59288 193088 59294
rect 193036 59230 193088 59236
rect 193048 58750 193076 59230
rect 193036 58744 193088 58750
rect 193036 58686 193088 58692
rect 192668 51060 192720 51066
rect 192668 51002 192720 51008
rect 193036 51060 193088 51066
rect 193036 51002 193088 51008
rect 193048 50454 193076 51002
rect 193036 50448 193088 50454
rect 193036 50390 193088 50396
rect 191930 39944 191986 39953
rect 191930 39879 191986 39888
rect 193034 39944 193090 39953
rect 193034 39879 193090 39888
rect 193048 39273 193076 39879
rect 193034 39264 193090 39273
rect 193034 39199 193090 39208
rect 189736 16546 189856 16574
rect 191852 16546 192064 16574
rect 188344 4140 188396 4146
rect 188344 4082 188396 4088
rect 188264 3454 188568 3482
rect 188540 480 188568 3454
rect 189828 3398 189856 16546
rect 190828 3528 190880 3534
rect 190828 3470 190880 3476
rect 189724 3392 189776 3398
rect 189724 3334 189776 3340
rect 189816 3392 189868 3398
rect 189816 3334 189868 3340
rect 189736 480 189764 3334
rect 190840 480 190868 3470
rect 192036 480 192064 16546
rect 193140 3330 193168 71538
rect 193232 56370 193260 195502
rect 193324 60654 193352 196930
rect 193416 64802 193444 200194
rect 193496 196920 193548 196926
rect 193496 196862 193548 196868
rect 193508 69766 193536 196862
rect 193588 146260 193640 146266
rect 193588 146202 193640 146208
rect 193496 69760 193548 69766
rect 193496 69702 193548 69708
rect 193404 64796 193456 64802
rect 193404 64738 193456 64744
rect 193416 64326 193444 64738
rect 193404 64320 193456 64326
rect 193404 64262 193456 64268
rect 193312 60648 193364 60654
rect 193312 60590 193364 60596
rect 193220 56364 193272 56370
rect 193220 56306 193272 56312
rect 193600 52193 193628 146202
rect 193692 141370 193720 261190
rect 193784 144362 193812 263638
rect 193956 263220 194008 263226
rect 193956 263162 194008 263168
rect 193864 260092 193916 260098
rect 193864 260034 193916 260040
rect 193772 144356 193824 144362
rect 193772 144298 193824 144304
rect 193876 141914 193904 260034
rect 193968 146198 193996 263162
rect 194048 262812 194100 262818
rect 194048 262754 194100 262760
rect 193956 146192 194008 146198
rect 193956 146134 194008 146140
rect 193956 142044 194008 142050
rect 193956 141986 194008 141992
rect 193864 141908 193916 141914
rect 193864 141850 193916 141856
rect 193680 141364 193732 141370
rect 193680 141306 193732 141312
rect 193680 140752 193732 140758
rect 193678 140720 193680 140729
rect 193732 140720 193734 140729
rect 193678 140655 193734 140664
rect 193772 140276 193824 140282
rect 193772 140218 193824 140224
rect 193784 68406 193812 140218
rect 193862 139360 193918 139369
rect 193862 139295 193918 139304
rect 193876 71466 193904 139295
rect 193968 72554 193996 141986
rect 194060 141409 194088 262754
rect 194598 197160 194654 197169
rect 194598 197095 194654 197104
rect 194232 146056 194284 146062
rect 194232 145998 194284 146004
rect 194046 141400 194102 141409
rect 194046 141335 194102 141344
rect 194046 140040 194102 140049
rect 194046 139975 194102 139984
rect 194060 77722 194088 139975
rect 194048 77716 194100 77722
rect 194048 77658 194100 77664
rect 194046 75168 194102 75177
rect 194046 75103 194102 75112
rect 193956 72548 194008 72554
rect 193956 72490 194008 72496
rect 193864 71460 193916 71466
rect 193864 71402 193916 71408
rect 193772 68400 193824 68406
rect 193772 68342 193824 68348
rect 193678 60616 193734 60625
rect 193678 60551 193680 60560
rect 193732 60551 193734 60560
rect 193680 60522 193732 60528
rect 193586 52184 193642 52193
rect 193586 52119 193642 52128
rect 193310 50280 193366 50289
rect 193310 50215 193366 50224
rect 193324 16574 193352 50215
rect 193324 16546 193996 16574
rect 193864 4140 193916 4146
rect 193864 4082 193916 4088
rect 193876 3534 193904 4082
rect 193864 3528 193916 3534
rect 193864 3470 193916 3476
rect 193968 3482 193996 16546
rect 194060 4146 194088 75103
rect 194244 72146 194272 145998
rect 194508 144832 194560 144838
rect 194508 144774 194560 144780
rect 194520 138145 194548 144774
rect 194506 138136 194562 138145
rect 194506 138071 194562 138080
rect 194232 72140 194284 72146
rect 194232 72082 194284 72088
rect 194508 60648 194560 60654
rect 194508 60590 194560 60596
rect 194416 60580 194468 60586
rect 194416 60522 194468 60528
rect 194428 59430 194456 60522
rect 194520 60042 194548 60590
rect 194508 60036 194560 60042
rect 194508 59978 194560 59984
rect 194416 59424 194468 59430
rect 194416 59366 194468 59372
rect 194508 56364 194560 56370
rect 194508 56306 194560 56312
rect 194520 56098 194548 56306
rect 194508 56092 194560 56098
rect 194508 56034 194560 56040
rect 194612 54913 194640 197095
rect 194692 195424 194744 195430
rect 194692 195366 194744 195372
rect 194704 57866 194732 195366
rect 194796 139670 194824 265134
rect 194888 144158 194916 265610
rect 196256 265600 196308 265606
rect 196256 265542 196308 265548
rect 196164 265464 196216 265470
rect 196164 265406 196216 265412
rect 194968 262472 195020 262478
rect 194968 262414 195020 262420
rect 194980 146130 195008 262414
rect 195060 261180 195112 261186
rect 195060 261122 195112 261128
rect 195072 150414 195100 261122
rect 195978 195800 196034 195809
rect 195978 195735 196034 195744
rect 195426 152688 195482 152697
rect 195426 152623 195482 152632
rect 195060 150408 195112 150414
rect 195060 150350 195112 150356
rect 195060 149048 195112 149054
rect 195060 148990 195112 148996
rect 194968 146124 195020 146130
rect 194968 146066 195020 146072
rect 194876 144152 194928 144158
rect 194876 144094 194928 144100
rect 194784 139664 194836 139670
rect 194784 139606 194836 139612
rect 195072 70378 195100 148990
rect 195152 148504 195204 148510
rect 195152 148446 195204 148452
rect 195164 80374 195192 148446
rect 195242 139224 195298 139233
rect 195242 139159 195298 139168
rect 195152 80368 195204 80374
rect 195152 80310 195204 80316
rect 195256 77858 195284 139159
rect 195336 138916 195388 138922
rect 195336 138858 195388 138864
rect 195348 80442 195376 138858
rect 195440 124914 195468 152623
rect 195612 148844 195664 148850
rect 195612 148786 195664 148792
rect 195518 145616 195574 145625
rect 195518 145551 195574 145560
rect 195428 124908 195480 124914
rect 195428 124850 195480 124856
rect 195336 80436 195388 80442
rect 195336 80378 195388 80384
rect 195244 77852 195296 77858
rect 195244 77794 195296 77800
rect 195532 71194 195560 145551
rect 195624 71262 195652 148786
rect 195704 147348 195756 147354
rect 195704 147290 195756 147296
rect 195716 76362 195744 147290
rect 195704 76356 195756 76362
rect 195704 76298 195756 76304
rect 195612 71256 195664 71262
rect 195612 71198 195664 71204
rect 195520 71188 195572 71194
rect 195520 71130 195572 71136
rect 195060 70372 195112 70378
rect 195060 70314 195112 70320
rect 195072 69698 195100 70314
rect 195060 69692 195112 69698
rect 195060 69634 195112 69640
rect 194692 57860 194744 57866
rect 194692 57802 194744 57808
rect 195060 57860 195112 57866
rect 195060 57802 195112 57808
rect 195072 57322 195100 57802
rect 195060 57316 195112 57322
rect 195060 57258 195112 57264
rect 194598 54904 194654 54913
rect 194598 54839 194654 54848
rect 194612 54641 194640 54839
rect 194598 54632 194654 54641
rect 194598 54567 194654 54576
rect 195992 49473 196020 195735
rect 196072 195696 196124 195702
rect 196072 195638 196124 195644
rect 196084 53689 196112 195638
rect 196176 144770 196204 265406
rect 196268 144906 196296 265542
rect 197360 265532 197412 265538
rect 197360 265474 197412 265480
rect 196440 261044 196492 261050
rect 196440 260986 196492 260992
rect 196348 260908 196400 260914
rect 196348 260850 196400 260856
rect 196256 144900 196308 144906
rect 196256 144842 196308 144848
rect 196164 144764 196216 144770
rect 196164 144706 196216 144712
rect 196360 143274 196388 260850
rect 196452 147626 196480 260986
rect 196624 259820 196676 259826
rect 196624 259762 196676 259768
rect 196532 259480 196584 259486
rect 196532 259422 196584 259428
rect 196440 147620 196492 147626
rect 196440 147562 196492 147568
rect 196544 145586 196572 259422
rect 196636 157894 196664 259762
rect 196624 157888 196676 157894
rect 196624 157830 196676 157836
rect 196900 148776 196952 148782
rect 196900 148718 196952 148724
rect 196714 146976 196770 146985
rect 196714 146911 196770 146920
rect 196532 145580 196584 145586
rect 196532 145522 196584 145528
rect 196348 143268 196400 143274
rect 196348 143210 196400 143216
rect 196532 141296 196584 141302
rect 196532 141238 196584 141244
rect 196440 138848 196492 138854
rect 196440 138790 196492 138796
rect 196162 82240 196218 82249
rect 196162 82175 196218 82184
rect 196176 82142 196204 82175
rect 196164 82136 196216 82142
rect 196164 82078 196216 82084
rect 196164 76968 196216 76974
rect 196164 76910 196216 76916
rect 196176 76566 196204 76910
rect 196164 76560 196216 76566
rect 196164 76502 196216 76508
rect 196452 70242 196480 138790
rect 196544 72690 196572 141238
rect 196622 138680 196678 138689
rect 196622 138615 196678 138624
rect 196532 72684 196584 72690
rect 196532 72626 196584 72632
rect 196636 72350 196664 138615
rect 196728 80714 196756 146911
rect 196806 113928 196862 113937
rect 196806 113863 196862 113872
rect 196716 80708 196768 80714
rect 196716 80650 196768 80656
rect 196820 76566 196848 113863
rect 196808 76560 196860 76566
rect 196808 76502 196860 76508
rect 196624 72344 196676 72350
rect 196624 72286 196676 72292
rect 196440 70236 196492 70242
rect 196440 70178 196492 70184
rect 196624 69896 196676 69902
rect 196624 69838 196676 69844
rect 196164 67244 196216 67250
rect 196164 67186 196216 67192
rect 196176 66910 196204 67186
rect 196164 66904 196216 66910
rect 196164 66846 196216 66852
rect 196070 53680 196126 53689
rect 196070 53615 196126 53624
rect 195978 49464 196034 49473
rect 195978 49399 196034 49408
rect 195992 49201 196020 49399
rect 195978 49192 196034 49201
rect 195978 49127 196034 49136
rect 196636 4146 196664 69838
rect 196912 66910 196940 148718
rect 197372 146878 197400 265474
rect 199016 265396 199068 265402
rect 199016 265338 199068 265344
rect 198004 265260 198056 265266
rect 198004 265202 198056 265208
rect 197912 265124 197964 265130
rect 197912 265066 197964 265072
rect 197820 261384 197872 261390
rect 197820 261326 197872 261332
rect 197728 197260 197780 197266
rect 197728 197202 197780 197208
rect 197450 197024 197506 197033
rect 197450 196959 197506 196968
rect 197360 146872 197412 146878
rect 197360 146814 197412 146820
rect 196992 145920 197044 145926
rect 196992 145862 197044 145868
rect 197004 69970 197032 145862
rect 197084 145784 197136 145790
rect 197084 145726 197136 145732
rect 197096 70174 197124 145726
rect 197268 79416 197320 79422
rect 197268 79358 197320 79364
rect 197360 79416 197412 79422
rect 197360 79358 197412 79364
rect 197280 77874 197308 79358
rect 197372 78033 197400 79358
rect 197358 78024 197414 78033
rect 197358 77959 197414 77968
rect 197280 77846 197400 77874
rect 197084 70168 197136 70174
rect 197084 70110 197136 70116
rect 196992 69964 197044 69970
rect 196992 69906 197044 69912
rect 196900 66904 196952 66910
rect 196900 66846 196952 66852
rect 197372 16574 197400 77846
rect 197464 52562 197492 196959
rect 197636 196852 197688 196858
rect 197636 196794 197688 196800
rect 197544 196784 197596 196790
rect 197544 196726 197596 196732
rect 197452 52556 197504 52562
rect 197452 52498 197504 52504
rect 197450 52456 197506 52465
rect 197556 52442 197584 196726
rect 197648 62898 197676 196794
rect 197636 62892 197688 62898
rect 197636 62834 197688 62840
rect 197740 62778 197768 197202
rect 197832 147422 197860 261326
rect 197924 158710 197952 265066
rect 197912 158704 197964 158710
rect 197912 158646 197964 158652
rect 198016 157962 198044 265202
rect 198738 197296 198794 197305
rect 198738 197231 198794 197240
rect 198004 157956 198056 157962
rect 198004 157898 198056 157904
rect 198372 148912 198424 148918
rect 198372 148854 198424 148860
rect 197820 147416 197872 147422
rect 197820 147358 197872 147364
rect 197912 146940 197964 146946
rect 197912 146882 197964 146888
rect 197818 138952 197874 138961
rect 197818 138887 197874 138896
rect 197832 68474 197860 138887
rect 197924 86834 197952 146882
rect 198004 141228 198056 141234
rect 198004 141170 198056 141176
rect 197912 86828 197964 86834
rect 197912 86770 197964 86776
rect 198016 86714 198044 141170
rect 198188 138168 198240 138174
rect 198188 138110 198240 138116
rect 198094 114472 198150 114481
rect 198094 114407 198150 114416
rect 197924 86686 198044 86714
rect 197924 79082 197952 86686
rect 198004 86624 198056 86630
rect 198004 86566 198056 86572
rect 197912 79076 197964 79082
rect 197912 79018 197964 79024
rect 197910 78568 197966 78577
rect 197910 78503 197966 78512
rect 197924 78470 197952 78503
rect 197912 78464 197964 78470
rect 197912 78406 197964 78412
rect 197924 77382 197952 78406
rect 198016 77926 198044 86566
rect 198004 77920 198056 77926
rect 198004 77862 198056 77868
rect 197912 77376 197964 77382
rect 197912 77318 197964 77324
rect 198004 76628 198056 76634
rect 198004 76570 198056 76576
rect 197820 68468 197872 68474
rect 197820 68410 197872 68416
rect 197820 62892 197872 62898
rect 197820 62834 197872 62840
rect 197648 62750 197768 62778
rect 197648 62014 197676 62750
rect 197636 62008 197688 62014
rect 197636 61950 197688 61956
rect 197648 61470 197676 61950
rect 197636 61464 197688 61470
rect 197636 61406 197688 61412
rect 197832 61282 197860 62834
rect 197648 61254 197860 61282
rect 197648 56438 197676 61254
rect 197636 56432 197688 56438
rect 197636 56374 197688 56380
rect 197648 56030 197676 56374
rect 197636 56024 197688 56030
rect 197636 55966 197688 55972
rect 197636 52556 197688 52562
rect 197636 52498 197688 52504
rect 197506 52414 197584 52442
rect 197450 52391 197506 52400
rect 197464 52057 197492 52391
rect 197450 52048 197506 52057
rect 197450 51983 197506 51992
rect 197450 48104 197506 48113
rect 197648 48090 197676 52498
rect 197506 48062 197676 48090
rect 197450 48039 197506 48048
rect 197464 47841 197492 48039
rect 197450 47832 197506 47841
rect 197450 47767 197506 47776
rect 197372 16546 197952 16574
rect 194048 4140 194100 4146
rect 194048 4082 194100 4088
rect 195612 4140 195664 4146
rect 195612 4082 195664 4088
rect 196624 4140 196676 4146
rect 196624 4082 196676 4088
rect 193968 3454 194456 3482
rect 193220 3392 193272 3398
rect 193220 3334 193272 3340
rect 193128 3324 193180 3330
rect 193128 3266 193180 3272
rect 193232 480 193260 3334
rect 194428 480 194456 3454
rect 195624 480 195652 4082
rect 196808 3528 196860 3534
rect 196808 3470 196860 3476
rect 196820 480 196848 3470
rect 197924 480 197952 16546
rect 198016 3534 198044 76570
rect 198108 53718 198136 114407
rect 198200 79354 198228 138110
rect 198188 79348 198240 79354
rect 198188 79290 198240 79296
rect 198384 69562 198412 148854
rect 198372 69556 198424 69562
rect 198372 69498 198424 69504
rect 198096 53712 198148 53718
rect 198096 53654 198148 53660
rect 198108 53174 198136 53654
rect 198096 53168 198148 53174
rect 198096 53110 198148 53116
rect 198752 50697 198780 197231
rect 198832 197192 198884 197198
rect 198832 197134 198884 197140
rect 198844 55214 198872 197134
rect 198924 195492 198976 195498
rect 198924 195434 198976 195440
rect 198936 66094 198964 195434
rect 199028 139738 199056 265338
rect 199200 265328 199252 265334
rect 199200 265270 199252 265276
rect 199108 261112 199160 261118
rect 199108 261054 199160 261060
rect 199120 142118 199148 261054
rect 199212 147558 199240 265270
rect 203248 264988 203300 264994
rect 203248 264930 203300 264936
rect 199292 263832 199344 263838
rect 199292 263774 199344 263780
rect 199200 147552 199252 147558
rect 199200 147494 199252 147500
rect 199304 147490 199332 263774
rect 200580 260160 200632 260166
rect 200580 260102 200632 260108
rect 200120 198620 200172 198626
rect 200120 198562 200172 198568
rect 199476 151428 199528 151434
rect 199476 151370 199528 151376
rect 199292 147484 199344 147490
rect 199292 147426 199344 147432
rect 199292 147280 199344 147286
rect 199292 147222 199344 147228
rect 199108 142112 199160 142118
rect 199108 142054 199160 142060
rect 199016 139732 199068 139738
rect 199016 139674 199068 139680
rect 199106 139088 199162 139097
rect 199106 139023 199162 139032
rect 199014 78568 199070 78577
rect 199014 78503 199070 78512
rect 199028 78402 199056 78503
rect 199016 78396 199068 78402
rect 199016 78338 199068 78344
rect 199028 77314 199056 78338
rect 199016 77308 199068 77314
rect 199016 77250 199068 77256
rect 198924 66088 198976 66094
rect 198924 66030 198976 66036
rect 198936 65550 198964 66030
rect 198924 65544 198976 65550
rect 198924 65486 198976 65492
rect 199120 62121 199148 139023
rect 199304 76430 199332 147222
rect 199384 138780 199436 138786
rect 199384 138722 199436 138728
rect 199292 76424 199344 76430
rect 199292 76366 199344 76372
rect 199396 70038 199424 138722
rect 199488 81569 199516 151370
rect 199752 148708 199804 148714
rect 199752 148650 199804 148656
rect 199660 148300 199712 148306
rect 199660 148242 199712 148248
rect 199566 138816 199622 138825
rect 199566 138751 199622 138760
rect 199474 81560 199530 81569
rect 199474 81495 199530 81504
rect 199580 71398 199608 138751
rect 199568 71392 199620 71398
rect 199568 71334 199620 71340
rect 199384 70032 199436 70038
rect 199384 69974 199436 69980
rect 199672 67386 199700 148242
rect 199764 70106 199792 148650
rect 200132 79642 200160 198562
rect 200394 196752 200450 196761
rect 200394 196687 200450 196696
rect 200304 195832 200356 195838
rect 200304 195774 200356 195780
rect 200212 193180 200264 193186
rect 200212 193122 200264 193128
rect 200040 79614 200160 79642
rect 200040 79286 200068 79614
rect 200028 79280 200080 79286
rect 200028 79222 200080 79228
rect 200120 71052 200172 71058
rect 200120 70994 200172 71000
rect 199752 70100 199804 70106
rect 199752 70042 199804 70048
rect 199660 67380 199712 67386
rect 199660 67322 199712 67328
rect 199106 62112 199162 62121
rect 199106 62047 199162 62056
rect 199842 62112 199898 62121
rect 199842 62047 199898 62056
rect 199856 61577 199884 62047
rect 199842 61568 199898 61577
rect 199842 61503 199898 61512
rect 198832 55208 198884 55214
rect 198832 55150 198884 55156
rect 198844 54602 198872 55150
rect 198832 54596 198884 54602
rect 198832 54538 198884 54544
rect 198738 50688 198794 50697
rect 198738 50623 198794 50632
rect 198740 44872 198792 44878
rect 198740 44814 198792 44820
rect 198004 3528 198056 3534
rect 198004 3470 198056 3476
rect 198096 3460 198148 3466
rect 198096 3402 198148 3408
rect 198108 3330 198136 3402
rect 198096 3324 198148 3330
rect 198096 3266 198148 3272
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 44814
rect 200132 16574 200160 70994
rect 200224 45393 200252 193122
rect 200316 57769 200344 195774
rect 200408 63073 200436 196687
rect 200488 191208 200540 191214
rect 200488 191150 200540 191156
rect 200500 78198 200528 191150
rect 200592 155650 200620 260102
rect 202880 200388 202932 200394
rect 202880 200330 202932 200336
rect 201776 196716 201828 196722
rect 201776 196658 201828 196664
rect 201684 193112 201736 193118
rect 201684 193054 201736 193060
rect 201500 191276 201552 191282
rect 201500 191218 201552 191224
rect 201224 158568 201276 158574
rect 201224 158510 201276 158516
rect 200580 155644 200632 155650
rect 200580 155586 200632 155592
rect 200672 155440 200724 155446
rect 200672 155382 200724 155388
rect 200488 78192 200540 78198
rect 200488 78134 200540 78140
rect 200684 68814 200712 155382
rect 200764 155372 200816 155378
rect 200764 155314 200816 155320
rect 200776 74322 200804 155314
rect 200856 148436 200908 148442
rect 200856 148378 200908 148384
rect 200764 74316 200816 74322
rect 200764 74258 200816 74264
rect 200672 68808 200724 68814
rect 200672 68750 200724 68756
rect 200868 68134 200896 148378
rect 200946 137864 201002 137873
rect 200946 137799 201002 137808
rect 200960 72894 200988 137799
rect 200948 72888 201000 72894
rect 200948 72830 201000 72836
rect 201236 68678 201264 158510
rect 201314 80064 201370 80073
rect 201314 79999 201370 80008
rect 201328 79150 201356 79999
rect 201408 79484 201460 79490
rect 201408 79426 201460 79432
rect 201316 79144 201368 79150
rect 201316 79086 201368 79092
rect 201328 78742 201356 79086
rect 201316 78736 201368 78742
rect 201316 78678 201368 78684
rect 201420 78169 201448 79426
rect 201406 78160 201462 78169
rect 201406 78095 201462 78104
rect 201224 68672 201276 68678
rect 201224 68614 201276 68620
rect 200856 68128 200908 68134
rect 200856 68070 200908 68076
rect 201512 63306 201540 191218
rect 201500 63300 201552 63306
rect 201500 63242 201552 63248
rect 200394 63064 200450 63073
rect 200394 62999 200450 63008
rect 200302 57760 200358 57769
rect 200302 57695 200358 57704
rect 201696 52329 201724 193054
rect 201788 59362 201816 196658
rect 202420 192432 202472 192438
rect 202420 192374 202472 192380
rect 202328 190120 202380 190126
rect 202328 190062 202380 190068
rect 201866 158128 201922 158137
rect 201866 158063 201922 158072
rect 201776 59356 201828 59362
rect 201776 59298 201828 59304
rect 201880 56506 201908 158063
rect 201958 151056 202014 151065
rect 201958 150991 202014 151000
rect 201972 76838 202000 150991
rect 202052 148640 202104 148646
rect 202052 148582 202104 148588
rect 202064 78130 202092 148582
rect 202144 137828 202196 137834
rect 202144 137770 202196 137776
rect 202052 78124 202104 78130
rect 202052 78066 202104 78072
rect 201960 76832 202012 76838
rect 201960 76774 202012 76780
rect 201960 75200 202012 75206
rect 201960 75142 202012 75148
rect 201868 56500 201920 56506
rect 201868 56442 201920 56448
rect 201682 52320 201738 52329
rect 201682 52255 201738 52264
rect 201592 49156 201644 49162
rect 201592 49098 201644 49104
rect 200210 45384 200266 45393
rect 200210 45319 200266 45328
rect 201406 45384 201462 45393
rect 201406 45319 201462 45328
rect 201420 44985 201448 45319
rect 201406 44976 201462 44985
rect 201406 44911 201462 44920
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201604 2774 201632 49098
rect 201972 16574 202000 75142
rect 202156 71602 202184 137770
rect 202236 136740 202288 136746
rect 202236 136682 202288 136688
rect 202248 75818 202276 136682
rect 202340 136610 202368 190062
rect 202328 136604 202380 136610
rect 202328 136546 202380 136552
rect 202328 122120 202380 122126
rect 202328 122062 202380 122068
rect 202340 78334 202368 122062
rect 202328 78328 202380 78334
rect 202328 78270 202380 78276
rect 202236 75812 202288 75818
rect 202236 75754 202288 75760
rect 202144 71596 202196 71602
rect 202144 71538 202196 71544
rect 202432 49609 202460 192374
rect 202788 75812 202840 75818
rect 202788 75754 202840 75760
rect 202800 75274 202828 75754
rect 202788 75268 202840 75274
rect 202788 75210 202840 75216
rect 202788 59356 202840 59362
rect 202788 59298 202840 59304
rect 202800 58682 202828 59298
rect 202788 58676 202840 58682
rect 202788 58618 202840 58624
rect 202788 56500 202840 56506
rect 202788 56442 202840 56448
rect 202800 55962 202828 56442
rect 202788 55956 202840 55962
rect 202788 55898 202840 55904
rect 202892 55146 202920 200330
rect 203156 197056 203208 197062
rect 203156 196998 203208 197004
rect 203064 192976 203116 192982
rect 203064 192918 203116 192924
rect 202970 192808 203026 192817
rect 202970 192743 203026 192752
rect 202880 55140 202932 55146
rect 202880 55082 202932 55088
rect 202892 54534 202920 55082
rect 202880 54528 202932 54534
rect 202880 54470 202932 54476
rect 202786 52320 202842 52329
rect 202786 52255 202842 52264
rect 202800 51921 202828 52255
rect 202786 51912 202842 51921
rect 202786 51847 202842 51856
rect 202418 49600 202474 49609
rect 202418 49535 202474 49544
rect 202786 49600 202842 49609
rect 202786 49535 202842 49544
rect 202800 49065 202828 49535
rect 202786 49056 202842 49065
rect 202786 48991 202842 49000
rect 202984 47977 203012 192743
rect 203076 64734 203104 192918
rect 203168 73710 203196 196998
rect 203260 154018 203288 264930
rect 204812 264240 204864 264246
rect 204812 264182 204864 264188
rect 204824 263634 204852 264182
rect 204812 263628 204864 263634
rect 204812 263570 204864 263576
rect 204628 262676 204680 262682
rect 204628 262618 204680 262624
rect 203340 259888 203392 259894
rect 203340 259830 203392 259836
rect 203352 157826 203380 259830
rect 204260 193044 204312 193050
rect 204260 192986 204312 192992
rect 203432 158500 203484 158506
rect 203432 158442 203484 158448
rect 203340 157820 203392 157826
rect 203340 157762 203392 157768
rect 203338 155544 203394 155553
rect 203338 155479 203394 155488
rect 203248 154012 203300 154018
rect 203248 153954 203300 153960
rect 203246 148336 203302 148345
rect 203246 148271 203302 148280
rect 203156 73704 203208 73710
rect 203156 73646 203208 73652
rect 203064 64728 203116 64734
rect 203064 64670 203116 64676
rect 203076 64258 203104 64670
rect 203064 64252 203116 64258
rect 203064 64194 203116 64200
rect 203260 57934 203288 148271
rect 203248 57928 203300 57934
rect 203248 57870 203300 57876
rect 203352 48249 203380 155479
rect 203444 68746 203472 158442
rect 203524 151292 203576 151298
rect 203524 151234 203576 151240
rect 203536 71330 203564 151234
rect 203708 148572 203760 148578
rect 203708 148514 203760 148520
rect 203616 138712 203668 138718
rect 203616 138654 203668 138660
rect 203524 71324 203576 71330
rect 203524 71266 203576 71272
rect 203432 68740 203484 68746
rect 203432 68682 203484 68688
rect 203524 67108 203576 67114
rect 203524 67050 203576 67056
rect 203338 48240 203394 48249
rect 203338 48175 203394 48184
rect 202970 47968 203026 47977
rect 202970 47903 203026 47912
rect 201972 16546 202736 16574
rect 201512 2746 201632 2774
rect 201512 480 201540 2746
rect 202708 480 202736 16546
rect 203536 2922 203564 67050
rect 203628 63442 203656 138654
rect 203720 82822 203748 148514
rect 203708 82816 203760 82822
rect 203708 82758 203760 82764
rect 203616 63436 203668 63442
rect 203616 63378 203668 63384
rect 204168 57928 204220 57934
rect 204168 57870 204220 57876
rect 204180 57254 204208 57870
rect 204168 57248 204220 57254
rect 204168 57190 204220 57196
rect 204272 53786 204300 192986
rect 204444 192908 204496 192914
rect 204444 192850 204496 192856
rect 204352 192772 204404 192778
rect 204352 192714 204404 192720
rect 204364 70990 204392 192714
rect 204456 74186 204484 192850
rect 204536 192704 204588 192710
rect 204536 192646 204588 192652
rect 204548 75546 204576 192646
rect 204640 153950 204668 262618
rect 204824 258074 204852 263570
rect 206008 262744 206060 262750
rect 206008 262686 206060 262692
rect 204732 258046 204852 258074
rect 204732 158302 204760 258046
rect 205640 192840 205692 192846
rect 205640 192782 205692 192788
rect 204720 158296 204772 158302
rect 204720 158238 204772 158244
rect 204628 153944 204680 153950
rect 204628 153886 204680 153892
rect 204904 150272 204956 150278
rect 204904 150214 204956 150220
rect 204718 147112 204774 147121
rect 204718 147047 204774 147056
rect 204628 141500 204680 141506
rect 204628 141442 204680 141448
rect 204536 75540 204588 75546
rect 204536 75482 204588 75488
rect 204444 74180 204496 74186
rect 204444 74122 204496 74128
rect 204352 70984 204404 70990
rect 204352 70926 204404 70932
rect 204260 53780 204312 53786
rect 204260 53722 204312 53728
rect 204272 53106 204300 53722
rect 204260 53100 204312 53106
rect 204260 53042 204312 53048
rect 204166 48240 204222 48249
rect 204166 48175 204222 48184
rect 204074 47968 204130 47977
rect 204074 47903 204130 47912
rect 204088 47569 204116 47903
rect 204180 47705 204208 48175
rect 204166 47696 204222 47705
rect 204166 47631 204222 47640
rect 204260 47660 204312 47666
rect 204260 47602 204312 47608
rect 204074 47560 204130 47569
rect 204074 47495 204130 47504
rect 204272 16574 204300 47602
rect 204640 45554 204668 141442
rect 204732 46209 204760 147047
rect 204812 124908 204864 124914
rect 204812 124850 204864 124856
rect 204718 46200 204774 46209
rect 204718 46135 204774 46144
rect 204640 45526 204760 45554
rect 204732 41313 204760 45526
rect 204718 41304 204774 41313
rect 204718 41239 204774 41248
rect 204732 40633 204760 41239
rect 204718 40624 204774 40633
rect 204718 40559 204774 40568
rect 204824 35873 204852 124850
rect 204916 74089 204944 150214
rect 204996 149864 205048 149870
rect 204996 149806 205048 149812
rect 205008 80889 205036 149806
rect 205088 147008 205140 147014
rect 205088 146950 205140 146956
rect 204994 80880 205050 80889
rect 205100 80850 205128 146950
rect 204994 80815 205050 80824
rect 205088 80844 205140 80850
rect 205088 80786 205140 80792
rect 205546 75848 205602 75857
rect 205546 75783 205602 75792
rect 205560 75750 205588 75783
rect 205548 75744 205600 75750
rect 205548 75686 205600 75692
rect 204902 74080 204958 74089
rect 204902 74015 204958 74024
rect 205652 68202 205680 192782
rect 205914 192672 205970 192681
rect 205824 192636 205876 192642
rect 205914 192607 205970 192616
rect 205824 192578 205876 192584
rect 205732 190392 205784 190398
rect 205732 190334 205784 190340
rect 205640 68196 205692 68202
rect 205640 68138 205692 68144
rect 204902 67552 204958 67561
rect 204902 67487 204958 67496
rect 204916 67182 204944 67487
rect 204904 67176 204956 67182
rect 204904 67118 204956 67124
rect 204916 66298 204944 67118
rect 204904 66292 204956 66298
rect 204904 66234 204956 66240
rect 205744 66026 205772 190334
rect 205836 68542 205864 192578
rect 205928 75410 205956 192607
rect 206020 151366 206048 262686
rect 206100 260296 206152 260302
rect 206100 260238 206152 260244
rect 206008 151360 206060 151366
rect 206008 151302 206060 151308
rect 206112 151230 206140 260238
rect 207020 190052 207072 190058
rect 207020 189994 207072 190000
rect 206100 151224 206152 151230
rect 206100 151166 206152 151172
rect 206192 150204 206244 150210
rect 206192 150146 206244 150152
rect 206100 149728 206152 149734
rect 206100 149670 206152 149676
rect 206008 140140 206060 140146
rect 206008 140082 206060 140088
rect 205916 75404 205968 75410
rect 205916 75346 205968 75352
rect 205928 75206 205956 75346
rect 205916 75200 205968 75206
rect 205916 75142 205968 75148
rect 205824 68536 205876 68542
rect 205824 68478 205876 68484
rect 205732 66020 205784 66026
rect 205732 65962 205784 65968
rect 205916 45552 205968 45558
rect 205914 45520 205916 45529
rect 205968 45520 205970 45529
rect 205914 45455 205970 45464
rect 205928 44198 205956 45455
rect 205916 44192 205968 44198
rect 205916 44134 205968 44140
rect 205640 36916 205692 36922
rect 205640 36858 205692 36864
rect 204810 35864 204866 35873
rect 204810 35799 204866 35808
rect 204824 35329 204852 35799
rect 204810 35320 204866 35329
rect 204810 35255 204866 35264
rect 205652 16574 205680 36858
rect 206020 30297 206048 140082
rect 206112 74254 206140 149670
rect 206100 74248 206152 74254
rect 206100 74190 206152 74196
rect 206204 74118 206232 150146
rect 206284 150068 206336 150074
rect 206284 150010 206336 150016
rect 206296 76770 206324 150010
rect 206376 147144 206428 147150
rect 206376 147086 206428 147092
rect 206388 80753 206416 147086
rect 206468 136604 206520 136610
rect 206468 136546 206520 136552
rect 206374 80744 206430 80753
rect 206374 80679 206430 80688
rect 206284 76764 206336 76770
rect 206284 76706 206336 76712
rect 206480 75886 206508 136546
rect 206468 75880 206520 75886
rect 206282 75848 206338 75857
rect 206468 75822 206520 75828
rect 206282 75783 206338 75792
rect 206296 75682 206324 75783
rect 206376 75744 206428 75750
rect 206376 75686 206428 75692
rect 206284 75676 206336 75682
rect 206284 75618 206336 75624
rect 206296 74662 206324 75618
rect 206284 74656 206336 74662
rect 206284 74598 206336 74604
rect 206388 74594 206416 75686
rect 206376 74588 206428 74594
rect 206376 74530 206428 74536
rect 206192 74112 206244 74118
rect 206192 74054 206244 74060
rect 205730 30288 205786 30297
rect 205730 30223 205786 30232
rect 206006 30288 206062 30297
rect 206006 30223 206062 30232
rect 205744 29617 205772 30223
rect 205730 29608 205786 29617
rect 205730 29543 205786 29552
rect 207032 21865 207060 189994
rect 207124 151094 207152 277366
rect 234632 273970 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 699718 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 265624 699712 265676 699718
rect 265624 699654 265676 699660
rect 267648 699712 267700 699718
rect 267648 699654 267700 699660
rect 265636 284986 265664 699654
rect 265624 284980 265676 284986
rect 265624 284922 265676 284928
rect 234620 273964 234672 273970
rect 234620 273906 234672 273912
rect 207572 267028 207624 267034
rect 207572 266970 207624 266976
rect 207584 266490 207612 266970
rect 207572 266484 207624 266490
rect 207572 266426 207624 266432
rect 207294 200288 207350 200297
rect 207294 200223 207350 200232
rect 207204 194404 207256 194410
rect 207204 194346 207256 194352
rect 207112 151088 207164 151094
rect 207112 151030 207164 151036
rect 207110 75304 207166 75313
rect 207110 75239 207166 75248
rect 207124 75041 207152 75239
rect 207110 75032 207166 75041
rect 207110 74967 207166 74976
rect 207216 68270 207244 194346
rect 207308 75478 207336 200223
rect 207388 194200 207440 194206
rect 207388 194142 207440 194148
rect 207296 75472 207348 75478
rect 207296 75414 207348 75420
rect 207400 75177 207428 194142
rect 207480 192568 207532 192574
rect 207480 192510 207532 192516
rect 207492 75313 207520 192510
rect 207584 151162 207612 266426
rect 282932 262886 282960 702406
rect 299492 267034 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 331232 275330 331260 702986
rect 348804 699718 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 347044 699712 347096 699718
rect 347044 699654 347096 699660
rect 348792 699712 348844 699718
rect 348792 699654 348844 699660
rect 347056 290465 347084 699654
rect 347042 290456 347098 290465
rect 347042 290391 347098 290400
rect 364352 283626 364380 702406
rect 397472 699718 397500 703520
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 364340 283620 364392 283626
rect 364340 283562 364392 283568
rect 396736 282169 396764 699654
rect 396722 282160 396778 282169
rect 396722 282095 396778 282104
rect 331220 275324 331272 275330
rect 331220 275266 331272 275272
rect 299480 267028 299532 267034
rect 299480 266970 299532 266976
rect 282920 262880 282972 262886
rect 412652 262857 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 699718 429884 703520
rect 428464 699712 428516 699718
rect 428464 699654 428516 699660
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 428476 264246 428504 699654
rect 462332 660346 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 660340 462372 660346
rect 462320 660282 462372 660288
rect 477512 287706 477540 702406
rect 477500 287700 477552 287706
rect 477500 287642 477552 287648
rect 494072 271182 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 280838 527220 703520
rect 543476 700330 543504 703520
rect 559668 700330 559696 703520
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 543004 700256 543056 700262
rect 543004 700198 543056 700204
rect 527180 280832 527232 280838
rect 527180 280774 527232 280780
rect 494060 271176 494112 271182
rect 494060 271118 494112 271124
rect 543016 269822 543044 700198
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580262 365120 580318 365129
rect 580262 365055 580318 365064
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 543004 269816 543056 269822
rect 543004 269758 543056 269764
rect 428464 264240 428516 264246
rect 428464 264182 428516 264188
rect 580276 263566 580304 365055
rect 580264 263560 580316 263566
rect 580264 263502 580316 263508
rect 580540 263084 580592 263090
rect 580540 263026 580592 263032
rect 580356 263016 580408 263022
rect 580356 262958 580408 262964
rect 282920 262822 282972 262828
rect 412638 262848 412694 262857
rect 412638 262783 412694 262792
rect 472624 261316 472676 261322
rect 472624 261258 472676 261264
rect 471242 259584 471298 259593
rect 207664 259548 207716 259554
rect 471242 259519 471298 259528
rect 207664 259490 207716 259496
rect 207676 152386 207704 259490
rect 471256 206990 471284 259519
rect 472636 245614 472664 261258
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 472624 245608 472676 245614
rect 579712 245608 579764 245614
rect 472624 245550 472676 245556
rect 579710 245576 579712 245585
rect 579764 245576 579766 245585
rect 579710 245511 579766 245520
rect 471244 206984 471296 206990
rect 471244 206926 471296 206932
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 216956 200184 217008 200190
rect 209962 200152 210018 200161
rect 216956 200126 217008 200132
rect 209962 200087 210018 200096
rect 208676 194336 208728 194342
rect 208676 194278 208728 194284
rect 208490 194032 208546 194041
rect 208490 193967 208546 193976
rect 208398 190088 208454 190097
rect 208398 190023 208454 190032
rect 207940 152924 207992 152930
rect 207940 152866 207992 152872
rect 207664 152380 207716 152386
rect 207664 152322 207716 152328
rect 207572 151156 207624 151162
rect 207572 151098 207624 151104
rect 207572 150136 207624 150142
rect 207572 150078 207624 150084
rect 207478 75304 207534 75313
rect 207478 75239 207534 75248
rect 207386 75168 207442 75177
rect 207386 75103 207442 75112
rect 207584 73778 207612 150078
rect 207756 150000 207808 150006
rect 207756 149942 207808 149948
rect 207664 149932 207716 149938
rect 207664 149874 207716 149880
rect 207676 79218 207704 149874
rect 207768 81025 207796 149942
rect 207848 149796 207900 149802
rect 207848 149738 207900 149744
rect 207860 81161 207888 149738
rect 207846 81152 207902 81161
rect 207846 81087 207902 81096
rect 207754 81016 207810 81025
rect 207754 80951 207810 80960
rect 207664 79212 207716 79218
rect 207664 79154 207716 79160
rect 207664 73908 207716 73914
rect 207664 73850 207716 73856
rect 207572 73772 207624 73778
rect 207572 73714 207624 73720
rect 207204 68264 207256 68270
rect 207204 68206 207256 68212
rect 207018 21856 207074 21865
rect 207018 21791 207074 21800
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 203892 4140 203944 4146
rect 203892 4082 203944 4088
rect 203984 4140 204036 4146
rect 203984 4082 204036 4088
rect 203524 2916 203576 2922
rect 203524 2858 203576 2864
rect 203904 480 203932 4082
rect 203996 3534 204024 4082
rect 203984 3528 204036 3534
rect 203984 3470 204036 3476
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 207676 3398 207704 73850
rect 207952 72593 207980 152866
rect 207938 72584 207994 72593
rect 207938 72519 207994 72528
rect 208412 44169 208440 190023
rect 208504 51785 208532 193967
rect 208584 190324 208636 190330
rect 208584 190266 208636 190272
rect 208596 58585 208624 190266
rect 208688 69630 208716 194278
rect 208768 194132 208820 194138
rect 208768 194074 208820 194080
rect 208780 72729 208808 194074
rect 209870 191176 209926 191185
rect 209870 191111 209926 191120
rect 209778 189952 209834 189961
rect 209778 189887 209834 189896
rect 208952 187400 209004 187406
rect 208952 187342 209004 187348
rect 208860 187332 208912 187338
rect 208860 187274 208912 187280
rect 208872 77042 208900 187274
rect 208964 78946 208992 187342
rect 209136 152856 209188 152862
rect 209136 152798 209188 152804
rect 209044 152788 209096 152794
rect 209044 152730 209096 152736
rect 208952 78940 209004 78946
rect 208952 78882 209004 78888
rect 208860 77036 208912 77042
rect 208860 76978 208912 76984
rect 208766 72720 208822 72729
rect 208766 72655 208822 72664
rect 208676 69624 208728 69630
rect 208676 69566 208728 69572
rect 208582 58576 208638 58585
rect 208582 58511 208638 58520
rect 208490 51776 208546 51785
rect 208490 51711 208546 51720
rect 208492 50992 208544 50998
rect 208492 50934 208544 50940
rect 208504 50386 208532 50934
rect 208492 50380 208544 50386
rect 208492 50322 208544 50328
rect 209056 46918 209084 152730
rect 209148 50386 209176 152798
rect 209228 152652 209280 152658
rect 209228 152594 209280 152600
rect 209240 73030 209268 152594
rect 209228 73024 209280 73030
rect 209228 72966 209280 72972
rect 209136 50380 209188 50386
rect 209136 50322 209188 50328
rect 208492 46912 208544 46918
rect 208492 46854 208544 46860
rect 209044 46912 209096 46918
rect 209044 46854 209096 46860
rect 208504 46238 208532 46854
rect 208492 46232 208544 46238
rect 208492 46174 208544 46180
rect 208398 44160 208454 44169
rect 208398 44095 208454 44104
rect 208412 43489 208440 44095
rect 208398 43480 208454 43489
rect 208398 43415 208454 43424
rect 208398 30968 208454 30977
rect 208398 30903 208454 30912
rect 208412 16574 208440 30903
rect 209792 21321 209820 189887
rect 209884 33017 209912 191111
rect 209976 68882 210004 200087
rect 215392 199776 215444 199782
rect 215392 199718 215444 199724
rect 215300 199028 215352 199034
rect 215300 198970 215352 198976
rect 211436 198484 211488 198490
rect 211436 198426 211488 198432
rect 211252 198348 211304 198354
rect 211252 198290 211304 198296
rect 210332 195356 210384 195362
rect 210332 195298 210384 195304
rect 210148 194268 210200 194274
rect 210148 194210 210200 194216
rect 210056 187128 210108 187134
rect 210056 187070 210108 187076
rect 209964 68876 210016 68882
rect 209964 68818 210016 68824
rect 209964 65612 210016 65618
rect 209964 65554 210016 65560
rect 209870 33008 209926 33017
rect 209870 32943 209926 32952
rect 209778 21312 209834 21321
rect 209778 21247 209834 21256
rect 208412 16546 208624 16574
rect 207664 3392 207716 3398
rect 207664 3334 207716 3340
rect 207388 2916 207440 2922
rect 207388 2858 207440 2864
rect 207400 480 207428 2858
rect 208596 480 208624 16546
rect 209976 11694 210004 65554
rect 210068 55185 210096 187070
rect 210054 55176 210110 55185
rect 210054 55111 210110 55120
rect 210054 54496 210110 54505
rect 210054 54431 210110 54440
rect 209964 11688 210016 11694
rect 209964 11630 210016 11636
rect 210068 6914 210096 54431
rect 210160 48929 210188 194210
rect 210240 190256 210292 190262
rect 210240 190198 210292 190204
rect 210252 66230 210280 190198
rect 210344 72865 210372 195298
rect 210516 193996 210568 194002
rect 210516 193938 210568 193944
rect 210424 187468 210476 187474
rect 210424 187410 210476 187416
rect 210330 72856 210386 72865
rect 210330 72791 210386 72800
rect 210436 69494 210464 187410
rect 210528 76945 210556 193938
rect 211158 189816 211214 189825
rect 211158 189751 211214 189760
rect 210608 158636 210660 158642
rect 210608 158578 210660 158584
rect 210514 76936 210570 76945
rect 210514 76871 210570 76880
rect 210620 75070 210648 158578
rect 211066 76936 211122 76945
rect 211066 76871 211122 76880
rect 211080 76537 211108 76871
rect 211066 76528 211122 76537
rect 211066 76463 211122 76472
rect 210608 75064 210660 75070
rect 210608 75006 210660 75012
rect 210424 69488 210476 69494
rect 210424 69430 210476 69436
rect 211068 68876 211120 68882
rect 211068 68818 211120 68824
rect 211080 68338 211108 68818
rect 211068 68332 211120 68338
rect 211068 68274 211120 68280
rect 210240 66224 210292 66230
rect 210240 66166 210292 66172
rect 210146 48920 210202 48929
rect 210146 48855 210202 48864
rect 210146 44160 210202 44169
rect 210146 44095 210148 44104
rect 210200 44095 210202 44104
rect 211068 44124 211120 44130
rect 210148 44066 210200 44072
rect 211068 44066 211120 44072
rect 211080 42838 211108 44066
rect 211068 42832 211120 42838
rect 211068 42774 211120 42780
rect 211172 17921 211200 189751
rect 211264 55049 211292 198290
rect 211344 195628 211396 195634
rect 211344 195570 211396 195576
rect 211356 67318 211384 195570
rect 211448 71505 211476 198426
rect 212816 198416 212868 198422
rect 212538 198384 212594 198393
rect 212816 198358 212868 198364
rect 212538 198319 212594 198328
rect 211528 198280 211580 198286
rect 211528 198222 211580 198228
rect 211540 71738 211568 198222
rect 211804 194064 211856 194070
rect 211804 194006 211856 194012
rect 211620 191140 211672 191146
rect 211620 191082 211672 191088
rect 211528 71732 211580 71738
rect 211528 71674 211580 71680
rect 211434 71496 211490 71505
rect 211434 71431 211490 71440
rect 211632 67590 211660 191082
rect 211712 190188 211764 190194
rect 211712 190130 211764 190136
rect 211620 67584 211672 67590
rect 211620 67526 211672 67532
rect 211344 67312 211396 67318
rect 211344 67254 211396 67260
rect 211724 66162 211752 190130
rect 211816 76906 211844 194006
rect 211896 155304 211948 155310
rect 211896 155246 211948 155252
rect 211804 76900 211856 76906
rect 211804 76842 211856 76848
rect 211908 68950 211936 155246
rect 211988 142928 212040 142934
rect 211988 142870 212040 142876
rect 212000 79422 212028 142870
rect 212172 79552 212224 79558
rect 212172 79494 212224 79500
rect 212184 79422 212212 79494
rect 211988 79416 212040 79422
rect 211988 79358 212040 79364
rect 212172 79416 212224 79422
rect 212172 79358 212224 79364
rect 212448 71732 212500 71738
rect 212448 71674 212500 71680
rect 212460 71058 212488 71674
rect 212448 71052 212500 71058
rect 212448 70994 212500 71000
rect 211896 68944 211948 68950
rect 211896 68886 211948 68892
rect 211712 66156 211764 66162
rect 211712 66098 211764 66104
rect 212552 62082 212580 198319
rect 212630 193896 212686 193905
rect 212630 193831 212686 193840
rect 212540 62076 212592 62082
rect 212540 62018 212592 62024
rect 212644 60489 212672 193831
rect 212724 187536 212776 187542
rect 212724 187478 212776 187484
rect 212736 67522 212764 187478
rect 212828 79014 212856 198358
rect 213918 198248 213974 198257
rect 212908 198212 212960 198218
rect 213918 198183 213974 198192
rect 212908 198154 212960 198160
rect 212920 79490 212948 198154
rect 213000 155236 213052 155242
rect 213000 155178 213052 155184
rect 212908 79484 212960 79490
rect 212908 79426 212960 79432
rect 212816 79008 212868 79014
rect 212816 78950 212868 78956
rect 213012 70310 213040 155178
rect 213092 142860 213144 142866
rect 213092 142802 213144 142808
rect 213104 79898 213132 142802
rect 213184 141432 213236 141438
rect 213184 141374 213236 141380
rect 213196 80782 213224 141374
rect 213184 80776 213236 80782
rect 213184 80718 213236 80724
rect 213092 79892 213144 79898
rect 213092 79834 213144 79840
rect 213104 78878 213132 79834
rect 213736 79416 213788 79422
rect 213736 79358 213788 79364
rect 213748 79014 213776 79358
rect 213736 79008 213788 79014
rect 213736 78950 213788 78956
rect 213092 78872 213144 78878
rect 213092 78814 213144 78820
rect 213000 70304 213052 70310
rect 213000 70246 213052 70252
rect 212724 67516 212776 67522
rect 212724 67458 212776 67464
rect 213828 62076 213880 62082
rect 213828 62018 213880 62024
rect 213840 61402 213868 62018
rect 213828 61396 213880 61402
rect 213828 61338 213880 61344
rect 212630 60480 212686 60489
rect 212630 60415 212686 60424
rect 213826 60480 213882 60489
rect 213826 60415 213882 60424
rect 213840 59945 213868 60415
rect 213826 59936 213882 59945
rect 213826 59871 213882 59880
rect 211250 55040 211306 55049
rect 211250 54975 211306 54984
rect 211264 54505 211292 54975
rect 211250 54496 211306 54505
rect 211250 54431 211306 54440
rect 213932 40050 213960 198183
rect 214288 198144 214340 198150
rect 214010 198112 214066 198121
rect 214288 198086 214340 198092
rect 214010 198047 214066 198056
rect 214024 66065 214052 198047
rect 214194 197976 214250 197985
rect 214194 197911 214250 197920
rect 214102 186960 214158 186969
rect 214102 186895 214158 186904
rect 214010 66056 214066 66065
rect 214010 65991 214066 66000
rect 214010 62792 214066 62801
rect 214010 62727 214066 62736
rect 213920 40044 213972 40050
rect 213920 39986 213972 39992
rect 212538 28248 212594 28257
rect 212538 28183 212594 28192
rect 211158 17912 211214 17921
rect 211158 17847 211214 17856
rect 212446 17912 212502 17921
rect 212446 17847 212502 17856
rect 212460 17241 212488 17847
rect 212446 17232 212502 17241
rect 212446 17167 212502 17176
rect 212552 16574 212580 28183
rect 214024 16574 214052 62727
rect 214116 35737 214144 186895
rect 214208 58721 214236 197911
rect 214300 65521 214328 198086
rect 214472 198076 214524 198082
rect 214472 198018 214524 198024
rect 214380 193928 214432 193934
rect 214380 193870 214432 193876
rect 214286 65512 214342 65521
rect 214286 65447 214342 65456
rect 214392 64870 214420 193870
rect 214484 69737 214512 198018
rect 214656 198008 214708 198014
rect 214656 197950 214708 197956
rect 214564 195288 214616 195294
rect 214564 195230 214616 195236
rect 214470 69728 214526 69737
rect 214470 69663 214526 69672
rect 214576 69018 214604 195230
rect 214668 74534 214696 197950
rect 214748 153876 214800 153882
rect 214748 153818 214800 153824
rect 214760 78062 214788 153818
rect 214748 78056 214800 78062
rect 214748 77998 214800 78004
rect 214668 74506 214788 74534
rect 214760 71777 214788 74506
rect 214746 71768 214802 71777
rect 214746 71703 214802 71712
rect 214760 71369 214788 71703
rect 214746 71360 214802 71369
rect 214746 71295 214802 71304
rect 214564 69012 214616 69018
rect 214564 68954 214616 68960
rect 214576 68542 214604 68954
rect 214564 68536 214616 68542
rect 214564 68478 214616 68484
rect 214380 64864 214432 64870
rect 214380 64806 214432 64812
rect 214392 64190 214420 64806
rect 214380 64184 214432 64190
rect 214380 64126 214432 64132
rect 214194 58712 214250 58721
rect 214194 58647 214250 58656
rect 215312 53825 215340 198970
rect 215404 59129 215432 199718
rect 215852 199708 215904 199714
rect 215852 199650 215904 199656
rect 215484 199164 215536 199170
rect 215484 199106 215536 199112
rect 215496 63510 215524 199106
rect 215758 195392 215814 195401
rect 215758 195327 215814 195336
rect 215668 187264 215720 187270
rect 215668 187206 215720 187212
rect 215574 155272 215630 155281
rect 215574 155207 215630 155216
rect 215484 63504 215536 63510
rect 215484 63446 215536 63452
rect 215496 62898 215524 63446
rect 215484 62892 215536 62898
rect 215484 62834 215536 62840
rect 215390 59120 215446 59129
rect 215390 59055 215446 59064
rect 215298 53816 215354 53825
rect 215298 53751 215354 53760
rect 215312 53417 215340 53751
rect 215298 53408 215354 53417
rect 215298 53343 215354 53352
rect 215300 47592 215352 47598
rect 215300 47534 215352 47540
rect 214380 40044 214432 40050
rect 214380 39986 214432 39992
rect 214392 39506 214420 39986
rect 214380 39500 214432 39506
rect 214380 39442 214432 39448
rect 214102 35728 214158 35737
rect 214102 35663 214158 35672
rect 214116 35193 214144 35663
rect 214102 35184 214158 35193
rect 214102 35119 214158 35128
rect 212552 16546 213408 16574
rect 214024 16546 214512 16574
rect 210976 11688 211028 11694
rect 210976 11630 211028 11636
rect 209792 6886 210096 6914
rect 209792 480 209820 6886
rect 210988 480 211016 11630
rect 212172 4072 212224 4078
rect 212172 4014 212224 4020
rect 212184 480 212212 4014
rect 213380 480 213408 16546
rect 214484 480 214512 16546
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 47534
rect 215588 33153 215616 155207
rect 215680 66201 215708 187206
rect 215772 74225 215800 195327
rect 215864 81122 215892 199650
rect 215944 199096 215996 199102
rect 215944 199038 215996 199044
rect 215852 81116 215904 81122
rect 215852 81058 215904 81064
rect 215956 81002 215984 199038
rect 216678 192536 216734 192545
rect 216678 192471 216734 192480
rect 216864 192500 216916 192506
rect 216036 158432 216088 158438
rect 216036 158374 216088 158380
rect 215864 80974 215984 81002
rect 215864 80102 215892 80974
rect 215852 80096 215904 80102
rect 215852 80038 215904 80044
rect 215864 78606 215892 80038
rect 216048 79626 216076 158374
rect 216128 81116 216180 81122
rect 216128 81058 216180 81064
rect 216036 79620 216088 79626
rect 216036 79562 216088 79568
rect 215852 78600 215904 78606
rect 215852 78542 215904 78548
rect 216140 78062 216168 81058
rect 215852 78056 215904 78062
rect 215852 77998 215904 78004
rect 216128 78056 216180 78062
rect 216128 77998 216180 78004
rect 215864 77654 215892 77998
rect 215852 77648 215904 77654
rect 215852 77590 215904 77596
rect 215758 74216 215814 74225
rect 215758 74151 215814 74160
rect 215666 66192 215722 66201
rect 215666 66127 215722 66136
rect 215574 33144 215630 33153
rect 215574 33079 215630 33088
rect 215588 32473 215616 33079
rect 215574 32464 215630 32473
rect 215574 32399 215630 32408
rect 216692 22001 216720 192471
rect 216864 192442 216916 192448
rect 216772 79824 216824 79830
rect 216772 79766 216824 79772
rect 216784 78810 216812 79766
rect 216772 78804 216824 78810
rect 216772 78746 216824 78752
rect 216772 75336 216824 75342
rect 216772 75278 216824 75284
rect 216678 21992 216734 22001
rect 216678 21927 216734 21936
rect 216784 16574 216812 75278
rect 216876 38593 216904 192442
rect 216968 50969 216996 200126
rect 217600 199640 217652 199646
rect 217600 199582 217652 199588
rect 217048 199572 217100 199578
rect 217048 199514 217100 199520
rect 217060 59265 217088 199514
rect 217322 198792 217378 198801
rect 217322 198727 217378 198736
rect 217138 195664 217194 195673
rect 217138 195599 217194 195608
rect 217046 59256 217102 59265
rect 217046 59191 217102 59200
rect 217152 59106 217180 195599
rect 217230 195528 217286 195537
rect 217230 195463 217286 195472
rect 217060 59078 217180 59106
rect 217060 56574 217088 59078
rect 217244 57905 217272 195463
rect 217336 63345 217364 198727
rect 217416 186992 217468 186998
rect 217416 186934 217468 186940
rect 217428 79830 217456 186934
rect 217508 158364 217560 158370
rect 217508 158306 217560 158312
rect 217416 79824 217468 79830
rect 217416 79766 217468 79772
rect 217520 79694 217548 158306
rect 217508 79688 217560 79694
rect 217508 79630 217560 79636
rect 217612 63481 217640 199582
rect 219532 199232 219584 199238
rect 219532 199174 219584 199180
rect 218150 196616 218206 196625
rect 218150 196551 218206 196560
rect 218060 158024 218112 158030
rect 218060 157966 218112 157972
rect 218072 77330 218100 157966
rect 217980 77302 218100 77330
rect 217980 76945 218008 77302
rect 218060 77240 218112 77246
rect 218060 77182 218112 77188
rect 217966 76936 218022 76945
rect 217966 76871 218022 76880
rect 218072 76702 218100 77182
rect 218060 76696 218112 76702
rect 218060 76638 218112 76644
rect 218164 74361 218192 196551
rect 219438 191040 219494 191049
rect 219438 190975 219494 190984
rect 218244 187060 218296 187066
rect 218244 187002 218296 187008
rect 218256 74458 218284 187002
rect 218428 152992 218480 152998
rect 218428 152934 218480 152940
rect 218336 152584 218388 152590
rect 218336 152526 218388 152532
rect 218348 77246 218376 152526
rect 218336 77240 218388 77246
rect 218336 77182 218388 77188
rect 218440 77178 218468 152934
rect 218518 152552 218574 152561
rect 218518 152487 218574 152496
rect 218612 152516 218664 152522
rect 218428 77172 218480 77178
rect 218428 77114 218480 77120
rect 218334 77072 218390 77081
rect 218334 77007 218390 77016
rect 218348 76673 218376 77007
rect 218440 76770 218468 77114
rect 218532 77081 218560 152487
rect 218612 152458 218664 152464
rect 218518 77072 218574 77081
rect 218518 77007 218574 77016
rect 218518 76936 218574 76945
rect 218518 76871 218574 76880
rect 218428 76764 218480 76770
rect 218428 76706 218480 76712
rect 218334 76664 218390 76673
rect 218334 76599 218390 76608
rect 218532 76401 218560 76871
rect 218624 76702 218652 152458
rect 218702 78840 218758 78849
rect 218702 78775 218758 78784
rect 218612 76696 218664 76702
rect 218612 76638 218664 76644
rect 218518 76392 218574 76401
rect 218518 76327 218574 76336
rect 218244 74452 218296 74458
rect 218244 74394 218296 74400
rect 218150 74352 218206 74361
rect 218150 74287 218206 74296
rect 218164 73953 218192 74287
rect 218150 73944 218206 73953
rect 218256 73914 218284 74394
rect 218150 73879 218206 73888
rect 218244 73908 218296 73914
rect 218244 73850 218296 73856
rect 217598 63472 217654 63481
rect 217598 63407 217654 63416
rect 217322 63336 217378 63345
rect 217322 63271 217378 63280
rect 217336 62801 217364 63271
rect 217322 62792 217378 62801
rect 217322 62727 217378 62736
rect 217230 57896 217286 57905
rect 217230 57831 217286 57840
rect 217244 57225 217272 57831
rect 217230 57216 217286 57225
rect 217230 57151 217286 57160
rect 217048 56568 217100 56574
rect 217048 56510 217100 56516
rect 217060 55894 217088 56510
rect 217048 55888 217100 55894
rect 217048 55830 217100 55836
rect 217324 51740 217376 51746
rect 217324 51682 217376 51688
rect 216954 50960 217010 50969
rect 216954 50895 217010 50904
rect 216862 38584 216918 38593
rect 216862 38519 216918 38528
rect 217046 38584 217102 38593
rect 217046 38519 217102 38528
rect 217060 37913 217088 38519
rect 217046 37904 217102 37913
rect 217046 37839 217102 37848
rect 216784 16546 216904 16574
rect 216876 480 216904 16546
rect 217336 3126 217364 51682
rect 218716 16574 218744 78775
rect 218888 77104 218940 77110
rect 218888 77046 218940 77052
rect 218900 76634 218928 77046
rect 218888 76628 218940 76634
rect 218888 76570 218940 76576
rect 219452 46753 219480 190975
rect 219544 60353 219572 199174
rect 220820 196648 220872 196654
rect 220820 196590 220872 196596
rect 219624 189984 219676 189990
rect 219624 189926 219676 189932
rect 219636 73001 219664 189926
rect 219716 187196 219768 187202
rect 219716 187138 219768 187144
rect 219728 74050 219756 187138
rect 219900 158228 219952 158234
rect 219900 158170 219952 158176
rect 219808 158092 219860 158098
rect 219808 158034 219860 158040
rect 219716 74044 219768 74050
rect 219716 73986 219768 73992
rect 219622 72992 219678 73001
rect 219622 72927 219678 72936
rect 219820 70854 219848 158034
rect 219912 75138 219940 158170
rect 219992 158160 220044 158166
rect 219992 158102 220044 158108
rect 220004 79762 220032 158102
rect 219992 79756 220044 79762
rect 219992 79698 220044 79704
rect 219900 75132 219952 75138
rect 219900 75074 219952 75080
rect 220832 74526 220860 196590
rect 220910 195256 220966 195265
rect 220910 195191 220966 195200
rect 220820 74520 220872 74526
rect 220820 74462 220872 74468
rect 220832 74050 220860 74462
rect 220820 74044 220872 74050
rect 220820 73986 220872 73992
rect 219808 70848 219860 70854
rect 219808 70790 219860 70796
rect 220820 68604 220872 68610
rect 220820 68546 220872 68552
rect 219530 60344 219586 60353
rect 219530 60279 219586 60288
rect 220084 56228 220136 56234
rect 220084 56170 220136 56176
rect 219438 46744 219494 46753
rect 219438 46679 219494 46688
rect 219440 17468 219492 17474
rect 219440 17410 219492 17416
rect 219452 16574 219480 17410
rect 218716 16546 219296 16574
rect 219452 16546 220032 16574
rect 217324 3120 217376 3126
rect 217324 3062 217376 3068
rect 218060 3120 218112 3126
rect 218060 3062 218112 3068
rect 218072 480 218100 3062
rect 219268 480 219296 16546
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220096 3194 220124 56170
rect 220832 16574 220860 68546
rect 220924 46889 220952 195191
rect 221372 193860 221424 193866
rect 221372 193802 221424 193808
rect 221096 189916 221148 189922
rect 221096 189858 221148 189864
rect 221004 189848 221056 189854
rect 221004 189790 221056 189796
rect 221016 73137 221044 189790
rect 221002 73128 221058 73137
rect 221108 73098 221136 189858
rect 221188 189780 221240 189786
rect 221188 189722 221240 189728
rect 221200 79286 221228 189722
rect 221278 189680 221334 189689
rect 221278 189615 221334 189624
rect 221188 79280 221240 79286
rect 221188 79222 221240 79228
rect 221292 73681 221320 189615
rect 221384 93854 221412 193802
rect 580368 192545 580396 262958
rect 580448 262404 580500 262410
rect 580448 262346 580500 262352
rect 580460 219065 580488 262346
rect 580552 232393 580580 263026
rect 580538 232384 580594 232393
rect 580538 232319 580594 232328
rect 580446 219056 580502 219065
rect 580446 218991 580502 219000
rect 580354 192536 580410 192545
rect 580354 192471 580410 192480
rect 580354 179208 580410 179217
rect 580354 179143 580410 179152
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 580078 152688 580134 152697
rect 580078 152623 580134 152632
rect 580092 151842 580120 152623
rect 580080 151836 580132 151842
rect 580080 151778 580132 151784
rect 580262 150512 580318 150521
rect 580262 150447 580318 150456
rect 549904 142316 549956 142322
rect 549904 142258 549956 142264
rect 482282 141128 482338 141137
rect 482282 141063 482338 141072
rect 327724 139460 327776 139466
rect 327724 139402 327776 139408
rect 221384 93826 221504 93854
rect 221372 79280 221424 79286
rect 221372 79222 221424 79228
rect 221278 73672 221334 73681
rect 221278 73607 221334 73616
rect 221292 73273 221320 73607
rect 221278 73264 221334 73273
rect 221278 73199 221334 73208
rect 221002 73063 221058 73072
rect 221096 73092 221148 73098
rect 221096 73034 221148 73040
rect 221384 72826 221412 79222
rect 221476 78033 221504 93826
rect 302240 80776 302292 80782
rect 302240 80718 302292 80724
rect 288440 80096 288492 80102
rect 288440 80038 288492 80044
rect 238760 79892 238812 79898
rect 238760 79834 238812 79840
rect 234618 78704 234674 78713
rect 234618 78639 234674 78648
rect 221462 78024 221518 78033
rect 221462 77959 221518 77968
rect 222106 78024 222162 78033
rect 222106 77959 222162 77968
rect 222120 77353 222148 77959
rect 222106 77344 222162 77353
rect 222106 77279 222162 77288
rect 224222 73264 224278 73273
rect 224222 73199 224278 73208
rect 222108 73092 222160 73098
rect 222108 73034 222160 73040
rect 221372 72820 221424 72826
rect 221372 72762 221424 72768
rect 221384 72282 221412 72762
rect 222120 72690 222148 73034
rect 222108 72684 222160 72690
rect 222108 72626 222160 72632
rect 221372 72276 221424 72282
rect 221372 72218 221424 72224
rect 220910 46880 220966 46889
rect 220910 46815 220966 46824
rect 220832 16546 221136 16574
rect 220084 3188 220136 3194
rect 220084 3130 220136 3136
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 224236 4078 224264 73199
rect 227718 66872 227774 66881
rect 227718 66807 227774 66816
rect 224960 64456 225012 64462
rect 224960 64398 225012 64404
rect 224972 16574 225000 64398
rect 225604 32564 225656 32570
rect 225604 32506 225656 32512
rect 224972 16546 225184 16574
rect 224224 4072 224276 4078
rect 224224 4014 224276 4020
rect 223948 3392 224000 3398
rect 223948 3334 224000 3340
rect 222752 3188 222804 3194
rect 222752 3130 222804 3136
rect 222764 480 222792 3130
rect 223960 480 223988 3334
rect 225156 480 225184 16546
rect 225616 3398 225644 32506
rect 227732 16574 227760 66807
rect 230478 61704 230534 61713
rect 230478 61639 230534 61648
rect 229098 40760 229154 40769
rect 229098 40695 229154 40704
rect 229112 16574 229140 40695
rect 230492 16574 230520 61639
rect 233240 46300 233292 46306
rect 233240 46242 233292 46248
rect 231858 45248 231914 45257
rect 231858 45183 231914 45192
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 227536 16176 227588 16182
rect 227536 16118 227588 16124
rect 225604 3392 225656 3398
rect 225604 3334 225656 3340
rect 226340 3392 226392 3398
rect 226340 3334 226392 3340
rect 226352 480 226380 3334
rect 227548 480 227576 16118
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 45183
rect 233252 16574 233280 46242
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 11694 234660 78639
rect 237378 74080 237434 74089
rect 237378 74015 237434 74024
rect 236000 39636 236052 39642
rect 236000 39578 236052 39584
rect 236012 16574 236040 39578
rect 237392 16574 237420 74015
rect 238772 16574 238800 79834
rect 252560 79824 252612 79830
rect 252560 79766 252612 79772
rect 247682 76936 247738 76945
rect 247682 76871 247738 76880
rect 245658 63200 245714 63209
rect 245658 63135 245714 63144
rect 242900 53236 242952 53242
rect 242900 53178 242952 53184
rect 239404 42356 239456 42362
rect 239404 42298 239456 42304
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 238772 16546 239352 16574
rect 234620 11688 234672 11694
rect 234620 11630 234672 11636
rect 235816 11688 235868 11694
rect 235816 11630 235868 11636
rect 234620 10600 234672 10606
rect 234620 10542 234672 10548
rect 234632 480 234660 10542
rect 235828 480 235856 11630
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239324 480 239352 16546
rect 239416 3398 239444 42298
rect 241704 12028 241756 12034
rect 241704 11970 241756 11976
rect 239404 3392 239456 3398
rect 239404 3334 239456 3340
rect 240508 3392 240560 3398
rect 240508 3334 240560 3340
rect 240520 480 240548 3334
rect 241716 480 241744 11970
rect 242912 480 242940 53178
rect 242992 32496 243044 32502
rect 242992 32438 243044 32444
rect 243004 16574 243032 32438
rect 245672 16574 245700 63135
rect 243004 16546 244136 16574
rect 245672 16546 245976 16574
rect 244108 480 244136 16546
rect 245200 5092 245252 5098
rect 245200 5034 245252 5040
rect 245212 480 245240 5034
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247696 4146 247724 76871
rect 248420 73840 248472 73846
rect 248420 73782 248472 73788
rect 247592 4140 247644 4146
rect 247592 4082 247644 4088
rect 247684 4140 247736 4146
rect 247684 4082 247736 4088
rect 247604 480 247632 4082
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 73782
rect 251180 61600 251232 61606
rect 251180 61542 251232 61548
rect 249798 58984 249854 58993
rect 249798 58919 249854 58928
rect 249812 16574 249840 58919
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 480 251220 61542
rect 252572 16574 252600 79766
rect 268382 78160 268438 78169
rect 268382 78095 268438 78104
rect 260838 76800 260894 76809
rect 260838 76735 260894 76744
rect 255318 73944 255374 73953
rect 255318 73879 255374 73888
rect 255332 16574 255360 73879
rect 256700 64388 256752 64394
rect 256700 64330 256752 64336
rect 252572 16546 253520 16574
rect 255332 16546 255912 16574
rect 252376 6588 252428 6594
rect 252376 6530 252428 6536
rect 252388 480 252416 6530
rect 253492 480 253520 16546
rect 254676 4140 254728 4146
rect 254676 4082 254728 4088
rect 254688 480 254716 4082
rect 255884 480 255912 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 354 256740 64330
rect 259460 60172 259512 60178
rect 259460 60114 259512 60120
rect 257344 38140 257396 38146
rect 257344 38082 257396 38088
rect 257356 4146 257384 38082
rect 259472 11694 259500 60114
rect 259550 46472 259606 46481
rect 259550 46407 259606 46416
rect 259460 11688 259512 11694
rect 259460 11630 259512 11636
rect 259564 6914 259592 46407
rect 260852 16574 260880 76735
rect 268396 73846 268424 78095
rect 270500 78056 270552 78062
rect 270500 77998 270552 78004
rect 269120 74044 269172 74050
rect 269120 73986 269172 73992
rect 268384 73840 268436 73846
rect 261482 73808 261538 73817
rect 268384 73782 268436 73788
rect 261482 73743 261538 73752
rect 260852 16546 261432 16574
rect 260656 11688 260708 11694
rect 260656 11630 260708 11636
rect 259472 6886 259592 6914
rect 257344 4140 257396 4146
rect 257344 4082 257396 4088
rect 258264 4140 258316 4146
rect 258264 4082 258316 4088
rect 258276 480 258304 4082
rect 259472 480 259500 6886
rect 260668 480 260696 11630
rect 261404 3482 261432 16546
rect 261496 4146 261524 73743
rect 263600 57452 263652 57458
rect 263600 57394 263652 57400
rect 263612 16574 263640 57394
rect 267740 43580 267792 43586
rect 267740 43522 267792 43528
rect 264980 31204 265032 31210
rect 264980 31146 265032 31152
rect 263612 16546 264192 16574
rect 261484 4140 261536 4146
rect 261484 4082 261536 4088
rect 262956 4140 263008 4146
rect 262956 4082 263008 4088
rect 261404 3454 261800 3482
rect 261772 480 261800 3454
rect 262968 480 262996 4082
rect 264164 480 264192 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 31146
rect 266358 18592 266414 18601
rect 266358 18527 266414 18536
rect 266372 16574 266400 18527
rect 266372 16546 266584 16574
rect 266556 480 266584 16546
rect 267752 480 267780 43522
rect 267832 36848 267884 36854
rect 267832 36790 267884 36796
rect 267844 16574 267872 36790
rect 269132 16574 269160 73986
rect 270512 16574 270540 77998
rect 287704 77376 287756 77382
rect 287704 77318 287756 77324
rect 283564 72752 283616 72758
rect 283564 72694 283616 72700
rect 274640 67040 274692 67046
rect 274640 66982 274692 66988
rect 273260 18828 273312 18834
rect 273260 18770 273312 18776
rect 267844 16546 268424 16574
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 270052 480 270080 16546
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272432 13388 272484 13394
rect 272432 13330 272484 13336
rect 272444 480 272472 13330
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 18770
rect 274652 16574 274680 66982
rect 277400 61532 277452 61538
rect 277400 61474 277452 61480
rect 276110 39264 276166 39273
rect 276110 39199 276166 39208
rect 275284 27192 275336 27198
rect 275284 27134 275336 27140
rect 274652 16546 274864 16574
rect 274836 480 274864 16546
rect 275296 3398 275324 27134
rect 276124 16574 276152 39199
rect 277412 16574 277440 61474
rect 281538 58848 281594 58857
rect 281538 58783 281594 58792
rect 278780 25832 278832 25838
rect 278780 25774 278832 25780
rect 278792 16574 278820 25774
rect 280160 20188 280212 20194
rect 280160 20130 280212 20136
rect 280172 16574 280200 20130
rect 276124 16546 276704 16574
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 275284 3392 275336 3398
rect 275284 3334 275336 3340
rect 276020 3392 276072 3398
rect 276020 3334 276072 3340
rect 276032 480 276060 3334
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 16546
rect 278332 480 278360 16546
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 58783
rect 282920 24336 282972 24342
rect 282920 24278 282972 24284
rect 282932 16574 282960 24278
rect 282932 16546 283144 16574
rect 283116 480 283144 16546
rect 283576 4146 283604 72694
rect 284390 53408 284446 53417
rect 284390 53343 284446 53352
rect 284404 16574 284432 53343
rect 285680 49020 285732 49026
rect 285680 48962 285732 48968
rect 285692 16574 285720 48962
rect 287716 20058 287744 77318
rect 287060 20052 287112 20058
rect 287060 19994 287112 20000
rect 287704 20052 287756 20058
rect 287704 19994 287756 20000
rect 287072 16574 287100 19994
rect 288452 16574 288480 80038
rect 289820 76764 289872 76770
rect 289820 76706 289872 76712
rect 284404 16546 284984 16574
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 288452 16546 289032 16574
rect 283564 4140 283616 4146
rect 283564 4082 283616 4088
rect 284300 4072 284352 4078
rect 284300 4014 284352 4020
rect 284312 480 284340 4014
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 354 284984 16546
rect 286612 480 286640 16546
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 289004 480 289032 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 76706
rect 296720 76696 296772 76702
rect 296720 76638 296772 76644
rect 295338 65784 295394 65793
rect 295338 65719 295394 65728
rect 292580 62892 292632 62898
rect 292580 62834 292632 62840
rect 291200 20120 291252 20126
rect 291200 20062 291252 20068
rect 291212 16574 291240 20062
rect 291212 16546 291424 16574
rect 291396 480 291424 16546
rect 292592 480 292620 62834
rect 293958 37904 294014 37913
rect 293958 37839 294014 37848
rect 293972 16574 294000 37839
rect 295352 16574 295380 65719
rect 296732 16574 296760 76638
rect 299480 60104 299532 60110
rect 299480 60046 299532 60052
rect 293972 16546 294920 16574
rect 295352 16546 295656 16574
rect 296732 16546 297312 16574
rect 293224 14748 293276 14754
rect 293224 14690 293276 14696
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 14690
rect 294892 480 294920 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 297284 480 297312 16546
rect 298468 4140 298520 4146
rect 298468 4082 298520 4088
rect 298480 480 298508 4082
rect 299492 3482 299520 60046
rect 299572 29844 299624 29850
rect 299572 29786 299624 29792
rect 299584 4078 299612 29786
rect 302252 16574 302280 80718
rect 306380 77988 306432 77994
rect 306380 77930 306432 77936
rect 305000 72616 305052 72622
rect 305000 72558 305052 72564
rect 303618 35320 303674 35329
rect 303618 35255 303674 35264
rect 303632 16574 303660 35255
rect 305012 16574 305040 72558
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 301964 9172 302016 9178
rect 301964 9114 302016 9120
rect 299572 4072 299624 4078
rect 299572 4014 299624 4020
rect 300768 4072 300820 4078
rect 300768 4014 300820 4020
rect 299492 3454 299704 3482
rect 299676 480 299704 3454
rect 300780 480 300808 4014
rect 301976 480 302004 9114
rect 303172 480 303200 16546
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 77930
rect 322940 73976 322992 73982
rect 322940 73918 322992 73924
rect 311164 72820 311216 72826
rect 311164 72762 311216 72768
rect 309140 57384 309192 57390
rect 309140 57326 309192 57332
rect 307024 40928 307076 40934
rect 307024 40870 307076 40876
rect 307036 3398 307064 40870
rect 309152 16574 309180 57326
rect 310520 23044 310572 23050
rect 310520 22986 310572 22992
rect 310532 16574 310560 22986
rect 309152 16546 309824 16574
rect 310532 16546 311112 16574
rect 307944 13320 307996 13326
rect 307944 13262 307996 13268
rect 307024 3392 307076 3398
rect 307024 3334 307076 3340
rect 307956 480 307984 13262
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311084 3482 311112 16546
rect 311176 4078 311204 72762
rect 318798 72584 318854 72593
rect 318798 72519 318854 72528
rect 317420 69828 317472 69834
rect 317420 69770 317472 69776
rect 313280 56160 313332 56166
rect 313280 56102 313332 56108
rect 313292 16574 313320 56102
rect 315302 54768 315358 54777
rect 315302 54703 315358 54712
rect 313292 16546 313872 16574
rect 311164 4072 311216 4078
rect 311164 4014 311216 4020
rect 312636 4072 312688 4078
rect 312636 4014 312688 4020
rect 311084 3454 311480 3482
rect 311452 480 311480 3454
rect 312648 480 312676 4014
rect 313844 480 313872 16546
rect 314660 14680 314712 14686
rect 314660 14622 314712 14628
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 354 314700 14622
rect 315316 3194 315344 54703
rect 316130 17232 316186 17241
rect 316130 17167 316186 17176
rect 316144 16574 316172 17167
rect 317432 16574 317460 69770
rect 318812 16574 318840 72519
rect 320180 51128 320232 51134
rect 320180 51070 320232 51076
rect 320192 16574 320220 51070
rect 321560 28484 321612 28490
rect 321560 28426 321612 28432
rect 321572 16574 321600 28426
rect 316144 16546 316264 16574
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 315304 3188 315356 3194
rect 315304 3130 315356 3136
rect 316236 480 316264 16546
rect 317328 3188 317380 3194
rect 317328 3130 317380 3136
rect 317340 480 317368 3130
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 73918
rect 327736 73166 327764 139402
rect 482296 86970 482324 141063
rect 549916 100706 549944 142258
rect 579804 142248 579856 142254
rect 579804 142190 579856 142196
rect 579816 139369 579844 142190
rect 579802 139360 579858 139369
rect 579802 139295 579858 139304
rect 549904 100700 549956 100706
rect 549904 100642 549956 100648
rect 579620 100700 579672 100706
rect 579620 100642 579672 100648
rect 579632 99521 579660 100642
rect 579618 99512 579674 99521
rect 579618 99447 579674 99456
rect 482284 86964 482336 86970
rect 482284 86906 482336 86912
rect 579620 86964 579672 86970
rect 579620 86906 579672 86912
rect 579632 86193 579660 86906
rect 579618 86184 579674 86193
rect 579618 86119 579674 86128
rect 380900 80708 380952 80714
rect 380900 80650 380952 80656
rect 376760 79620 376812 79626
rect 376760 79562 376812 79568
rect 342902 78024 342958 78033
rect 342902 77959 342958 77968
rect 327724 73160 327776 73166
rect 327724 73102 327776 73108
rect 324964 72684 325016 72690
rect 324964 72626 325016 72632
rect 324318 40624 324374 40633
rect 324318 40559 324374 40568
rect 324332 16574 324360 40559
rect 324332 16546 324452 16574
rect 324424 480 324452 16546
rect 324976 3058 325004 72626
rect 340880 72548 340932 72554
rect 340880 72490 340932 72496
rect 332598 72448 332654 72457
rect 332598 72383 332654 72392
rect 331220 62824 331272 62830
rect 331220 62766 331272 62772
rect 327080 58744 327132 58750
rect 327080 58686 327132 58692
rect 327092 16574 327120 58686
rect 329104 21412 329156 21418
rect 329104 21354 329156 21360
rect 327092 16546 328040 16574
rect 325608 9104 325660 9110
rect 325608 9046 325660 9052
rect 324964 3052 325016 3058
rect 324964 2994 325016 3000
rect 325620 480 325648 9046
rect 326804 3052 326856 3058
rect 326804 2994 326856 3000
rect 326816 480 326844 2994
rect 328012 480 328040 16546
rect 328736 11960 328788 11966
rect 328736 11902 328788 11908
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 354 328776 11902
rect 329116 3398 329144 21354
rect 329104 3392 329156 3398
rect 329104 3334 329156 3340
rect 330392 3392 330444 3398
rect 330392 3334 330444 3340
rect 330404 480 330432 3334
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 62766
rect 332612 3398 332640 72383
rect 332692 66972 332744 66978
rect 332692 66914 332744 66920
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 66914
rect 338120 50448 338172 50454
rect 338120 50390 338172 50396
rect 333978 29608 334034 29617
rect 333978 29543 334034 29552
rect 333992 16574 334020 29543
rect 336738 21584 336794 21593
rect 336738 21519 336794 21528
rect 336752 16574 336780 21519
rect 338132 16574 338160 50390
rect 339500 32428 339552 32434
rect 339500 32370 339552 32376
rect 333992 16546 334664 16574
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336280 10532 336332 10538
rect 336280 10474 336332 10480
rect 336292 480 336320 10474
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 32370
rect 340892 3210 340920 72490
rect 340972 64320 341024 64326
rect 340972 64262 341024 64268
rect 340984 3398 341012 64262
rect 342916 21418 342944 77959
rect 367098 76664 367154 76673
rect 353300 76628 353352 76634
rect 367098 76599 367154 76608
rect 353300 76570 353352 76576
rect 345020 69760 345072 69766
rect 345020 69702 345072 69708
rect 342994 21448 343050 21457
rect 342904 21412 342956 21418
rect 342994 21383 343050 21392
rect 342904 21354 342956 21360
rect 340972 3392 341024 3398
rect 340972 3334 341024 3340
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 340892 3182 341012 3210
rect 340984 480 341012 3182
rect 342180 480 342208 3334
rect 343008 3262 343036 21383
rect 345032 16574 345060 69702
rect 349160 60036 349212 60042
rect 349160 59978 349212 59984
rect 346400 34060 346452 34066
rect 346400 34002 346452 34008
rect 346412 16574 346440 34002
rect 347778 21312 347834 21321
rect 347778 21247 347834 21256
rect 347792 16574 347820 21247
rect 349172 16574 349200 59978
rect 351920 56092 351972 56098
rect 351920 56034 351972 56040
rect 350540 42288 350592 42294
rect 350540 42230 350592 42236
rect 350552 16574 350580 42230
rect 351932 16574 351960 56034
rect 353312 16574 353340 76570
rect 354680 73908 354732 73914
rect 354680 73850 354732 73856
rect 354692 16574 354720 73850
rect 358820 68536 358872 68542
rect 358820 68478 358872 68484
rect 356058 49328 356114 49337
rect 356058 49263 356114 49272
rect 356072 16574 356100 49263
rect 357440 31136 357492 31142
rect 357440 31078 357492 31084
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 349172 16546 349292 16574
rect 350552 16546 351224 16574
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 356072 16546 356376 16574
rect 343364 7880 343416 7886
rect 343364 7822 343416 7828
rect 342996 3256 343048 3262
rect 342996 3198 343048 3204
rect 343376 480 343404 7822
rect 344560 3256 344612 3262
rect 344560 3198 344612 3204
rect 344572 480 344600 3198
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349264 480 349292 16546
rect 350448 6520 350500 6526
rect 350448 6462 350500 6468
rect 350460 480 350488 6462
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352852 480 352880 16546
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356348 480 356376 16546
rect 357452 3210 357480 31078
rect 357532 19984 357584 19990
rect 357532 19926 357584 19932
rect 357544 3398 357572 19926
rect 358832 16574 358860 68478
rect 362960 57316 363012 57322
rect 362960 57258 363012 57264
rect 361580 36780 361632 36786
rect 361580 36722 361632 36728
rect 361592 16574 361620 36722
rect 362972 16574 363000 57258
rect 364982 54632 365038 54641
rect 364982 54567 365038 54576
rect 358832 16546 359504 16574
rect 361592 16546 361896 16574
rect 362972 16546 363552 16574
rect 357532 3392 357584 3398
rect 357532 3334 357584 3340
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 357452 3182 357572 3210
rect 357544 480 357572 3182
rect 358740 480 358768 3334
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 361120 16108 361172 16114
rect 361120 16050 361172 16056
rect 361132 480 361160 16050
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363524 480 363552 16546
rect 364616 16040 364668 16046
rect 364616 15982 364668 15988
rect 364628 480 364656 15982
rect 364996 3398 365024 54567
rect 367112 16574 367140 76599
rect 368480 69692 368532 69698
rect 368480 69634 368532 69640
rect 368492 16574 368520 69634
rect 375380 66904 375432 66910
rect 375380 66846 375432 66852
rect 369858 52184 369914 52193
rect 369858 52119 369914 52128
rect 369872 16574 369900 52119
rect 373998 50552 374054 50561
rect 373998 50487 374054 50496
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 369872 16546 370176 16574
rect 365812 7812 365864 7818
rect 365812 7754 365864 7760
rect 364984 3392 365036 3398
rect 364984 3334 365036 3340
rect 365824 480 365852 7754
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367020 480 367048 3334
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 372896 10464 372948 10470
rect 372896 10406 372948 10412
rect 371700 5024 371752 5030
rect 371700 4966 371752 4972
rect 371712 480 371740 4966
rect 372908 480 372936 10406
rect 374012 1170 374040 50487
rect 374092 27124 374144 27130
rect 374092 27066 374144 27072
rect 374104 3398 374132 27066
rect 375392 16574 375420 66846
rect 376772 16574 376800 79562
rect 378140 25764 378192 25770
rect 378140 25706 378192 25712
rect 378152 16574 378180 25706
rect 380912 16574 380940 80650
rect 480260 79552 480312 79558
rect 480260 79494 480312 79500
rect 453304 77308 453356 77314
rect 453304 77250 453356 77256
rect 389180 76560 389232 76566
rect 389180 76502 389232 76508
rect 382280 72480 382332 72486
rect 382280 72422 382332 72428
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 378152 16546 378456 16574
rect 380912 16546 381216 16574
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374012 1142 374132 1170
rect 374104 480 374132 1142
rect 375300 480 375328 3334
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 370566 -960 370678 326
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 379520 11892 379572 11898
rect 379520 11834 379572 11840
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 11834
rect 381188 480 381216 16546
rect 382292 1018 382320 72422
rect 382922 53272 382978 53281
rect 382922 53207 382978 53216
rect 382372 13252 382424 13258
rect 382372 13194 382424 13200
rect 382280 1012 382332 1018
rect 382280 954 382332 960
rect 382384 480 382412 13194
rect 382936 3058 382964 53207
rect 387798 49192 387854 49201
rect 387798 49127 387854 49136
rect 385960 14612 386012 14618
rect 385960 14554 386012 14560
rect 382924 3052 382976 3058
rect 382924 2994 382976 3000
rect 384764 3052 384816 3058
rect 384764 2994 384816 3000
rect 383568 1012 383620 1018
rect 383568 954 383620 960
rect 383580 480 383608 954
rect 384776 480 384804 2994
rect 385972 480 386000 14554
rect 386696 13184 386748 13190
rect 386696 13126 386748 13132
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386708 354 386736 13126
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 49127
rect 389192 16574 389220 76502
rect 396080 68468 396132 68474
rect 396080 68410 396132 68416
rect 394700 61464 394752 61470
rect 394700 61406 394752 61412
rect 390558 45112 390614 45121
rect 390558 45047 390614 45056
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 3398 390600 45047
rect 390650 32600 390706 32609
rect 390650 32535 390706 32544
rect 390560 3392 390612 3398
rect 390560 3334 390612 3340
rect 390664 480 390692 32535
rect 391940 24268 391992 24274
rect 391940 24210 391992 24216
rect 391952 16574 391980 24210
rect 394712 16574 394740 61406
rect 391952 16546 392624 16574
rect 394712 16546 395384 16574
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391860 480 391888 3334
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394240 4004 394292 4010
rect 394240 3946 394292 3952
rect 394252 480 394280 3946
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 68410
rect 440240 68400 440292 68406
rect 440240 68342 440292 68348
rect 418804 65544 418856 65550
rect 418804 65486 418856 65492
rect 412638 60072 412694 60081
rect 412638 60007 412694 60016
rect 398840 56024 398892 56030
rect 398840 55966 398892 55972
rect 397736 4956 397788 4962
rect 397736 4898 397788 4904
rect 397748 480 397776 4898
rect 398852 3210 398880 55966
rect 402980 53168 403032 53174
rect 402980 53110 403032 53116
rect 400862 52048 400918 52057
rect 400862 51983 400918 51992
rect 398932 22976 398984 22982
rect 398932 22918 398984 22924
rect 398944 3398 398972 22918
rect 400876 3398 400904 51983
rect 402992 16574 403020 53110
rect 405738 47832 405794 47841
rect 405738 47767 405794 47776
rect 405752 16574 405780 47767
rect 408500 43512 408552 43518
rect 408500 43454 408552 43460
rect 407212 29776 407264 29782
rect 407212 29718 407264 29724
rect 402992 16546 403664 16574
rect 405752 16546 406056 16574
rect 401324 3936 401376 3942
rect 401324 3878 401376 3884
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400864 3392 400916 3398
rect 400864 3334 400916 3340
rect 398852 3182 398972 3210
rect 398944 480 398972 3182
rect 400140 480 400168 3334
rect 401336 480 401364 3878
rect 402520 3392 402572 3398
rect 402520 3334 402572 3340
rect 402532 480 402560 3334
rect 403636 480 403664 16546
rect 404360 14544 404412 14550
rect 404360 14486 404412 14492
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 14486
rect 406028 480 406056 16546
rect 407224 480 407252 29718
rect 408512 16574 408540 43454
rect 409880 39568 409932 39574
rect 409880 39510 409932 39516
rect 409892 16574 409920 39510
rect 410524 27056 410576 27062
rect 410524 26998 410576 27004
rect 408512 16546 409184 16574
rect 409892 16546 410472 16574
rect 408408 3868 408460 3874
rect 408408 3810 408460 3816
rect 408420 480 408448 3810
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410444 3482 410472 16546
rect 410536 3874 410564 26998
rect 410524 3868 410576 3874
rect 410524 3810 410576 3816
rect 411904 3868 411956 3874
rect 411904 3810 411956 3816
rect 410444 3454 410840 3482
rect 410812 480 410840 3454
rect 411916 480 411944 3810
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 60007
rect 414664 54596 414716 54602
rect 414664 54538 414716 54544
rect 414296 9036 414348 9042
rect 414296 8978 414348 8984
rect 414308 480 414336 8978
rect 414676 3398 414704 54538
rect 418160 25696 418212 25702
rect 418160 25638 418212 25644
rect 418172 16574 418200 25638
rect 418172 16546 418568 16574
rect 417424 11824 417476 11830
rect 417424 11766 417476 11772
rect 415492 3800 415544 3806
rect 415492 3742 415544 3748
rect 414664 3392 414716 3398
rect 414664 3334 414716 3340
rect 415504 480 415532 3742
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416700 480 416728 3334
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 11766
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 418816 3398 418844 65486
rect 430578 63064 430634 63073
rect 430578 62999 430634 63008
rect 422942 61568 422998 61577
rect 422942 61503 422998 61512
rect 420920 15972 420972 15978
rect 420920 15914 420972 15920
rect 418804 3392 418856 3398
rect 418804 3334 418856 3340
rect 420184 3392 420236 3398
rect 420184 3334 420236 3340
rect 420196 480 420224 3334
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 15914
rect 422576 3732 422628 3738
rect 422576 3674 422628 3680
rect 422588 480 422616 3674
rect 422956 3398 422984 61503
rect 423770 50416 423826 50425
rect 423770 50351 423826 50360
rect 422944 3392 422996 3398
rect 422944 3334 422996 3340
rect 423784 480 423812 50351
rect 425058 46336 425114 46345
rect 425058 46271 425114 46280
rect 425072 16574 425100 46271
rect 426440 42220 426492 42226
rect 426440 42162 426492 42168
rect 426452 16574 426480 42162
rect 427820 28416 427872 28422
rect 427820 28358 427872 28364
rect 427832 16574 427860 28358
rect 430592 16574 430620 62999
rect 432602 57352 432658 57361
rect 432602 57287 432658 57296
rect 431960 18760 432012 18766
rect 431960 18702 432012 18708
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 424980 480 425008 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 429660 3664 429712 3670
rect 429660 3606 429712 3612
rect 429672 480 429700 3606
rect 430868 480 430896 16546
rect 431972 3670 432000 18702
rect 432052 10396 432104 10402
rect 432052 10338 432104 10344
rect 431960 3664 432012 3670
rect 431960 3606 432012 3612
rect 432064 480 432092 10338
rect 432616 3398 432644 57287
rect 437478 53136 437534 53145
rect 437478 53071 437534 53080
rect 435548 7744 435600 7750
rect 435548 7686 435600 7692
rect 433248 3664 433300 3670
rect 433248 3606 433300 3612
rect 432604 3392 432656 3398
rect 432604 3334 432656 3340
rect 433260 480 433288 3606
rect 434444 3392 434496 3398
rect 434444 3334 434496 3340
rect 434456 480 434484 3334
rect 435560 480 435588 7686
rect 436744 6452 436796 6458
rect 436744 6394 436796 6400
rect 436756 480 436784 6394
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437492 354 437520 53071
rect 438860 42152 438912 42158
rect 438860 42094 438912 42100
rect 438872 16574 438900 42094
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 3398 440280 68342
rect 448520 58676 448572 58682
rect 448520 58618 448572 58624
rect 444378 44976 444434 44985
rect 444378 44911 444434 44920
rect 440332 22908 440384 22914
rect 440332 22850 440384 22856
rect 440240 3392 440292 3398
rect 440240 3334 440292 3340
rect 440344 480 440372 22850
rect 444392 16574 444420 44911
rect 446404 33992 446456 33998
rect 446404 33934 446456 33940
rect 445760 17400 445812 17406
rect 445760 17342 445812 17348
rect 444392 16546 445064 16574
rect 442632 7676 442684 7682
rect 442632 7618 442684 7624
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 441540 480 441568 3334
rect 442644 480 442672 7618
rect 443828 6384 443880 6390
rect 443828 6326 443880 6332
rect 443840 480 443868 6326
rect 445036 480 445064 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 17342
rect 446416 3398 446444 33934
rect 446404 3392 446456 3398
rect 446404 3334 446456 3340
rect 447416 3392 447468 3398
rect 447416 3334 447468 3340
rect 447428 480 447456 3334
rect 448532 3210 448560 58618
rect 448612 55956 448664 55962
rect 448612 55898 448664 55904
rect 448624 3398 448652 55898
rect 450542 51912 450598 51921
rect 450542 51847 450598 51856
rect 450556 4146 450584 51847
rect 450912 6316 450964 6322
rect 450912 6258 450964 6264
rect 450544 4140 450596 4146
rect 450544 4082 450596 4088
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 6258
rect 453316 6254 453344 77250
rect 454684 75268 454736 75274
rect 454684 75210 454736 75216
rect 454038 35184 454094 35193
rect 454038 35119 454094 35128
rect 453212 6248 453264 6254
rect 453212 6190 453264 6196
rect 453304 6248 453356 6254
rect 453304 6190 453356 6196
rect 452108 4140 452160 4146
rect 452108 4082 452160 4088
rect 452120 480 452148 4082
rect 453224 3210 453252 6190
rect 453224 3182 453344 3210
rect 453316 480 453344 3182
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454052 354 454080 35119
rect 454696 3670 454724 75210
rect 475384 74656 475436 74662
rect 475384 74598 475436 74604
rect 472624 64252 472676 64258
rect 472624 64194 472676 64200
rect 459560 59424 459612 59430
rect 459560 59366 459612 59372
rect 455418 49056 455474 49065
rect 455418 48991 455474 49000
rect 455432 16574 455460 48991
rect 458180 43444 458232 43450
rect 458180 43386 458232 43392
rect 456798 32464 456854 32473
rect 456798 32399 456854 32408
rect 455432 16546 455736 16574
rect 454684 3664 454736 3670
rect 454684 3606 454736 3612
rect 455708 480 455736 16546
rect 456812 3210 456840 32399
rect 456892 20052 456944 20058
rect 456892 19994 456944 20000
rect 456904 3398 456932 19994
rect 458192 16574 458220 43386
rect 459572 16574 459600 59366
rect 464344 54528 464396 54534
rect 464344 54470 464396 54476
rect 462320 40860 462372 40866
rect 462320 40802 462372 40808
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 456892 3392 456944 3398
rect 456892 3334 456944 3340
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 456812 3182 456932 3210
rect 456904 480 456932 3182
rect 458100 480 458128 3334
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461584 3596 461636 3602
rect 461584 3538 461636 3544
rect 461596 480 461624 3538
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 40802
rect 463700 38072 463752 38078
rect 463700 38014 463752 38020
rect 463712 16574 463740 38014
rect 463712 16546 464016 16574
rect 463988 480 464016 16546
rect 464356 3058 464384 54470
rect 466458 47696 466514 47705
rect 466458 47631 466514 47640
rect 466472 16574 466500 47631
rect 468482 47560 468538 47569
rect 468482 47495 468538 47504
rect 467840 35284 467892 35290
rect 467840 35226 467892 35232
rect 467852 16574 467880 35226
rect 466472 16546 467512 16574
rect 467852 16546 468248 16574
rect 465172 3460 465224 3466
rect 465172 3402 465224 3408
rect 464344 3052 464396 3058
rect 464344 2994 464396 3000
rect 465184 480 465212 3402
rect 466276 3052 466328 3058
rect 466276 2994 466328 3000
rect 466288 480 466316 2994
rect 467484 480 467512 16546
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 468496 3466 468524 47495
rect 470600 31068 470652 31074
rect 470600 31010 470652 31016
rect 468484 3460 468536 3466
rect 468484 3402 468536 3408
rect 469864 3460 469916 3466
rect 469864 3402 469916 3408
rect 469876 480 469904 3402
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 31010
rect 471980 21412 472032 21418
rect 471980 21354 472032 21360
rect 471992 16574 472020 21354
rect 471992 16546 472296 16574
rect 472268 480 472296 16546
rect 472636 3534 472664 64194
rect 473452 57248 473504 57254
rect 473452 57190 473504 57196
rect 473464 16574 473492 57190
rect 473464 16546 474136 16574
rect 472624 3528 472676 3534
rect 472624 3470 472676 3476
rect 473452 3528 473504 3534
rect 473452 3470 473504 3476
rect 473464 480 473492 3470
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475396 3534 475424 74598
rect 476120 38004 476172 38010
rect 476120 37946 476172 37952
rect 476132 16574 476160 37946
rect 477500 17332 477552 17338
rect 477500 17274 477552 17280
rect 477512 16574 477540 17274
rect 480272 16574 480300 79494
rect 500960 79484 501012 79490
rect 500960 79426 501012 79432
rect 486422 77888 486478 77897
rect 486422 77823 486478 77832
rect 480904 71052 480956 71058
rect 480904 70994 480956 71000
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 480272 16546 480576 16574
rect 475384 3528 475436 3534
rect 475384 3470 475436 3476
rect 475752 3460 475804 3466
rect 475752 3402 475804 3408
rect 475764 480 475792 3402
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478156 480 478184 16546
rect 479340 6248 479392 6254
rect 479340 6190 479392 6196
rect 479352 480 479380 6190
rect 480548 480 480576 16546
rect 480916 2922 480944 70994
rect 484398 46200 484454 46209
rect 484398 46135 484454 46144
rect 481640 36712 481692 36718
rect 481640 36654 481692 36660
rect 481652 16574 481680 36654
rect 484412 16574 484440 46135
rect 481652 16546 481772 16574
rect 484412 16546 484808 16574
rect 480904 2916 480956 2922
rect 480904 2858 480956 2864
rect 481744 480 481772 16546
rect 482836 4888 482888 4894
rect 482836 4830 482888 4836
rect 482848 480 482876 4830
rect 484032 2916 484084 2922
rect 484032 2858 484084 2864
rect 484044 480 484072 2858
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486436 13122 486464 77823
rect 493322 75304 493378 75313
rect 493322 75239 493378 75248
rect 489182 58712 489238 58721
rect 489182 58647 489238 58656
rect 486514 54496 486570 54505
rect 486514 54431 486570 54440
rect 486332 13116 486384 13122
rect 486332 13058 486384 13064
rect 486424 13116 486476 13122
rect 486424 13058 486476 13064
rect 486344 6914 486372 13058
rect 486344 6886 486464 6914
rect 486436 480 486464 6886
rect 486528 3534 486556 54431
rect 488540 33924 488592 33930
rect 488540 33866 488592 33872
rect 488552 16574 488580 33866
rect 488552 16546 488856 16574
rect 486516 3528 486568 3534
rect 486516 3470 486568 3476
rect 487620 3528 487672 3534
rect 487620 3470 487672 3476
rect 487632 480 487660 3470
rect 488828 480 488856 16546
rect 489196 3738 489224 58647
rect 490012 53100 490064 53106
rect 490012 53042 490064 53048
rect 490024 6914 490052 53042
rect 491300 29708 491352 29714
rect 491300 29650 491352 29656
rect 491312 16574 491340 29650
rect 491312 16546 492352 16574
rect 489932 6886 490052 6914
rect 489184 3732 489236 3738
rect 489184 3674 489236 3680
rect 489932 480 489960 6886
rect 491116 3732 491168 3738
rect 491116 3674 491168 3680
rect 491128 480 491156 3674
rect 492324 480 492352 16546
rect 493048 14476 493100 14482
rect 493048 14418 493100 14424
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 354 493088 14418
rect 493336 3534 493364 75239
rect 499580 75200 499632 75206
rect 499580 75142 499632 75148
rect 494058 71360 494114 71369
rect 494058 71295 494114 71304
rect 494072 16574 494100 71295
rect 498198 65648 498254 65657
rect 498198 65583 498254 65592
rect 495440 42084 495492 42090
rect 495440 42026 495492 42032
rect 494072 16546 494744 16574
rect 493324 3528 493376 3534
rect 493324 3470 493376 3476
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 42026
rect 497096 3664 497148 3670
rect 497096 3606 497148 3612
rect 497108 480 497136 3606
rect 498212 480 498240 65583
rect 498292 40792 498344 40798
rect 498292 40734 498344 40740
rect 498304 16574 498332 40734
rect 499592 16574 499620 75142
rect 500972 16574 501000 79426
rect 525800 79416 525852 79422
rect 525800 79358 525852 79364
rect 523132 79348 523184 79354
rect 523132 79290 523184 79296
rect 521658 75168 521714 75177
rect 521658 75103 521714 75112
rect 511264 74588 511316 74594
rect 511264 74530 511316 74536
rect 502982 69728 503038 69737
rect 502982 69663 503038 69672
rect 502340 28348 502392 28354
rect 502340 28290 502392 28296
rect 498304 16546 498976 16574
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500604 480 500632 16546
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502352 6914 502380 28290
rect 502996 16574 503024 69663
rect 507858 65512 507914 65521
rect 507858 65447 507914 65456
rect 503720 36644 503772 36650
rect 503720 36586 503772 36592
rect 502996 16546 503116 16574
rect 502352 6886 503024 6914
rect 502996 480 503024 6886
rect 503088 3058 503116 16546
rect 503076 3052 503128 3058
rect 503076 2994 503128 3000
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 36586
rect 506572 26988 506624 26994
rect 506572 26930 506624 26936
rect 506584 6914 506612 26930
rect 507872 16574 507900 65447
rect 510620 26920 510672 26926
rect 510620 26862 510672 26868
rect 509240 25628 509292 25634
rect 509240 25570 509292 25576
rect 509252 16574 509280 25570
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 506492 6886 506612 6914
rect 505376 3052 505428 3058
rect 505376 2994 505428 3000
rect 505388 480 505416 2994
rect 506492 480 506520 6886
rect 507676 3460 507728 3466
rect 507676 3402 507728 3408
rect 507688 480 507716 3402
rect 508884 480 508912 16546
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 510632 6914 510660 26862
rect 511276 16574 511304 74530
rect 511998 64152 512054 64161
rect 511998 64087 512054 64096
rect 511276 16546 511396 16574
rect 510632 6886 511304 6914
rect 511276 480 511304 6886
rect 511368 3466 511396 16546
rect 511356 3460 511408 3466
rect 511356 3402 511408 3408
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 64087
rect 514022 62928 514078 62937
rect 514022 62863 514078 62872
rect 513380 24200 513432 24206
rect 513380 24142 513432 24148
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 24142
rect 514036 3534 514064 62863
rect 520924 44192 520976 44198
rect 520924 44134 520976 44140
rect 518900 39500 518952 39506
rect 518900 39442 518952 39448
rect 516140 39432 516192 39438
rect 516140 39374 516192 39380
rect 516152 16574 516180 39374
rect 518912 16574 518940 39442
rect 520280 22840 520332 22846
rect 520280 22782 520332 22788
rect 516152 16546 517192 16574
rect 518912 16546 519584 16574
rect 514024 3528 514076 3534
rect 514024 3470 514076 3476
rect 515956 3528 516008 3534
rect 515956 3470 516008 3476
rect 514760 3460 514812 3466
rect 514760 3402 514812 3408
rect 514772 480 514800 3402
rect 515968 480 515996 3470
rect 517164 480 517192 16546
rect 518348 3392 518400 3398
rect 518348 3334 518400 3340
rect 518360 480 518388 3334
rect 519556 480 519584 16546
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 354 520320 22782
rect 520936 3330 520964 44134
rect 520924 3324 520976 3330
rect 520924 3266 520976 3272
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 75103
rect 523144 6914 523172 79290
rect 525064 37936 525116 37942
rect 525064 37878 525116 37884
rect 524420 25560 524472 25566
rect 524420 25502 524472 25508
rect 524432 16574 524460 25502
rect 524432 16546 525012 16574
rect 523052 6886 523172 6914
rect 523052 480 523080 6886
rect 524984 3482 525012 16546
rect 525076 3602 525104 37878
rect 525812 16574 525840 79358
rect 539692 78736 539744 78742
rect 539692 78678 539744 78684
rect 531318 71224 531374 71233
rect 531318 71159 531374 71168
rect 529940 61396 529992 61402
rect 529940 61338 529992 61344
rect 527822 59936 527878 59945
rect 527822 59871 527878 59880
rect 527836 16574 527864 59871
rect 528558 44840 528614 44849
rect 528558 44775 528614 44784
rect 525812 16546 526208 16574
rect 527836 16546 527956 16574
rect 525064 3596 525116 3602
rect 525064 3538 525116 3544
rect 524984 3454 525472 3482
rect 524236 3324 524288 3330
rect 524236 3266 524288 3272
rect 524248 480 524276 3266
rect 525444 480 525472 3454
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527824 3596 527876 3602
rect 527824 3538 527876 3544
rect 527836 480 527864 3538
rect 527928 3466 527956 16546
rect 527916 3460 527968 3466
rect 527916 3402 527968 3408
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 44775
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 61338
rect 531332 480 531360 71159
rect 536840 68332 536892 68338
rect 536840 68274 536892 68280
rect 535460 40724 535512 40730
rect 535460 40666 535512 40672
rect 534080 36576 534132 36582
rect 534080 36518 534132 36524
rect 531412 24132 531464 24138
rect 531412 24074 531464 24080
rect 531424 16574 531452 24074
rect 534092 16574 534120 36518
rect 535472 16574 535500 40666
rect 536852 16574 536880 68274
rect 538862 58576 538918 58585
rect 538862 58511 538918 58520
rect 531424 16546 532096 16574
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533712 3460 533764 3466
rect 533712 3402 533764 3408
rect 533724 480 533752 3402
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 538404 7608 538456 7614
rect 538404 7550 538456 7556
rect 538416 480 538444 7550
rect 538876 3194 538904 58511
rect 538956 22772 539008 22778
rect 538956 22714 539008 22720
rect 538968 3466 538996 22714
rect 539704 16574 539732 78678
rect 552662 76528 552718 76537
rect 552662 76463 552718 76472
rect 547878 71088 547934 71097
rect 547878 71023 547934 71032
rect 543740 64184 543792 64190
rect 543740 64126 543792 64132
rect 542358 51776 542414 51785
rect 542358 51711 542414 51720
rect 542372 16574 542400 51711
rect 543752 16574 543780 64126
rect 545762 57216 545818 57225
rect 545762 57151 545818 57160
rect 539704 16546 540376 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 538956 3460 539008 3466
rect 538956 3402 539008 3408
rect 539600 3460 539652 3466
rect 539600 3402 539652 3408
rect 538864 3188 538916 3194
rect 538864 3130 538916 3136
rect 539612 480 539640 3402
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540348 354 540376 16546
rect 541992 11756 542044 11762
rect 541992 11698 542044 11704
rect 542004 480 542032 11698
rect 540766 354 540878 480
rect 540348 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545488 4820 545540 4826
rect 545488 4762 545540 4768
rect 545500 480 545528 4762
rect 545776 3534 545804 57151
rect 545764 3528 545816 3534
rect 545764 3470 545816 3476
rect 546684 3188 546736 3194
rect 546684 3130 546736 3136
rect 546696 480 546724 3130
rect 547892 480 547920 71023
rect 549258 43480 549314 43489
rect 549258 43415 549314 43424
rect 549272 16574 549300 43415
rect 552020 35216 552072 35222
rect 552020 35158 552072 35164
rect 549272 16546 550312 16574
rect 548616 10328 548668 10334
rect 548616 10270 548668 10276
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548628 354 548656 10270
rect 550284 480 550312 16546
rect 552032 6914 552060 35158
rect 552676 16574 552704 76463
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 557538 69592 557594 69601
rect 557538 69527 557594 69536
rect 554044 66292 554096 66298
rect 554044 66234 554096 66240
rect 552676 16546 552796 16574
rect 552032 6886 552704 6914
rect 551468 3528 551520 3534
rect 551468 3470 551520 3476
rect 551480 480 551508 3470
rect 552676 480 552704 6886
rect 552768 3262 552796 16546
rect 554056 3534 554084 66234
rect 556158 48920 556214 48929
rect 556158 48855 556214 48864
rect 556172 16574 556200 48855
rect 557552 16574 557580 69527
rect 574742 68232 574798 68241
rect 574742 68167 574798 68176
rect 561678 62792 561734 62801
rect 561678 62727 561734 62736
rect 560942 50280 560998 50289
rect 560942 50215 560998 50224
rect 558920 39364 558972 39370
rect 558920 39306 558972 39312
rect 558932 16574 558960 39306
rect 556172 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 556160 8968 556212 8974
rect 556160 8910 556212 8916
rect 554044 3528 554096 3534
rect 554044 3470 554096 3476
rect 554964 3528 555016 3534
rect 554964 3470 555016 3476
rect 552756 3256 552808 3262
rect 552756 3198 552808 3204
rect 553768 3256 553820 3262
rect 553768 3198 553820 3204
rect 553780 480 553808 3198
rect 554976 480 555004 3470
rect 556172 480 556200 8910
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 560392 15904 560444 15910
rect 560392 15846 560444 15852
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 15846
rect 560956 3534 560984 50215
rect 561692 16574 561720 62727
rect 563702 61432 563758 61441
rect 563702 61367 563758 61376
rect 561692 16546 562088 16574
rect 560944 3528 560996 3534
rect 560944 3470 560996 3476
rect 562060 480 562088 16546
rect 563244 6180 563296 6186
rect 563244 6122 563296 6128
rect 563256 480 563284 6122
rect 563716 4146 563744 61367
rect 564532 55888 564584 55894
rect 564532 55830 564584 55836
rect 564544 16574 564572 55830
rect 569960 50380 570012 50386
rect 569960 50322 570012 50328
rect 565820 33856 565872 33862
rect 565820 33798 565872 33804
rect 565832 16574 565860 33798
rect 567200 18692 567252 18698
rect 567200 18634 567252 18640
rect 567212 16574 567240 18634
rect 569972 16574 570000 50322
rect 571984 46232 572036 46238
rect 571984 46174 572036 46180
rect 571340 18624 571392 18630
rect 571340 18566 571392 18572
rect 570604 17264 570656 17270
rect 570604 17206 570656 17212
rect 564544 16546 565216 16574
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 569972 16546 570368 16574
rect 563704 4140 563756 4146
rect 563704 4082 563756 4088
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564452 480 564480 3470
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 569132 4140 569184 4146
rect 569132 4082 569184 4088
rect 569144 480 569172 4082
rect 570340 480 570368 16546
rect 570616 3466 570644 17206
rect 570604 3460 570656 3466
rect 570604 3402 570656 3408
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 18566
rect 571996 3534 572024 46174
rect 574100 29640 574152 29646
rect 574100 29582 574152 29588
rect 574112 16574 574140 29582
rect 574112 16546 574692 16574
rect 571984 3528 572036 3534
rect 571984 3470 572036 3476
rect 573916 3528 573968 3534
rect 573916 3470 573968 3476
rect 574664 3482 574692 16546
rect 574756 3602 574784 68167
rect 576860 42832 576912 42838
rect 576860 42774 576912 42780
rect 576872 16574 576900 42774
rect 578240 33788 578292 33794
rect 578240 33730 578292 33736
rect 578252 16574 578280 33730
rect 576872 16546 576992 16574
rect 578252 16546 578648 16574
rect 574744 3596 574796 3602
rect 574744 3538 574796 3544
rect 576308 3596 576360 3602
rect 576308 3538 576360 3544
rect 572720 3460 572772 3466
rect 572720 3402 572772 3408
rect 572732 480 572760 3402
rect 573928 480 573956 3470
rect 574664 3454 575152 3482
rect 575124 480 575152 3454
rect 576320 480 576348 3538
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576964 354 576992 16546
rect 578620 480 578648 16546
rect 580276 6633 580304 150447
rect 580368 144226 580396 179143
rect 580540 150476 580592 150482
rect 580540 150418 580592 150424
rect 580356 144220 580408 144226
rect 580356 144162 580408 144168
rect 580354 142216 580410 142225
rect 580354 142151 580410 142160
rect 580368 19825 580396 142151
rect 580446 140856 580502 140865
rect 580446 140791 580502 140800
rect 580460 33153 580488 140791
rect 580552 46345 580580 150418
rect 580632 149116 580684 149122
rect 580632 149058 580684 149064
rect 580644 59673 580672 149058
rect 580816 142180 580868 142186
rect 580816 142122 580868 142128
rect 580722 140992 580778 141001
rect 580722 140927 580778 140936
rect 580736 112849 580764 140927
rect 580828 126041 580856 142122
rect 580814 126032 580870 126041
rect 580814 125967 580870 125976
rect 580722 112840 580778 112849
rect 580722 112775 580778 112784
rect 581000 73840 581052 73846
rect 581000 73782 581052 73788
rect 580630 59664 580686 59673
rect 580630 59599 580686 59608
rect 580538 46336 580594 46345
rect 580538 46271 580594 46280
rect 580446 33144 580502 33153
rect 580446 33079 580502 33088
rect 580354 19816 580410 19825
rect 580354 19751 580410 19760
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 581012 480 581040 73782
rect 582380 28280 582432 28286
rect 582380 28222 582432 28228
rect 582392 16574 582420 28222
rect 582392 16546 583432 16574
rect 581736 13116 581788 13122
rect 581736 13058 581788 13064
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 13058
rect 583404 480 583432 16546
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 2778 514820 2834 514856
rect 2778 514800 2780 514820
rect 2780 514800 2832 514820
rect 2832 514800 2834 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3146 449520 3202 449576
rect 2870 410488 2926 410544
rect 3146 358400 3202 358456
rect 3330 319232 3386 319288
rect 3514 462576 3570 462632
rect 3514 423544 3570 423600
rect 3514 397468 3516 397488
rect 3516 397468 3568 397488
rect 3568 397468 3570 397488
rect 3514 397432 3570 397468
rect 3514 371320 3570 371376
rect 3514 345344 3570 345400
rect 3514 306176 3570 306232
rect 3514 293120 3570 293176
rect 3054 267144 3110 267200
rect 3330 241068 3332 241088
rect 3332 241068 3384 241088
rect 3384 241068 3386 241088
rect 3330 241032 3386 241068
rect 2778 214920 2834 214976
rect 111430 262792 111486 262848
rect 3606 254088 3662 254144
rect 3514 201864 3570 201920
rect 3422 188808 3478 188864
rect 3514 162832 3570 162888
rect 3146 149776 3202 149832
rect 3238 136720 3294 136776
rect 2778 110608 2834 110664
rect 2778 77832 2834 77888
rect 3514 84632 3570 84688
rect 7562 75112 7618 75168
rect 3514 71612 3516 71632
rect 3516 71612 3568 71632
rect 3568 71612 3570 71632
rect 3514 71576 3570 71612
rect 4802 64096 4858 64152
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 8298 72392 8354 72448
rect 7654 66816 7710 66872
rect 17222 139440 17278 139496
rect 13082 76472 13138 76528
rect 9678 71168 9734 71224
rect 9034 71032 9090 71088
rect 12438 55800 12494 55856
rect 14462 73752 14518 73808
rect 18602 69536 18658 69592
rect 17958 53080 18014 53136
rect 26238 68176 26294 68232
rect 23478 61376 23534 61432
rect 25502 57160 25558 57216
rect 30378 50224 30434 50280
rect 39302 48864 39358 48920
rect 41418 54440 41474 54496
rect 44270 47504 44326 47560
rect 66258 76608 66314 76664
rect 49698 46144 49754 46200
rect 54482 73888 54538 73944
rect 59358 65592 59414 65648
rect 57978 65456 58034 65512
rect 57242 64232 57298 64288
rect 56598 55936 56654 55992
rect 63498 43424 63554 43480
rect 75182 61512 75238 61568
rect 74538 40568 74594 40624
rect 80058 57296 80114 57352
rect 84198 54576 84254 54632
rect 81438 51720 81494 51776
rect 92478 53760 92534 53816
rect 93858 58520 93914 58576
rect 95238 44784 95294 44840
rect 97538 192480 97594 192536
rect 96526 153720 96582 153776
rect 96250 41248 96306 41304
rect 96526 41248 96582 41304
rect 96526 40568 96582 40624
rect 96434 37168 96490 37224
rect 97354 75112 97410 75168
rect 97262 70216 97318 70272
rect 97722 192616 97778 192672
rect 103150 199280 103206 199336
rect 99286 199144 99342 199200
rect 98458 71576 98514 71632
rect 98458 71168 98514 71224
rect 97906 64776 97962 64832
rect 98734 76880 98790 76936
rect 98734 76472 98790 76528
rect 100574 195200 100630 195256
rect 99930 72936 99986 72992
rect 100206 151000 100262 151056
rect 100666 190984 100722 191040
rect 100298 62056 100354 62112
rect 100298 61376 100354 61432
rect 101218 138624 101274 138680
rect 101586 148280 101642 148336
rect 99470 50904 99526 50960
rect 100666 50904 100722 50960
rect 99470 50224 99526 50280
rect 100758 49544 100814 49600
rect 100758 48864 100814 48920
rect 102046 187040 102102 187096
rect 101954 55120 102010 55176
rect 101954 54440 102010 54496
rect 102598 138760 102654 138816
rect 102690 112376 102746 112432
rect 102046 49544 102102 49600
rect 100758 46824 100814 46880
rect 101586 46824 101642 46880
rect 100758 46144 100814 46200
rect 102782 69808 102838 69864
rect 102782 69556 102838 69592
rect 102782 69536 102784 69556
rect 102784 69536 102836 69556
rect 102836 69536 102838 69556
rect 102138 44104 102194 44160
rect 102690 44104 102746 44160
rect 102138 43424 102194 43480
rect 102138 37168 102194 37224
rect 102138 36488 102194 36544
rect 103058 76744 103114 76800
rect 103150 68856 103206 68912
rect 103150 68176 103206 68232
rect 103426 192888 103482 192944
rect 103978 113736 104034 113792
rect 103978 81096 104034 81152
rect 104622 195336 104678 195392
rect 104714 73072 104770 73128
rect 104622 72528 104678 72584
rect 104438 66156 104494 66192
rect 104438 66136 104440 66156
rect 104440 66136 104492 66156
rect 104492 66136 104494 66156
rect 104438 65592 104494 65648
rect 103794 64232 103850 64288
rect 103978 64096 104034 64152
rect 105542 189624 105598 189680
rect 105174 81368 105230 81424
rect 104898 71052 104954 71088
rect 104898 71032 104900 71052
rect 104900 71032 104952 71052
rect 104952 71032 104954 71052
rect 106002 191256 106058 191312
rect 106002 61512 106058 61568
rect 107198 190032 107254 190088
rect 107014 189896 107070 189952
rect 106186 187584 106242 187640
rect 106830 138896 106886 138952
rect 106278 73888 106334 73944
rect 106186 57840 106242 57896
rect 105450 53760 105506 53816
rect 107106 189760 107162 189816
rect 108118 79192 108174 79248
rect 108670 79192 108726 79248
rect 109498 123392 109554 123448
rect 109958 196560 110014 196616
rect 110142 66136 110198 66192
rect 111246 77152 111302 77208
rect 111154 75112 111210 75168
rect 110694 65864 110750 65920
rect 109590 54576 109646 54632
rect 112350 139304 112406 139360
rect 112258 80688 112314 80744
rect 112534 138488 112590 138544
rect 112718 75520 112774 75576
rect 112442 72664 112498 72720
rect 112810 71712 112866 71768
rect 113546 147464 113602 147520
rect 113178 138896 113234 138952
rect 113178 138352 113234 138408
rect 113270 74568 113326 74624
rect 113822 80824 113878 80880
rect 114466 75656 114522 75712
rect 115018 144472 115074 144528
rect 115018 110608 115074 110664
rect 115202 139168 115258 139224
rect 115202 75384 115258 75440
rect 116306 79464 116362 79520
rect 116214 78920 116270 78976
rect 116674 74160 116730 74216
rect 117870 150456 117926 150512
rect 117870 142024 117926 142080
rect 117778 80960 117834 81016
rect 117870 79056 117926 79112
rect 117686 74024 117742 74080
rect 119710 262656 119766 262712
rect 118330 141480 118386 141536
rect 118238 72664 118294 72720
rect 116858 71440 116914 71496
rect 118422 75248 118478 75304
rect 118330 68584 118386 68640
rect 119158 137808 119214 137864
rect 119158 80144 119214 80200
rect 120078 80552 120134 80608
rect 119802 78376 119858 78432
rect 117226 65456 117282 65512
rect 120814 262384 120870 262440
rect 120722 194520 120778 194576
rect 120814 138080 120870 138136
rect 120630 80416 120686 80472
rect 120630 72800 120686 72856
rect 116950 61784 117006 61840
rect 123758 259528 123814 259584
rect 135258 260208 135314 260264
rect 136224 260208 136280 260264
rect 140226 262520 140282 262576
rect 141422 263744 141478 263800
rect 142250 262792 142306 262848
rect 142802 262792 142858 262848
rect 143630 265104 143686 265160
rect 144182 265104 144238 265160
rect 143538 260208 143594 260264
rect 144504 260208 144560 260264
rect 145562 264968 145618 265024
rect 144918 259936 144974 259992
rect 146206 263608 146262 263664
rect 147770 260072 147826 260128
rect 150438 281560 150494 281616
rect 149702 262656 149758 262712
rect 152186 262792 152242 262848
rect 152186 262384 152242 262440
rect 149242 259800 149298 259856
rect 153290 289856 153346 289912
rect 153290 263608 153346 263664
rect 153290 263472 153346 263528
rect 155958 260208 156014 260264
rect 156648 260208 156704 260264
rect 146482 259664 146538 259720
rect 156786 259664 156842 259720
rect 160098 259936 160154 259992
rect 163410 263064 163466 263120
rect 162030 262520 162086 262576
rect 161478 260752 161534 260808
rect 160926 259936 160982 259992
rect 163410 262384 163466 262440
rect 162674 260752 162730 260808
rect 162582 259800 162638 259856
rect 163594 263064 163650 263120
rect 164376 260072 164432 260128
rect 167550 264968 167606 265024
rect 131394 259528 131450 259584
rect 185674 260208 185730 260264
rect 185674 259664 185730 259720
rect 185674 259392 185730 259448
rect 128726 200504 128782 200560
rect 127622 200096 127678 200152
rect 122102 199008 122158 199064
rect 122194 195608 122250 195664
rect 122102 138760 122158 138816
rect 122378 195744 122434 195800
rect 123574 148824 123630 148880
rect 122470 140800 122526 140856
rect 122378 139712 122434 139768
rect 122746 138760 122802 138816
rect 122286 138488 122342 138544
rect 123666 142024 123722 142080
rect 123942 138760 123998 138816
rect 123574 138352 123630 138408
rect 124862 142568 124918 142624
rect 124862 142160 124918 142216
rect 124218 140800 124274 140856
rect 124678 140800 124734 140856
rect 126426 195472 126482 195528
rect 126334 140528 126390 140584
rect 126610 194112 126666 194168
rect 127162 198192 127218 198248
rect 127438 141072 127494 141128
rect 127530 140936 127586 140992
rect 128726 199824 128782 199880
rect 127622 140256 127678 140312
rect 131946 200640 132002 200696
rect 129186 198736 129242 198792
rect 129278 198056 129334 198112
rect 129646 195336 129702 195392
rect 129738 193024 129794 193080
rect 130566 193160 130622 193216
rect 131854 199280 131910 199336
rect 130474 140256 130530 140312
rect 132222 200540 132224 200560
rect 132224 200540 132276 200560
rect 132276 200540 132278 200560
rect 132222 200504 132278 200540
rect 177946 200368 178002 200424
rect 132222 198872 132278 198928
rect 132038 193840 132094 193896
rect 131854 146240 131910 146296
rect 132406 198328 132462 198384
rect 133280 199824 133336 199880
rect 132130 148688 132186 148744
rect 132866 187176 132922 187232
rect 133648 199824 133704 199880
rect 133832 199824 133888 199880
rect 134016 199858 134072 199914
rect 133326 191120 133382 191176
rect 133786 199688 133842 199744
rect 134568 199824 134624 199880
rect 134752 199824 134808 199880
rect 133694 191392 133750 191448
rect 133878 199416 133934 199472
rect 133878 192888 133934 192944
rect 134384 199724 134386 199744
rect 134386 199724 134438 199744
rect 134438 199724 134440 199744
rect 134384 199688 134440 199724
rect 134522 199688 134578 199744
rect 134154 196424 134210 196480
rect 134614 195200 134670 195256
rect 134890 199688 134946 199744
rect 135120 199858 135176 199914
rect 135488 199858 135544 199914
rect 135764 199858 135820 199914
rect 135074 199552 135130 199608
rect 134982 199416 135038 199472
rect 131670 139984 131726 140040
rect 135534 196968 135590 197024
rect 135442 196832 135498 196888
rect 136408 199858 136464 199914
rect 135902 196016 135958 196072
rect 136454 199688 136510 199744
rect 136776 199858 136832 199914
rect 136730 199724 136732 199744
rect 136732 199724 136784 199744
rect 136784 199724 136786 199744
rect 136730 199688 136786 199724
rect 136454 198328 136510 198384
rect 136362 196696 136418 196752
rect 136178 195880 136234 195936
rect 136638 199552 136694 199608
rect 136822 198872 136878 198928
rect 137006 190304 137062 190360
rect 136822 190168 136878 190224
rect 137420 199858 137476 199914
rect 137374 196696 137430 196752
rect 137696 199858 137752 199914
rect 137650 199552 137706 199608
rect 138110 199588 138112 199608
rect 138112 199588 138164 199608
rect 138164 199588 138166 199608
rect 138110 199552 138166 199588
rect 138018 198872 138074 198928
rect 138616 199858 138672 199914
rect 138478 198600 138534 198656
rect 138662 199688 138718 199744
rect 138984 199858 139040 199914
rect 138570 198328 138626 198384
rect 136730 141344 136786 141400
rect 138846 198872 138902 198928
rect 139168 199858 139224 199914
rect 139030 199552 139086 199608
rect 139398 199708 139454 199744
rect 139812 199858 139868 199914
rect 139398 199688 139400 199708
rect 139400 199688 139452 199708
rect 139452 199688 139454 199708
rect 139398 199552 139454 199608
rect 139398 191528 139454 191584
rect 139582 199416 139638 199472
rect 140180 199858 140236 199914
rect 140456 199858 140512 199914
rect 139674 196696 139730 196752
rect 140042 196968 140098 197024
rect 140226 199688 140282 199744
rect 140226 196016 140282 196072
rect 140410 199688 140466 199744
rect 140640 199858 140696 199914
rect 140916 199858 140972 199914
rect 140410 196832 140466 196888
rect 140594 196832 140650 196888
rect 138662 147600 138718 147656
rect 140778 196424 140834 196480
rect 141468 199858 141524 199914
rect 141652 199858 141708 199914
rect 141606 199416 141662 199472
rect 141698 198192 141754 198248
rect 141514 196832 141570 196888
rect 142066 199688 142122 199744
rect 142250 199724 142252 199744
rect 142252 199724 142304 199744
rect 142304 199724 142306 199744
rect 142250 199688 142306 199724
rect 142664 199858 142720 199914
rect 142848 199858 142904 199914
rect 142158 199300 142214 199336
rect 142158 199280 142160 199300
rect 142160 199280 142212 199300
rect 142212 199280 142214 199300
rect 142158 199144 142214 199200
rect 139490 141480 139546 141536
rect 143032 199858 143088 199914
rect 142802 197376 142858 197432
rect 142710 196560 142766 196616
rect 143860 199858 143916 199914
rect 144412 199858 144468 199914
rect 142986 197376 143042 197432
rect 143354 199552 143410 199608
rect 143354 195608 143410 195664
rect 144688 199858 144744 199914
rect 143722 199436 143778 199472
rect 143722 199416 143724 199436
rect 143724 199416 143776 199436
rect 143776 199416 143778 199436
rect 143630 199144 143686 199200
rect 143630 199008 143686 199064
rect 143538 147328 143594 147384
rect 142158 147056 142214 147112
rect 144182 199416 144238 199472
rect 144550 198872 144606 198928
rect 144274 196016 144330 196072
rect 145010 199688 145066 199744
rect 144918 199144 144974 199200
rect 145424 199858 145480 199914
rect 145884 199858 145940 199914
rect 146068 199858 146124 199914
rect 145194 195744 145250 195800
rect 145378 199164 145434 199200
rect 145378 199144 145380 199164
rect 145380 199144 145432 199164
rect 145432 199144 145434 199164
rect 145746 199688 145802 199744
rect 146528 199858 146584 199914
rect 146896 199858 146952 199914
rect 146574 199688 146630 199744
rect 145746 198600 145802 198656
rect 146114 199144 146170 199200
rect 146482 199552 146538 199608
rect 146574 199416 146630 199472
rect 147264 199858 147320 199914
rect 147586 199688 147642 199744
rect 147126 199416 147182 199472
rect 142250 146104 142306 146160
rect 144366 145968 144422 146024
rect 146758 145832 146814 145888
rect 146298 145560 146354 145616
rect 145562 144744 145618 144800
rect 145102 143384 145158 143440
rect 146666 142976 146722 143032
rect 147494 196424 147550 196480
rect 147678 199280 147734 199336
rect 147586 195608 147642 195664
rect 147862 199416 147918 199472
rect 147586 186360 147642 186416
rect 146942 143248 146998 143304
rect 148644 199688 148700 199744
rect 148138 198464 148194 198520
rect 148874 199688 148930 199744
rect 149334 198328 149390 198384
rect 148322 143112 148378 143168
rect 150576 199858 150632 199914
rect 150438 199688 150494 199744
rect 151496 199858 151552 199914
rect 150898 198056 150954 198112
rect 149978 142840 150034 142896
rect 150806 148552 150862 148608
rect 151082 144608 151138 144664
rect 151450 199688 151506 199744
rect 151818 196968 151874 197024
rect 151726 195336 151782 195392
rect 151634 189488 151690 189544
rect 151910 144336 151966 144392
rect 152600 199858 152656 199914
rect 152370 198736 152426 198792
rect 152002 144064 152058 144120
rect 152554 195200 152610 195256
rect 153060 199858 153116 199914
rect 153428 199858 153484 199914
rect 153106 195472 153162 195528
rect 152830 186904 152886 186960
rect 153888 199858 153944 199914
rect 154348 199858 154404 199914
rect 153566 192752 153622 192808
rect 153382 148416 153438 148472
rect 153290 145696 153346 145752
rect 152462 144200 152518 144256
rect 152646 144064 152702 144120
rect 154118 199688 154174 199744
rect 153934 196560 153990 196616
rect 153750 187312 153806 187368
rect 154302 199688 154358 199744
rect 154808 199858 154864 199914
rect 155084 199858 155140 199914
rect 154118 192888 154174 192944
rect 154762 199688 154818 199744
rect 154394 193296 154450 193352
rect 154578 144336 154634 144392
rect 154302 144200 154358 144256
rect 154026 140120 154082 140176
rect 154854 193976 154910 194032
rect 156096 199858 156152 199914
rect 155590 199280 155646 199336
rect 156050 199688 156106 199744
rect 156326 199552 156382 199608
rect 157108 199858 157164 199914
rect 157752 199858 157808 199914
rect 158028 199858 158084 199914
rect 157016 199688 157072 199744
rect 156878 198056 156934 198112
rect 157062 199552 157118 199608
rect 158304 199858 158360 199914
rect 157798 199552 157854 199608
rect 157982 199688 158038 199744
rect 158672 199858 158728 199914
rect 157798 196016 157854 196072
rect 158396 199688 158452 199744
rect 159316 199858 159372 199914
rect 158810 199552 158866 199608
rect 158626 192480 158682 192536
rect 159086 199688 159142 199744
rect 159086 198328 159142 198384
rect 158994 195880 159050 195936
rect 160052 199858 160108 199914
rect 160420 199858 160476 199914
rect 159454 193160 159510 193216
rect 160098 199008 160154 199064
rect 160006 197920 160062 197976
rect 160282 196832 160338 196888
rect 161064 199858 161120 199914
rect 161248 199824 161304 199880
rect 160926 198736 160982 198792
rect 160834 197104 160890 197160
rect 161570 199688 161626 199744
rect 161110 196832 161166 196888
rect 160926 196696 160982 196752
rect 161570 195880 161626 195936
rect 157246 142840 157302 142896
rect 162168 199824 162224 199880
rect 162214 199688 162270 199744
rect 162720 199858 162776 199914
rect 162306 199552 162362 199608
rect 162030 198464 162086 198520
rect 162306 195628 162362 195664
rect 162306 195608 162308 195628
rect 162308 195608 162360 195628
rect 162360 195608 162362 195628
rect 162582 199688 162638 199744
rect 163180 199858 163236 199914
rect 162214 143112 162270 143168
rect 161110 141344 161166 141400
rect 163134 199688 163190 199744
rect 162858 196832 162914 196888
rect 163318 198872 163374 198928
rect 164008 199824 164064 199880
rect 163778 199552 163834 199608
rect 163686 196968 163742 197024
rect 163778 195744 163834 195800
rect 162766 144472 162822 144528
rect 162674 141480 162730 141536
rect 164146 199688 164202 199744
rect 164744 199858 164800 199914
rect 164422 199552 164478 199608
rect 165296 199858 165352 199914
rect 165480 199858 165536 199914
rect 165848 199824 165904 199880
rect 164606 199144 164662 199200
rect 165158 199552 165214 199608
rect 165342 199688 165398 199744
rect 166860 199824 166916 199880
rect 165894 199552 165950 199608
rect 163962 145832 164018 145888
rect 164146 144608 164202 144664
rect 163870 142976 163926 143032
rect 165986 196288 166042 196344
rect 166814 199588 166816 199608
rect 166816 199588 166868 199608
rect 166868 199588 166870 199608
rect 166814 199552 166870 199588
rect 166814 199144 166870 199200
rect 166998 198600 167054 198656
rect 167274 195880 167330 195936
rect 167964 199824 168020 199880
rect 167550 199008 167606 199064
rect 167918 199688 167974 199744
rect 167734 198600 167790 198656
rect 168240 199858 168296 199914
rect 167182 151136 167238 151192
rect 167090 148552 167146 148608
rect 166998 145696 167054 145752
rect 168608 199858 168664 199914
rect 168194 199552 168250 199608
rect 168884 199858 168940 199914
rect 169160 199858 169216 199914
rect 169436 199858 169492 199914
rect 168654 199724 168656 199744
rect 168656 199724 168708 199744
rect 168708 199724 168710 199744
rect 168654 199688 168710 199724
rect 168930 199688 168986 199744
rect 168746 197648 168802 197704
rect 169114 198872 169170 198928
rect 169206 198600 169262 198656
rect 168930 192752 168986 192808
rect 169390 198600 169446 198656
rect 169390 187040 169446 187096
rect 170080 199858 170136 199914
rect 170540 199858 170596 199914
rect 171000 199858 171056 199914
rect 171184 199858 171240 199914
rect 171644 199858 171700 199914
rect 170954 199552 171010 199608
rect 171138 198056 171194 198112
rect 170954 195880 171010 195936
rect 169942 147328 169998 147384
rect 171138 196424 171194 196480
rect 171138 193024 171194 193080
rect 171690 199416 171746 199472
rect 171690 199144 171746 199200
rect 171414 192616 171470 192672
rect 171782 196016 171838 196072
rect 172196 199858 172252 199914
rect 172380 199858 172436 199914
rect 172426 199688 172482 199744
rect 172058 198192 172114 198248
rect 171966 194112 172022 194168
rect 171230 147464 171286 147520
rect 171690 152360 171746 152416
rect 172932 199824 172988 199880
rect 172702 199688 172758 199744
rect 172426 197512 172482 197568
rect 171782 145968 171838 146024
rect 172978 199552 173034 199608
rect 173576 199858 173632 199914
rect 173760 199858 173816 199914
rect 174128 199858 174184 199914
rect 173990 199688 174046 199744
rect 174312 199858 174368 199914
rect 173530 194384 173586 194440
rect 173806 199552 173862 199608
rect 173714 199144 173770 199200
rect 173898 193840 173954 193896
rect 174680 199858 174736 199914
rect 174450 199572 174506 199608
rect 174450 199552 174452 199572
rect 174452 199552 174504 199572
rect 174504 199552 174506 199572
rect 174634 199552 174690 199608
rect 174358 199144 174414 199200
rect 175140 199858 175196 199914
rect 175002 198464 175058 198520
rect 174910 195880 174966 195936
rect 175968 199858 176024 199914
rect 176244 199858 176300 199914
rect 175186 195472 175242 195528
rect 172794 149776 172850 149832
rect 172610 149640 172666 149696
rect 175554 199008 175610 199064
rect 175830 198872 175886 198928
rect 176014 198736 176070 198792
rect 175646 152768 175702 152824
rect 175462 150048 175518 150104
rect 175278 149912 175334 149968
rect 176888 199858 176944 199914
rect 176290 195608 176346 195664
rect 176842 198464 176898 198520
rect 177670 198600 177726 198656
rect 177854 199416 177910 199472
rect 179510 199824 179566 199880
rect 178406 197784 178462 197840
rect 177026 157936 177082 157992
rect 176934 155352 176990 155408
rect 176842 152360 176898 152416
rect 179602 199280 179658 199336
rect 178774 140120 178830 140176
rect 180522 200096 180578 200152
rect 180522 199552 180578 199608
rect 180338 146104 180394 146160
rect 181350 199416 181406 199472
rect 180614 193976 180670 194032
rect 180430 144744 180486 144800
rect 181442 140392 181498 140448
rect 187146 200096 187202 200152
rect 182822 140256 182878 140312
rect 182638 139576 182694 139632
rect 183190 147600 183246 147656
rect 183466 142724 183522 142760
rect 183466 142704 183468 142724
rect 183468 142704 183520 142724
rect 183520 142704 183522 142724
rect 183650 141208 183706 141264
rect 183006 139440 183062 139496
rect 184846 141208 184902 141264
rect 185490 139848 185546 139904
rect 185398 139576 185454 139632
rect 185950 155760 186006 155816
rect 185766 139712 185822 139768
rect 126242 139304 126298 139360
rect 130566 139304 130622 139360
rect 149426 139304 149482 139360
rect 175002 139304 175058 139360
rect 184110 139304 184166 139360
rect 184386 139304 184442 139360
rect 187054 155624 187110 155680
rect 185950 139304 186006 139360
rect 187790 212472 187846 212528
rect 187698 144200 187754 144256
rect 186502 139340 186504 139360
rect 186504 139340 186556 139360
rect 186556 139340 186558 139360
rect 186502 139304 186558 139340
rect 187054 139304 187110 139360
rect 124034 138080 124090 138136
rect 189170 142840 189226 142896
rect 189538 260072 189594 260128
rect 189446 259936 189502 259992
rect 122746 137944 122802 138000
rect 188894 137944 188950 138000
rect 188158 137828 188214 137864
rect 188158 137808 188160 137828
rect 188160 137808 188212 137828
rect 188212 137808 188214 137828
rect 122746 128424 122802 128480
rect 122746 122848 122802 122904
rect 122746 84088 122802 84144
rect 122194 80552 122250 80608
rect 120906 71168 120962 71224
rect 122378 80144 122434 80200
rect 124034 81096 124090 81152
rect 124034 80552 124090 80608
rect 129002 80552 129058 80608
rect 122746 75792 122802 75848
rect 123114 75792 123170 75848
rect 128266 79872 128322 79928
rect 127806 79328 127862 79384
rect 127806 78784 127862 78840
rect 128174 78784 128230 78840
rect 127070 77968 127126 78024
rect 127162 77832 127218 77888
rect 128266 78512 128322 78568
rect 128634 76880 128690 76936
rect 181626 80552 181682 80608
rect 130290 80144 130346 80200
rect 129738 75112 129794 75168
rect 130382 73752 130438 73808
rect 130474 72936 130530 72992
rect 130750 77696 130806 77752
rect 130934 75112 130990 75168
rect 178222 80416 178278 80472
rect 178406 80416 178462 80472
rect 132314 79756 132370 79792
rect 132314 79736 132316 79756
rect 132316 79736 132368 79756
rect 132368 79736 132370 79756
rect 131762 73072 131818 73128
rect 132544 79872 132600 79928
rect 132912 79906 132968 79962
rect 132958 79736 133014 79792
rect 133556 79906 133612 79962
rect 133740 79906 133796 79962
rect 134016 79906 134072 79962
rect 134200 79906 134256 79962
rect 133326 79736 133382 79792
rect 132866 77560 132922 77616
rect 133740 79736 133796 79792
rect 133418 77424 133474 77480
rect 134154 79736 134210 79792
rect 133602 77288 133658 77344
rect 132866 71576 132922 71632
rect 134568 79906 134624 79962
rect 135028 79906 135084 79962
rect 135304 79872 135360 79928
rect 135580 79872 135636 79928
rect 133970 77968 134026 78024
rect 133970 72392 134026 72448
rect 134614 77288 134670 77344
rect 134706 76608 134762 76664
rect 136224 79838 136280 79894
rect 135810 77424 135866 77480
rect 136960 79906 137016 79962
rect 137144 79872 137200 79928
rect 136914 79772 136916 79792
rect 136916 79772 136968 79792
rect 136968 79772 136970 79792
rect 136914 79736 136970 79772
rect 137512 79872 137568 79928
rect 137466 79736 137522 79792
rect 136914 79600 136970 79656
rect 137006 79328 137062 79384
rect 136822 78240 136878 78296
rect 136822 78104 136878 78160
rect 137190 79600 137246 79656
rect 137374 78648 137430 78704
rect 137466 76744 137522 76800
rect 137880 79872 137936 79928
rect 138018 76064 138074 76120
rect 138110 75112 138166 75168
rect 138616 79872 138672 79928
rect 139076 79906 139132 79962
rect 138846 79464 138902 79520
rect 138662 76064 138718 76120
rect 139122 79636 139124 79656
rect 139124 79636 139176 79656
rect 139176 79636 139178 79656
rect 139122 79600 139178 79636
rect 139536 79872 139592 79928
rect 139904 79872 139960 79928
rect 139122 79328 139178 79384
rect 138938 77832 138994 77888
rect 138754 75792 138810 75848
rect 139306 78104 139362 78160
rect 139766 78240 139822 78296
rect 139674 76200 139730 76256
rect 140042 79600 140098 79656
rect 140364 79872 140420 79928
rect 140916 79872 140972 79928
rect 140686 79464 140742 79520
rect 140778 78648 140834 78704
rect 140870 77696 140926 77752
rect 141468 79906 141524 79962
rect 142296 79906 142352 79962
rect 141238 79192 141294 79248
rect 141422 79192 141478 79248
rect 141330 75112 141386 75168
rect 142664 79906 142720 79962
rect 142848 79906 142904 79962
rect 142250 79192 142306 79248
rect 142526 79484 142582 79520
rect 142802 79600 142858 79656
rect 143308 79906 143364 79962
rect 142526 79464 142528 79484
rect 142528 79464 142580 79484
rect 142580 79464 142582 79484
rect 142250 78260 142306 78296
rect 142250 78240 142252 78260
rect 142252 78240 142304 78260
rect 142304 78240 142306 78260
rect 142710 79364 142712 79384
rect 142712 79364 142764 79384
rect 142764 79364 142766 79384
rect 142710 79328 142766 79364
rect 143170 79600 143226 79656
rect 142434 77288 142490 77344
rect 142342 73752 142398 73808
rect 142986 77288 143042 77344
rect 143170 79464 143226 79520
rect 143768 79906 143824 79962
rect 144044 79906 144100 79962
rect 144228 79906 144284 79962
rect 144688 79892 144744 79928
rect 144688 79872 144690 79892
rect 144690 79872 144742 79892
rect 144742 79872 144744 79892
rect 143354 77016 143410 77072
rect 143722 79464 143778 79520
rect 144090 77424 144146 77480
rect 143998 77288 144054 77344
rect 145056 79906 145112 79962
rect 145424 79872 145480 79928
rect 144274 78376 144330 78432
rect 144458 77560 144514 77616
rect 145700 79906 145756 79962
rect 147264 79906 147320 79962
rect 145010 79464 145066 79520
rect 144734 76880 144790 76936
rect 144550 74976 144606 75032
rect 145194 78784 145250 78840
rect 145378 76200 145434 76256
rect 145746 78648 145802 78704
rect 146206 75112 146262 75168
rect 147448 79906 147504 79962
rect 147724 79906 147780 79962
rect 146666 79636 146668 79656
rect 146668 79636 146720 79656
rect 146720 79636 146722 79656
rect 146666 79600 146722 79636
rect 146482 75248 146538 75304
rect 146758 79192 146814 79248
rect 146482 71032 146538 71088
rect 147908 79906 147964 79962
rect 147494 76200 147550 76256
rect 147678 79600 147734 79656
rect 148046 79636 148048 79656
rect 148048 79636 148100 79656
rect 148100 79636 148102 79656
rect 148046 79600 148102 79636
rect 147770 79328 147826 79384
rect 147954 79328 148010 79384
rect 147586 75384 147642 75440
rect 147862 79228 147864 79248
rect 147864 79228 147916 79248
rect 147916 79228 147918 79248
rect 147862 79192 147918 79228
rect 147954 77424 148010 77480
rect 148414 77424 148470 77480
rect 148690 77288 148746 77344
rect 149012 79906 149068 79962
rect 149380 79906 149436 79962
rect 148966 79620 149022 79656
rect 148966 79600 148968 79620
rect 148968 79600 149020 79620
rect 149020 79600 149022 79620
rect 148874 79464 148930 79520
rect 149426 78376 149482 78432
rect 150208 79872 150264 79928
rect 150852 79872 150908 79928
rect 150530 79056 150586 79112
rect 150438 78648 150494 78704
rect 151312 79906 151368 79962
rect 150254 78512 150310 78568
rect 149794 56480 149850 56536
rect 151496 79736 151552 79792
rect 151772 79872 151828 79928
rect 151450 79500 151452 79520
rect 151452 79500 151504 79520
rect 151504 79500 151506 79520
rect 151450 79464 151506 79500
rect 150622 69672 150678 69728
rect 150622 68992 150678 69048
rect 151634 79328 151690 79384
rect 151726 79056 151782 79112
rect 151726 78648 151782 78704
rect 151450 68992 151506 69048
rect 152324 79872 152380 79928
rect 152600 79872 152656 79928
rect 152784 79906 152840 79962
rect 152278 79736 152334 79792
rect 152186 77152 152242 77208
rect 152554 79736 152610 79792
rect 153060 79872 153116 79928
rect 153612 79906 153668 79962
rect 152462 77696 152518 77752
rect 153290 79736 153346 79792
rect 152554 77288 152610 77344
rect 152002 73072 152058 73128
rect 151910 46144 151966 46200
rect 152738 79600 152794 79656
rect 152646 76744 152702 76800
rect 152554 74024 152610 74080
rect 152554 73072 152610 73128
rect 153106 77288 153162 77344
rect 152922 74704 152978 74760
rect 153888 79872 153944 79928
rect 154256 79906 154312 79962
rect 154026 79736 154082 79792
rect 154394 79736 154450 79792
rect 154716 79872 154772 79928
rect 155268 79906 155324 79962
rect 153566 67496 153622 67552
rect 153566 66272 153622 66328
rect 153198 64776 153254 64832
rect 154026 79464 154082 79520
rect 154026 74432 154082 74488
rect 154118 70080 154174 70136
rect 153934 66272 153990 66328
rect 154486 76336 154542 76392
rect 154486 74432 154542 74488
rect 154210 69944 154266 70000
rect 154210 68992 154266 69048
rect 154394 68992 154450 69048
rect 154302 64776 154358 64832
rect 154762 79600 154818 79656
rect 154670 77152 154726 77208
rect 155314 79736 155370 79792
rect 154854 64504 154910 64560
rect 155958 78920 156014 78976
rect 156464 79872 156520 79928
rect 156142 79464 156198 79520
rect 157016 79872 157072 79928
rect 157200 79872 157256 79928
rect 156970 78512 157026 78568
rect 156602 66000 156658 66056
rect 157568 79906 157624 79962
rect 157752 79872 157808 79928
rect 158396 79906 158452 79962
rect 158120 79770 158176 79826
rect 158304 79772 158306 79792
rect 158306 79772 158358 79792
rect 158358 79772 158360 79792
rect 157890 79600 157946 79656
rect 157798 79464 157854 79520
rect 158304 79736 158360 79772
rect 157982 79192 158038 79248
rect 158534 78512 158590 78568
rect 158856 79736 158912 79792
rect 158718 79464 158774 79520
rect 159086 79600 159142 79656
rect 158810 78512 158866 78568
rect 159592 79908 159594 79928
rect 159594 79908 159646 79928
rect 159646 79908 159648 79928
rect 159592 79872 159648 79908
rect 160052 79872 160108 79928
rect 159454 79600 159510 79656
rect 160420 79872 160476 79928
rect 160880 79872 160936 79928
rect 160834 79736 160890 79792
rect 160972 79736 161028 79792
rect 160834 79464 160890 79520
rect 160834 77016 160890 77072
rect 161110 77424 161166 77480
rect 161386 78512 161442 78568
rect 161110 15816 161166 15872
rect 160098 7520 160154 7576
rect 162260 79906 162316 79962
rect 162628 79906 162684 79962
rect 161478 67496 161534 67552
rect 162490 79636 162492 79656
rect 162492 79636 162544 79656
rect 162544 79636 162546 79656
rect 162490 79600 162546 79636
rect 162582 79192 162638 79248
rect 162858 79600 162914 79656
rect 162950 79192 163006 79248
rect 162766 77152 162822 77208
rect 162674 76472 162730 76528
rect 162490 67496 162546 67552
rect 163640 79906 163696 79962
rect 164008 79872 164064 79928
rect 163502 79600 163558 79656
rect 164284 79906 164340 79962
rect 164468 79906 164524 79962
rect 164928 79872 164984 79928
rect 163686 79464 163742 79520
rect 163870 75928 163926 75984
rect 164146 79056 164202 79112
rect 164698 78104 164754 78160
rect 164790 76880 164846 76936
rect 165664 79872 165720 79928
rect 165848 79872 165904 79928
rect 166124 79906 166180 79962
rect 164698 69944 164754 70000
rect 165526 79192 165582 79248
rect 165434 78920 165490 78976
rect 165618 78240 165674 78296
rect 166584 79736 166640 79792
rect 167228 79838 167284 79894
rect 165342 75928 165398 75984
rect 165802 75928 165858 75984
rect 166538 79600 166594 79656
rect 166630 78512 166686 78568
rect 166952 79736 167008 79792
rect 167688 79906 167744 79962
rect 166998 78512 167054 78568
rect 166998 75928 167054 75984
rect 167274 79600 167330 79656
rect 167274 79328 167330 79384
rect 167366 78376 167422 78432
rect 168056 79872 168112 79928
rect 168608 79872 168664 79928
rect 168792 79906 168848 79962
rect 167872 79736 167928 79792
rect 167734 75928 167790 75984
rect 168378 79736 168434 79792
rect 168562 79736 168618 79792
rect 169436 79872 169492 79928
rect 169620 79872 169676 79928
rect 169804 79872 169860 79928
rect 169022 79736 169078 79792
rect 168746 78920 168802 78976
rect 168930 79484 168986 79520
rect 168930 79464 168932 79484
rect 168932 79464 168984 79484
rect 168984 79464 168986 79484
rect 168838 78512 168894 78568
rect 168930 78240 168986 78296
rect 169390 79736 169446 79792
rect 169758 79736 169814 79792
rect 170080 79736 170136 79792
rect 169114 77832 169170 77888
rect 168930 75248 168986 75304
rect 170448 79906 170504 79962
rect 170632 79906 170688 79962
rect 171000 79872 171056 79928
rect 170954 79736 171010 79792
rect 171460 79872 171516 79928
rect 169574 77968 169630 78024
rect 169482 75248 169538 75304
rect 169114 72392 169170 72448
rect 168746 67360 168802 67416
rect 169666 67360 169722 67416
rect 170218 79600 170274 79656
rect 170126 78376 170182 78432
rect 170402 76608 170458 76664
rect 170126 76472 170182 76528
rect 170586 78512 170642 78568
rect 170494 76472 170550 76528
rect 170678 71712 170734 71768
rect 171230 79736 171286 79792
rect 171322 79600 171378 79656
rect 171046 76064 171102 76120
rect 171414 78512 171470 78568
rect 172150 79736 172206 79792
rect 171874 78104 171930 78160
rect 171966 77696 172022 77752
rect 171598 76472 171654 76528
rect 172150 76472 172206 76528
rect 172840 79872 172896 79928
rect 172702 79736 172758 79792
rect 172334 76472 172390 76528
rect 172242 75792 172298 75848
rect 172242 75248 172298 75304
rect 173116 79736 173172 79792
rect 172794 79600 172850 79656
rect 172702 78376 172758 78432
rect 173392 79736 173448 79792
rect 173668 79872 173724 79928
rect 174128 79906 174184 79962
rect 173852 79736 173908 79792
rect 174128 79770 174184 79826
rect 174404 79872 174460 79928
rect 174772 79872 174828 79928
rect 172886 78920 172942 78976
rect 173438 77696 173494 77752
rect 173254 75656 173310 75712
rect 173438 71576 173494 71632
rect 173714 78376 173770 78432
rect 173990 78376 174046 78432
rect 173162 22616 173218 22672
rect 174266 78920 174322 78976
rect 174266 72800 174322 72856
rect 175048 79872 175104 79928
rect 175600 79906 175656 79962
rect 176060 79906 176116 79962
rect 175784 79838 175840 79894
rect 176244 79872 176300 79928
rect 174634 79600 174690 79656
rect 174818 76880 174874 76936
rect 174726 76472 174782 76528
rect 174450 72800 174506 72856
rect 175232 79736 175288 79792
rect 175094 76472 175150 76528
rect 175186 75520 175242 75576
rect 175002 71304 175058 71360
rect 177440 79872 177496 79928
rect 175554 79600 175610 79656
rect 175738 79600 175794 79656
rect 176106 76880 176162 76936
rect 176198 76472 176254 76528
rect 176290 76200 176346 76256
rect 176106 75520 176162 75576
rect 175922 72800 175978 72856
rect 175554 70080 175610 70136
rect 176198 74840 176254 74896
rect 176290 74024 176346 74080
rect 176198 72528 176254 72584
rect 176382 72800 176438 72856
rect 176566 76472 176622 76528
rect 176474 72528 176530 72584
rect 177302 74840 177358 74896
rect 177578 78240 177634 78296
rect 177118 68856 177174 68912
rect 177946 77424 178002 77480
rect 177762 71440 177818 71496
rect 178222 78920 178278 78976
rect 181626 80280 181682 80336
rect 178314 78104 178370 78160
rect 178222 76880 178278 76936
rect 178038 74976 178094 75032
rect 178038 71032 178094 71088
rect 180522 79872 180578 79928
rect 181442 78512 181498 78568
rect 181626 78512 181682 78568
rect 180522 78376 180578 78432
rect 181442 78104 181498 78160
rect 183558 77424 183614 77480
rect 188894 80280 188950 80336
rect 188986 78512 189042 78568
rect 188342 65456 188398 65512
rect 189446 143112 189502 143168
rect 189538 110608 189594 110664
rect 189538 107072 189594 107128
rect 189630 51992 189686 52048
rect 191010 259800 191066 259856
rect 191010 142976 191066 143032
rect 191286 109112 191342 109168
rect 191838 43424 191894 43480
rect 192298 260208 192354 260264
rect 192482 72392 192538 72448
rect 191930 39888 191986 39944
rect 193034 39888 193090 39944
rect 193034 39208 193090 39264
rect 193678 140700 193680 140720
rect 193680 140700 193732 140720
rect 193732 140700 193734 140720
rect 193678 140664 193734 140700
rect 193862 139304 193918 139360
rect 194598 197104 194654 197160
rect 194046 141344 194102 141400
rect 194046 139984 194102 140040
rect 194046 75112 194102 75168
rect 193678 60580 193734 60616
rect 193678 60560 193680 60580
rect 193680 60560 193732 60580
rect 193732 60560 193734 60580
rect 193586 52128 193642 52184
rect 193310 50224 193366 50280
rect 194506 138080 194562 138136
rect 195978 195744 196034 195800
rect 195426 152632 195482 152688
rect 195242 139168 195298 139224
rect 195518 145560 195574 145616
rect 194598 54848 194654 54904
rect 194598 54576 194654 54632
rect 196714 146920 196770 146976
rect 196162 82184 196218 82240
rect 196622 138624 196678 138680
rect 196806 113872 196862 113928
rect 196070 53624 196126 53680
rect 195978 49408 196034 49464
rect 195978 49136 196034 49192
rect 197450 196968 197506 197024
rect 197358 77968 197414 78024
rect 197450 52400 197506 52456
rect 198738 197240 198794 197296
rect 197818 138896 197874 138952
rect 198094 114416 198150 114472
rect 197910 78512 197966 78568
rect 197450 51992 197506 52048
rect 197450 48048 197506 48104
rect 197450 47776 197506 47832
rect 199106 139032 199162 139088
rect 199014 78512 199070 78568
rect 199566 138760 199622 138816
rect 199474 81504 199530 81560
rect 200394 196696 200450 196752
rect 199106 62056 199162 62112
rect 199842 62056 199898 62112
rect 199842 61512 199898 61568
rect 198738 50632 198794 50688
rect 200946 137808 201002 137864
rect 201314 80008 201370 80064
rect 201406 78104 201462 78160
rect 200394 63008 200450 63064
rect 200302 57704 200358 57760
rect 201866 158072 201922 158128
rect 201958 151000 202014 151056
rect 201682 52264 201738 52320
rect 200210 45328 200266 45384
rect 201406 45328 201462 45384
rect 201406 44920 201462 44976
rect 202970 192752 203026 192808
rect 202786 52264 202842 52320
rect 202786 51856 202842 51912
rect 202418 49544 202474 49600
rect 202786 49544 202842 49600
rect 202786 49000 202842 49056
rect 203338 155488 203394 155544
rect 203246 148280 203302 148336
rect 203338 48184 203394 48240
rect 202970 47912 203026 47968
rect 204718 147056 204774 147112
rect 204166 48184 204222 48240
rect 204074 47912 204130 47968
rect 204166 47640 204222 47696
rect 204074 47504 204130 47560
rect 204718 46144 204774 46200
rect 204718 41248 204774 41304
rect 204718 40568 204774 40624
rect 204994 80824 205050 80880
rect 205546 75792 205602 75848
rect 204902 74024 204958 74080
rect 205914 192616 205970 192672
rect 204902 67496 204958 67552
rect 205914 45500 205916 45520
rect 205916 45500 205968 45520
rect 205968 45500 205970 45520
rect 205914 45464 205970 45500
rect 204810 35808 204866 35864
rect 204810 35264 204866 35320
rect 206374 80688 206430 80744
rect 206282 75792 206338 75848
rect 205730 30232 205786 30288
rect 206006 30232 206062 30288
rect 205730 29552 205786 29608
rect 207294 200232 207350 200288
rect 207110 75248 207166 75304
rect 207110 74976 207166 75032
rect 347042 290400 347098 290456
rect 396722 282104 396778 282160
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580262 365064 580318 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 325216 580226 325272
rect 579986 312024 580042 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 412638 262792 412694 262848
rect 471242 259528 471298 259584
rect 580170 258848 580226 258904
rect 579710 245556 579712 245576
rect 579712 245556 579764 245576
rect 579764 245556 579766 245576
rect 579710 245520 579766 245556
rect 580170 205672 580226 205728
rect 209962 200096 210018 200152
rect 208490 193976 208546 194032
rect 208398 190032 208454 190088
rect 207478 75248 207534 75304
rect 207386 75112 207442 75168
rect 207846 81096 207902 81152
rect 207754 80960 207810 81016
rect 207018 21800 207074 21856
rect 207938 72528 207994 72584
rect 209870 191120 209926 191176
rect 209778 189896 209834 189952
rect 208766 72664 208822 72720
rect 208582 58520 208638 58576
rect 208490 51720 208546 51776
rect 208398 44104 208454 44160
rect 208398 43424 208454 43480
rect 208398 30912 208454 30968
rect 209870 32952 209926 33008
rect 209778 21256 209834 21312
rect 210054 55120 210110 55176
rect 210054 54440 210110 54496
rect 210330 72800 210386 72856
rect 211158 189760 211214 189816
rect 210514 76880 210570 76936
rect 211066 76880 211122 76936
rect 211066 76472 211122 76528
rect 210146 48864 210202 48920
rect 210146 44124 210202 44160
rect 210146 44104 210148 44124
rect 210148 44104 210200 44124
rect 210200 44104 210202 44124
rect 212538 198328 212594 198384
rect 211434 71440 211490 71496
rect 212630 193840 212686 193896
rect 213918 198192 213974 198248
rect 212630 60424 212686 60480
rect 213826 60424 213882 60480
rect 213826 59880 213882 59936
rect 211250 54984 211306 55040
rect 211250 54440 211306 54496
rect 214010 198056 214066 198112
rect 214194 197920 214250 197976
rect 214102 186904 214158 186960
rect 214010 66000 214066 66056
rect 214010 62736 214066 62792
rect 212538 28192 212594 28248
rect 211158 17856 211214 17912
rect 212446 17856 212502 17912
rect 212446 17176 212502 17232
rect 214286 65456 214342 65512
rect 214470 69672 214526 69728
rect 214746 71712 214802 71768
rect 214746 71304 214802 71360
rect 214194 58656 214250 58712
rect 215758 195336 215814 195392
rect 215574 155216 215630 155272
rect 215390 59064 215446 59120
rect 215298 53760 215354 53816
rect 215298 53352 215354 53408
rect 214102 35672 214158 35728
rect 214102 35128 214158 35184
rect 216678 192480 216734 192536
rect 215758 74160 215814 74216
rect 215666 66136 215722 66192
rect 215574 33088 215630 33144
rect 215574 32408 215630 32464
rect 216678 21936 216734 21992
rect 217322 198736 217378 198792
rect 217138 195608 217194 195664
rect 217046 59200 217102 59256
rect 217230 195472 217286 195528
rect 218150 196560 218206 196616
rect 217966 76880 218022 76936
rect 219438 190984 219494 191040
rect 218518 152496 218574 152552
rect 218334 77016 218390 77072
rect 218518 77016 218574 77072
rect 218518 76880 218574 76936
rect 218334 76608 218390 76664
rect 218702 78784 218758 78840
rect 218518 76336 218574 76392
rect 218150 74296 218206 74352
rect 218150 73888 218206 73944
rect 217598 63416 217654 63472
rect 217322 63280 217378 63336
rect 217322 62736 217378 62792
rect 217230 57840 217286 57896
rect 217230 57160 217286 57216
rect 216954 50904 217010 50960
rect 216862 38528 216918 38584
rect 217046 38528 217102 38584
rect 217046 37848 217102 37904
rect 219622 72936 219678 72992
rect 220910 195200 220966 195256
rect 219530 60288 219586 60344
rect 219438 46688 219494 46744
rect 221002 73072 221058 73128
rect 221278 189624 221334 189680
rect 580538 232328 580594 232384
rect 580446 219000 580502 219056
rect 580354 192480 580410 192536
rect 580354 179152 580410 179208
rect 580170 165824 580226 165880
rect 580078 152632 580134 152688
rect 580262 150456 580318 150512
rect 482282 141072 482338 141128
rect 221278 73616 221334 73672
rect 221278 73208 221334 73264
rect 234618 78648 234674 78704
rect 221462 77968 221518 78024
rect 222106 77968 222162 78024
rect 222106 77288 222162 77344
rect 224222 73208 224278 73264
rect 220910 46824 220966 46880
rect 227718 66816 227774 66872
rect 230478 61648 230534 61704
rect 229098 40704 229154 40760
rect 231858 45192 231914 45248
rect 237378 74024 237434 74080
rect 247682 76880 247738 76936
rect 245658 63144 245714 63200
rect 249798 58928 249854 58984
rect 268382 78104 268438 78160
rect 260838 76744 260894 76800
rect 255318 73888 255374 73944
rect 259550 46416 259606 46472
rect 261482 73752 261538 73808
rect 266358 18536 266414 18592
rect 276110 39208 276166 39264
rect 281538 58792 281594 58848
rect 284390 53352 284446 53408
rect 295338 65728 295394 65784
rect 293958 37848 294014 37904
rect 303618 35264 303674 35320
rect 318798 72528 318854 72584
rect 315302 54712 315358 54768
rect 316130 17176 316186 17232
rect 579802 139304 579858 139360
rect 579618 99456 579674 99512
rect 579618 86128 579674 86184
rect 342902 77968 342958 78024
rect 324318 40568 324374 40624
rect 332598 72392 332654 72448
rect 333978 29552 334034 29608
rect 336738 21528 336794 21584
rect 367098 76608 367154 76664
rect 342994 21392 343050 21448
rect 347778 21256 347834 21312
rect 356058 49272 356114 49328
rect 364982 54576 365038 54632
rect 369858 52128 369914 52184
rect 373998 50496 374054 50552
rect 382922 53216 382978 53272
rect 387798 49136 387854 49192
rect 390558 45056 390614 45112
rect 390650 32544 390706 32600
rect 412638 60016 412694 60072
rect 400862 51992 400918 52048
rect 405738 47776 405794 47832
rect 430578 63008 430634 63064
rect 422942 61512 422998 61568
rect 423770 50360 423826 50416
rect 425058 46280 425114 46336
rect 432602 57296 432658 57352
rect 437478 53080 437534 53136
rect 444378 44920 444434 44976
rect 450542 51856 450598 51912
rect 454038 35128 454094 35184
rect 455418 49000 455474 49056
rect 456798 32408 456854 32464
rect 466458 47640 466514 47696
rect 468482 47504 468538 47560
rect 486422 77832 486478 77888
rect 484398 46144 484454 46200
rect 493322 75248 493378 75304
rect 489182 58656 489238 58712
rect 486514 54440 486570 54496
rect 494058 71304 494114 71360
rect 498198 65592 498254 65648
rect 521658 75112 521714 75168
rect 502982 69672 503038 69728
rect 507858 65456 507914 65512
rect 511998 64096 512054 64152
rect 514022 62872 514078 62928
rect 531318 71168 531374 71224
rect 527822 59880 527878 59936
rect 528558 44784 528614 44840
rect 538862 58520 538918 58576
rect 552662 76472 552718 76528
rect 547878 71032 547934 71088
rect 542358 51720 542414 51776
rect 545762 57160 545818 57216
rect 549258 43424 549314 43480
rect 580170 72936 580226 72992
rect 557538 69536 557594 69592
rect 556158 48864 556214 48920
rect 574742 68176 574798 68232
rect 561678 62736 561734 62792
rect 560942 50224 560998 50280
rect 563702 61376 563758 61432
rect 580354 142160 580410 142216
rect 580446 140800 580502 140856
rect 580722 140936 580778 140992
rect 580814 125976 580870 126032
rect 580722 112784 580778 112840
rect 580630 59608 580686 59664
rect 580538 46280 580594 46336
rect 580446 33088 580502 33144
rect 580354 19760 580410 19816
rect 580262 6568 580318 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 2773 514858 2839 514861
rect -960 514856 2839 514858
rect -960 514800 2778 514856
rect 2834 514800 2839 514856
rect -960 514798 2839 514800
rect -960 514708 480 514798
rect 2773 514795 2839 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect -960 371318 3575 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 580257 365122 580323 365125
rect 583520 365122 584960 365212
rect 580257 365120 584960 365122
rect 580257 365064 580262 365120
rect 580318 365064 584960 365120
rect 580257 365062 584960 365064
rect 580257 365059 580323 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3509 345402 3575 345405
rect -960 345400 3575 345402
rect -960 345344 3514 345400
rect 3570 345344 3575 345400
rect -960 345342 3575 345344
rect -960 345252 480 345342
rect 3509 345339 3575 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 347037 290458 347103 290461
rect 190410 290456 347103 290458
rect 190410 290400 347042 290456
rect 347098 290400 347103 290456
rect 190410 290398 347103 290400
rect 153285 289914 153351 289917
rect 189022 289914 189028 289916
rect 153285 289912 189028 289914
rect 153285 289856 153290 289912
rect 153346 289856 189028 289912
rect 153285 289854 189028 289856
rect 153285 289851 153351 289854
rect 189022 289852 189028 289854
rect 189092 289914 189098 289916
rect 190410 289914 190470 290398
rect 347037 290395 347103 290398
rect 189092 289854 190470 289914
rect 189092 289852 189098 289854
rect 583520 285276 584960 285516
rect 396717 282162 396783 282165
rect 190410 282160 396783 282162
rect 190410 282104 396722 282160
rect 396778 282104 396783 282160
rect 190410 282102 396783 282104
rect 150433 281618 150499 281621
rect 186998 281618 187004 281620
rect 150433 281616 187004 281618
rect 150433 281560 150438 281616
rect 150494 281560 187004 281616
rect 150433 281558 187004 281560
rect 150433 281555 150499 281558
rect 186998 281556 187004 281558
rect 187068 281618 187074 281620
rect 190410 281618 190470 282102
rect 396717 282099 396783 282102
rect 187068 281558 190470 281618
rect 187068 281556 187074 281558
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 111558 265100 111564 265164
rect 111628 265162 111634 265164
rect 143625 265162 143691 265165
rect 144177 265162 144243 265165
rect 111628 265160 144243 265162
rect 111628 265104 143630 265160
rect 143686 265104 144182 265160
rect 144238 265104 144243 265160
rect 111628 265102 144243 265104
rect 111628 265100 111634 265102
rect 143625 265099 143691 265102
rect 144177 265099 144243 265102
rect 111374 264964 111380 265028
rect 111444 265026 111450 265028
rect 145557 265026 145623 265029
rect 111444 265024 145623 265026
rect 111444 264968 145562 265024
rect 145618 264968 145623 265024
rect 111444 264966 145623 264968
rect 111444 264964 111450 264966
rect 145557 264963 145623 264966
rect 167545 265026 167611 265029
rect 198774 265026 198780 265028
rect 167545 265024 198780 265026
rect 167545 264968 167550 265024
rect 167606 264968 198780 265024
rect 167545 264966 198780 264968
rect 167545 264963 167611 264966
rect 198774 264964 198780 264966
rect 198844 264964 198850 265028
rect 115790 263740 115796 263804
rect 115860 263802 115866 263804
rect 141417 263802 141483 263805
rect 115860 263800 141483 263802
rect 115860 263744 141422 263800
rect 141478 263744 141483 263800
rect 115860 263742 141483 263744
rect 115860 263740 115866 263742
rect 141417 263739 141483 263742
rect 117078 263604 117084 263668
rect 117148 263666 117154 263668
rect 146201 263666 146267 263669
rect 117148 263664 146267 263666
rect 117148 263608 146206 263664
rect 146262 263608 146267 263664
rect 117148 263606 146267 263608
rect 117148 263604 117154 263606
rect 146201 263603 146267 263606
rect 153285 263666 153351 263669
rect 153285 263664 153394 263666
rect 153285 263608 153290 263664
rect 153346 263608 153394 263664
rect 153285 263603 153394 263608
rect 153334 263533 153394 263603
rect 153285 263528 153394 263533
rect 153285 263472 153290 263528
rect 153346 263472 153394 263528
rect 153285 263470 153394 263472
rect 153285 263467 153351 263470
rect 163405 263122 163471 263125
rect 163589 263122 163655 263125
rect 163405 263120 163655 263122
rect 163405 263064 163410 263120
rect 163466 263064 163594 263120
rect 163650 263064 163655 263120
rect 163405 263062 163655 263064
rect 163405 263059 163471 263062
rect 163589 263059 163655 263062
rect 111425 262850 111491 262853
rect 142245 262850 142311 262853
rect 142797 262850 142863 262853
rect 111425 262848 142863 262850
rect 111425 262792 111430 262848
rect 111486 262792 142250 262848
rect 142306 262792 142802 262848
rect 142858 262792 142863 262848
rect 111425 262790 142863 262792
rect 111425 262787 111491 262790
rect 142245 262787 142311 262790
rect 142797 262787 142863 262790
rect 152181 262850 152247 262853
rect 412633 262850 412699 262853
rect 152181 262848 412699 262850
rect 152181 262792 152186 262848
rect 152242 262792 412638 262848
rect 412694 262792 412699 262848
rect 152181 262790 412699 262792
rect 152181 262787 152247 262790
rect 412633 262787 412699 262790
rect 119705 262714 119771 262717
rect 149697 262714 149763 262717
rect 119705 262712 149763 262714
rect 119705 262656 119710 262712
rect 119766 262656 149702 262712
rect 149758 262656 149763 262712
rect 119705 262654 149763 262656
rect 119705 262651 119771 262654
rect 149697 262651 149763 262654
rect 109534 262516 109540 262580
rect 109604 262578 109610 262580
rect 140221 262578 140287 262581
rect 109604 262576 140287 262578
rect 109604 262520 140226 262576
rect 140282 262520 140287 262576
rect 109604 262518 140287 262520
rect 109604 262516 109610 262518
rect 140221 262515 140287 262518
rect 162025 262578 162091 262581
rect 193438 262578 193444 262580
rect 162025 262576 193444 262578
rect 162025 262520 162030 262576
rect 162086 262520 193444 262576
rect 162025 262518 193444 262520
rect 162025 262515 162091 262518
rect 193438 262516 193444 262518
rect 193508 262516 193514 262580
rect 120809 262442 120875 262445
rect 152181 262442 152247 262445
rect 120809 262440 152247 262442
rect 120809 262384 120814 262440
rect 120870 262384 152186 262440
rect 152242 262384 152247 262440
rect 120809 262382 152247 262384
rect 120809 262379 120875 262382
rect 152181 262379 152247 262382
rect 163405 262442 163471 262445
rect 193254 262442 193260 262444
rect 163405 262440 193260 262442
rect 163405 262384 163410 262440
rect 163466 262384 193260 262440
rect 163405 262382 193260 262384
rect 163405 262379 163471 262382
rect 193254 262380 193260 262382
rect 193324 262380 193330 262444
rect 161473 260810 161539 260813
rect 162669 260810 162735 260813
rect 161473 260808 162735 260810
rect 161473 260752 161478 260808
rect 161534 260752 162674 260808
rect 162730 260752 162735 260808
rect 161473 260750 162735 260752
rect 161473 260747 161539 260750
rect 162669 260747 162735 260750
rect 118366 260340 118372 260404
rect 118436 260402 118442 260404
rect 118436 260342 142170 260402
rect 118436 260340 118442 260342
rect 114134 260204 114140 260268
rect 114204 260266 114210 260268
rect 135253 260266 135319 260269
rect 136219 260266 136285 260269
rect 114204 260264 136285 260266
rect 114204 260208 135258 260264
rect 135314 260208 136224 260264
rect 136280 260208 136285 260264
rect 114204 260206 136285 260208
rect 142110 260266 142170 260342
rect 143533 260266 143599 260269
rect 144499 260266 144565 260269
rect 142110 260264 144565 260266
rect 142110 260208 143538 260264
rect 143594 260208 144504 260264
rect 144560 260208 144565 260264
rect 142110 260206 144565 260208
rect 114204 260204 114210 260206
rect 135253 260203 135319 260206
rect 136219 260203 136285 260206
rect 143533 260203 143599 260206
rect 144499 260203 144565 260206
rect 155953 260266 156019 260269
rect 156643 260266 156709 260269
rect 155953 260264 156709 260266
rect 155953 260208 155958 260264
rect 156014 260208 156648 260264
rect 156704 260208 156709 260264
rect 155953 260206 156709 260208
rect 155953 260203 156019 260206
rect 156643 260203 156709 260206
rect 185669 260266 185735 260269
rect 192293 260266 192359 260269
rect 185669 260264 192359 260266
rect 185669 260208 185674 260264
rect 185730 260208 192298 260264
rect 192354 260208 192359 260264
rect 185669 260206 192359 260208
rect 185669 260203 185735 260206
rect 192293 260203 192359 260206
rect 118550 260068 118556 260132
rect 118620 260130 118626 260132
rect 147765 260130 147831 260133
rect 118620 260128 147831 260130
rect 118620 260072 147770 260128
rect 147826 260072 147831 260128
rect 118620 260070 147831 260072
rect 118620 260068 118626 260070
rect 147765 260067 147831 260070
rect 164371 260130 164437 260133
rect 189533 260130 189599 260133
rect 164371 260128 189599 260130
rect 164371 260072 164376 260128
rect 164432 260072 189538 260128
rect 189594 260072 189599 260128
rect 164371 260070 189599 260072
rect 164371 260067 164437 260070
rect 189533 260067 189599 260070
rect 113030 259932 113036 259996
rect 113100 259994 113106 259996
rect 144913 259994 144979 259997
rect 113100 259992 144979 259994
rect 113100 259936 144918 259992
rect 144974 259936 144979 259992
rect 113100 259934 144979 259936
rect 113100 259932 113106 259934
rect 144913 259931 144979 259934
rect 160093 259994 160159 259997
rect 160921 259994 160987 259997
rect 189441 259994 189507 259997
rect 160093 259992 189507 259994
rect 160093 259936 160098 259992
rect 160154 259936 160926 259992
rect 160982 259936 189446 259992
rect 189502 259936 189507 259992
rect 160093 259934 189507 259936
rect 160093 259931 160159 259934
rect 160921 259931 160987 259934
rect 189441 259931 189507 259934
rect 116894 259796 116900 259860
rect 116964 259858 116970 259860
rect 149237 259858 149303 259861
rect 116964 259856 149303 259858
rect 116964 259800 149242 259856
rect 149298 259800 149303 259856
rect 116964 259798 149303 259800
rect 116964 259796 116970 259798
rect 149237 259795 149303 259798
rect 162577 259858 162643 259861
rect 191005 259858 191071 259861
rect 162577 259856 191071 259858
rect 162577 259800 162582 259856
rect 162638 259800 191010 259856
rect 191066 259800 191071 259856
rect 162577 259798 191071 259800
rect 162577 259795 162643 259798
rect 191005 259795 191071 259798
rect 113950 259660 113956 259724
rect 114020 259722 114026 259724
rect 146477 259722 146543 259725
rect 114020 259720 146543 259722
rect 114020 259664 146482 259720
rect 146538 259664 146543 259720
rect 114020 259662 146543 259664
rect 114020 259660 114026 259662
rect 146477 259659 146543 259662
rect 156781 259722 156847 259725
rect 185669 259722 185735 259725
rect 156781 259720 185735 259722
rect 156781 259664 156786 259720
rect 156842 259664 185674 259720
rect 185730 259664 185735 259720
rect 156781 259662 185735 259664
rect 156781 259659 156847 259662
rect 185669 259659 185735 259662
rect 111190 259524 111196 259588
rect 111260 259586 111266 259588
rect 123753 259586 123819 259589
rect 111260 259584 123819 259586
rect 111260 259528 123758 259584
rect 123814 259528 123819 259584
rect 111260 259526 123819 259528
rect 111260 259524 111266 259526
rect 123753 259523 123819 259526
rect 131389 259586 131455 259589
rect 471237 259586 471303 259589
rect 131389 259584 471303 259586
rect 131389 259528 131394 259584
rect 131450 259528 471242 259584
rect 471298 259528 471303 259584
rect 131389 259526 471303 259528
rect 131389 259523 131455 259526
rect 471237 259523 471303 259526
rect 185669 259450 185735 259453
rect 186078 259450 186084 259452
rect 185669 259448 186084 259450
rect 185669 259392 185674 259448
rect 185730 259392 186084 259448
rect 185669 259390 186084 259392
rect 185669 259387 185735 259390
rect 186078 259388 186084 259390
rect 186148 259388 186154 259452
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3601 254146 3667 254149
rect -960 254144 3667 254146
rect -960 254088 3606 254144
rect 3662 254088 3667 254144
rect -960 254086 3667 254088
rect -960 253996 480 254086
rect 3601 254083 3667 254086
rect 579705 245578 579771 245581
rect 583520 245578 584960 245668
rect 579705 245576 584960 245578
rect 579705 245520 579710 245576
rect 579766 245520 584960 245576
rect 579705 245518 584960 245520
rect 579705 245515 579771 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3325 241090 3391 241093
rect -960 241088 3391 241090
rect -960 241032 3330 241088
rect 3386 241032 3391 241088
rect -960 241030 3391 241032
rect -960 240940 480 241030
rect 3325 241027 3391 241030
rect 580533 232386 580599 232389
rect 583520 232386 584960 232476
rect 580533 232384 584960 232386
rect 580533 232328 580538 232384
rect 580594 232328 584960 232384
rect 580533 232326 584960 232328
rect 580533 232323 580599 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580441 219058 580507 219061
rect 583520 219058 584960 219148
rect 580441 219056 584960 219058
rect 580441 219000 580446 219056
rect 580502 219000 584960 219056
rect 580441 218998 584960 219000
rect 580441 218995 580507 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 2773 214978 2839 214981
rect -960 214976 2839 214978
rect -960 214920 2778 214976
rect 2834 214920 2839 214976
rect -960 214918 2839 214920
rect -960 214828 480 214918
rect 2773 214915 2839 214918
rect 186078 212468 186084 212532
rect 186148 212530 186154 212532
rect 187785 212530 187851 212533
rect 186148 212528 187851 212530
rect 186148 212472 187790 212528
rect 187846 212472 187851 212528
rect 186148 212470 187851 212472
rect 186148 212468 186154 212470
rect 187785 212467 187851 212470
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3509 201922 3575 201925
rect -960 201920 3575 201922
rect -960 201864 3514 201920
rect 3570 201864 3575 201920
rect -960 201862 3575 201864
rect -960 201772 480 201862
rect 3509 201859 3575 201862
rect 131941 200698 132007 200701
rect 137870 200698 137876 200700
rect 131941 200696 137876 200698
rect 131941 200640 131946 200696
rect 132002 200640 137876 200696
rect 131941 200638 137876 200640
rect 131941 200635 132007 200638
rect 137870 200636 137876 200638
rect 137940 200636 137946 200700
rect 103094 200500 103100 200564
rect 103164 200562 103170 200564
rect 128721 200562 128787 200565
rect 103164 200560 128787 200562
rect 103164 200504 128726 200560
rect 128782 200504 128787 200560
rect 103164 200502 128787 200504
rect 103164 200500 103170 200502
rect 128721 200499 128787 200502
rect 132217 200562 132283 200565
rect 136030 200562 136036 200564
rect 132217 200560 136036 200562
rect 132217 200504 132222 200560
rect 132278 200504 136036 200560
rect 132217 200502 136036 200504
rect 132217 200499 132283 200502
rect 136030 200500 136036 200502
rect 136100 200500 136106 200564
rect 102726 200364 102732 200428
rect 102796 200426 102802 200428
rect 102796 200366 118710 200426
rect 102796 200364 102802 200366
rect 118650 200290 118710 200366
rect 171358 200364 171364 200428
rect 171428 200426 171434 200428
rect 177941 200426 178007 200429
rect 171428 200424 178007 200426
rect 171428 200368 177946 200424
rect 178002 200368 178007 200424
rect 171428 200366 178007 200368
rect 171428 200364 171434 200366
rect 177941 200363 178007 200366
rect 207289 200290 207355 200293
rect 118650 200230 124230 200290
rect 124170 200018 124230 200230
rect 173988 200288 207355 200290
rect 173988 200232 207294 200288
rect 207350 200232 207355 200288
rect 173988 200230 207355 200232
rect 127617 200154 127683 200157
rect 127617 200152 152658 200154
rect 127617 200096 127622 200152
rect 127678 200096 152658 200152
rect 127617 200094 152658 200096
rect 127617 200091 127683 200094
rect 124170 199958 133522 200018
rect 128721 199882 128787 199885
rect 133275 199882 133341 199885
rect 128721 199880 133341 199882
rect 128721 199824 128726 199880
rect 128782 199824 133280 199880
rect 133336 199824 133341 199880
rect 128721 199822 133341 199824
rect 133462 199882 133522 199958
rect 139342 199956 139348 200020
rect 139412 199956 139418 200020
rect 134011 199914 134077 199919
rect 133643 199882 133709 199885
rect 133462 199880 133709 199882
rect 133462 199824 133648 199880
rect 133704 199824 133709 199880
rect 133462 199822 133709 199824
rect 128721 199819 128787 199822
rect 133275 199819 133341 199822
rect 133643 199819 133709 199822
rect 133827 199880 133893 199885
rect 133827 199824 133832 199880
rect 133888 199824 133893 199880
rect 134011 199858 134016 199914
rect 134072 199858 134077 199914
rect 135115 199914 135181 199919
rect 134011 199853 134077 199858
rect 134563 199880 134629 199885
rect 134747 199884 134813 199885
rect 133827 199819 133893 199824
rect 133830 199749 133890 199819
rect 133781 199744 133890 199749
rect 133781 199688 133786 199744
rect 133842 199688 133890 199744
rect 133781 199686 133890 199688
rect 133781 199683 133847 199686
rect 134014 199610 134074 199853
rect 134563 199824 134568 199880
rect 134624 199824 134629 199880
rect 134563 199819 134629 199824
rect 134742 199820 134748 199884
rect 134812 199882 134818 199884
rect 134812 199822 134904 199882
rect 135115 199858 135120 199914
rect 135176 199858 135181 199914
rect 135483 199914 135549 199919
rect 135483 199884 135488 199914
rect 135544 199884 135549 199914
rect 135759 199916 135825 199919
rect 135759 199914 135960 199916
rect 135115 199853 135181 199858
rect 134812 199820 134818 199822
rect 134747 199819 134813 199820
rect 134566 199749 134626 199819
rect 134190 199684 134196 199748
rect 134260 199746 134266 199748
rect 134379 199746 134445 199749
rect 134260 199744 134445 199746
rect 134260 199688 134384 199744
rect 134440 199688 134445 199744
rect 134260 199686 134445 199688
rect 134260 199684 134266 199686
rect 134379 199683 134445 199686
rect 134517 199744 134626 199749
rect 134885 199746 134951 199749
rect 134517 199688 134522 199744
rect 134578 199688 134626 199744
rect 134517 199686 134626 199688
rect 134750 199744 134951 199746
rect 134750 199688 134890 199744
rect 134946 199688 134951 199744
rect 134750 199686 134951 199688
rect 134517 199683 134583 199686
rect 125550 199550 134074 199610
rect 103145 199338 103211 199341
rect 125550 199338 125610 199550
rect 133873 199474 133939 199477
rect 134750 199474 134810 199686
rect 134885 199683 134951 199686
rect 135118 199613 135178 199853
rect 135478 199820 135484 199884
rect 135548 199882 135554 199884
rect 135548 199822 135606 199882
rect 135759 199858 135764 199914
rect 135820 199858 135960 199914
rect 136403 199914 136469 199919
rect 136403 199884 136408 199914
rect 136464 199884 136469 199914
rect 136771 199914 136837 199919
rect 137415 199916 137481 199919
rect 136771 199884 136776 199914
rect 136832 199884 136837 199914
rect 137142 199914 137481 199916
rect 135759 199856 135960 199858
rect 135759 199853 135825 199856
rect 135548 199820 135554 199822
rect 135069 199608 135178 199613
rect 135069 199552 135074 199608
rect 135130 199552 135178 199608
rect 135069 199550 135178 199552
rect 135069 199547 135135 199550
rect 133873 199472 134810 199474
rect 133873 199416 133878 199472
rect 133934 199416 134810 199472
rect 133873 199414 134810 199416
rect 134977 199474 135043 199477
rect 135900 199474 135960 199856
rect 136398 199820 136404 199884
rect 136468 199882 136474 199884
rect 136468 199822 136526 199882
rect 136468 199820 136474 199822
rect 136766 199820 136772 199884
rect 136836 199882 136842 199884
rect 136836 199822 136894 199882
rect 137142 199858 137420 199914
rect 137476 199858 137481 199914
rect 137142 199856 137481 199858
rect 136836 199820 136842 199822
rect 136030 199684 136036 199748
rect 136100 199746 136106 199748
rect 136449 199746 136515 199749
rect 136725 199746 136791 199749
rect 136100 199744 136515 199746
rect 136100 199688 136454 199744
rect 136510 199688 136515 199744
rect 136100 199686 136515 199688
rect 136100 199684 136106 199686
rect 136449 199683 136515 199686
rect 136590 199744 136791 199746
rect 136590 199688 136730 199744
rect 136786 199688 136791 199744
rect 136590 199686 136791 199688
rect 136590 199613 136650 199686
rect 136725 199683 136791 199686
rect 136590 199608 136699 199613
rect 136590 199552 136638 199608
rect 136694 199552 136699 199608
rect 136590 199550 136699 199552
rect 136633 199547 136699 199550
rect 134977 199472 135960 199474
rect 134977 199416 134982 199472
rect 135038 199416 135960 199472
rect 134977 199414 135960 199416
rect 133873 199411 133939 199414
rect 134977 199411 135043 199414
rect 103145 199336 125610 199338
rect 103145 199280 103150 199336
rect 103206 199280 125610 199336
rect 103145 199278 125610 199280
rect 131849 199338 131915 199341
rect 137142 199338 137202 199856
rect 137415 199853 137481 199856
rect 137691 199914 137757 199919
rect 137691 199858 137696 199914
rect 137752 199858 137757 199914
rect 138611 199914 138677 199919
rect 137691 199853 137757 199858
rect 137694 199613 137754 199853
rect 138238 199820 138244 199884
rect 138308 199882 138314 199884
rect 138611 199882 138616 199914
rect 138308 199858 138616 199882
rect 138672 199858 138677 199914
rect 138308 199853 138677 199858
rect 138979 199914 139045 199919
rect 138979 199858 138984 199914
rect 139040 199858 139045 199914
rect 139163 199914 139229 199919
rect 139163 199884 139168 199914
rect 139224 199884 139229 199914
rect 138979 199853 139045 199858
rect 138308 199822 138674 199853
rect 138308 199820 138314 199822
rect 138054 199684 138060 199748
rect 138124 199746 138130 199748
rect 138657 199746 138723 199749
rect 138124 199744 138723 199746
rect 138124 199688 138662 199744
rect 138718 199688 138723 199744
rect 138124 199686 138723 199688
rect 138124 199684 138130 199686
rect 138657 199683 138723 199686
rect 138982 199613 139042 199853
rect 139158 199820 139164 199884
rect 139228 199882 139234 199884
rect 139350 199882 139410 199956
rect 152598 199919 152658 200094
rect 166206 200092 166212 200156
rect 166276 200154 166282 200156
rect 166276 200094 171242 200154
rect 166276 200092 166282 200094
rect 161062 200018 161306 200052
rect 161062 199992 162456 200018
rect 161062 199919 161122 199992
rect 161246 199958 162456 199992
rect 139807 199916 139873 199919
rect 140175 199916 140241 199919
rect 139764 199914 139873 199916
rect 139764 199882 139812 199914
rect 139228 199822 139286 199882
rect 139350 199858 139812 199882
rect 139868 199858 139873 199914
rect 139350 199853 139873 199858
rect 140040 199914 140241 199916
rect 140040 199858 140180 199914
rect 140236 199858 140241 199914
rect 140040 199856 140241 199858
rect 139350 199822 139824 199853
rect 139228 199820 139234 199822
rect 139393 199746 139459 199749
rect 139258 199744 139459 199746
rect 139258 199688 139398 199744
rect 139454 199688 139459 199744
rect 139258 199686 139459 199688
rect 140040 199746 140100 199856
rect 140175 199853 140241 199856
rect 140451 199914 140517 199919
rect 140451 199858 140456 199914
rect 140512 199858 140517 199914
rect 140635 199914 140701 199919
rect 140635 199884 140640 199914
rect 140696 199884 140701 199914
rect 140911 199916 140977 199919
rect 141463 199918 141529 199919
rect 141458 199916 141464 199918
rect 140911 199914 141250 199916
rect 140451 199853 140517 199858
rect 140454 199749 140514 199853
rect 140630 199820 140636 199884
rect 140700 199882 140706 199884
rect 140700 199822 140758 199882
rect 140911 199858 140916 199914
rect 140972 199858 141250 199914
rect 140911 199856 141250 199858
rect 141372 199856 141464 199916
rect 140911 199853 140977 199856
rect 140700 199820 140706 199822
rect 140221 199746 140287 199749
rect 140040 199744 140287 199746
rect 140040 199688 140226 199744
rect 140282 199688 140287 199744
rect 140040 199686 140287 199688
rect 137645 199608 137754 199613
rect 137645 199552 137650 199608
rect 137706 199552 137754 199608
rect 137645 199550 137754 199552
rect 137645 199547 137711 199550
rect 137870 199548 137876 199612
rect 137940 199610 137946 199612
rect 138105 199610 138171 199613
rect 137940 199608 138171 199610
rect 137940 199552 138110 199608
rect 138166 199552 138171 199608
rect 137940 199550 138171 199552
rect 138982 199608 139091 199613
rect 138982 199552 139030 199608
rect 139086 199552 139091 199608
rect 138982 199550 139091 199552
rect 137940 199548 137946 199550
rect 138105 199547 138171 199550
rect 139025 199547 139091 199550
rect 139258 199474 139318 199686
rect 139393 199683 139459 199686
rect 140221 199683 140287 199686
rect 140405 199744 140514 199749
rect 140405 199688 140410 199744
rect 140466 199688 140514 199744
rect 140405 199686 140514 199688
rect 141190 199746 141250 199856
rect 141458 199854 141464 199856
rect 141528 199854 141534 199918
rect 141647 199916 141713 199919
rect 141647 199914 141986 199916
rect 141647 199858 141652 199914
rect 141708 199884 141986 199914
rect 142659 199914 142725 199919
rect 141708 199858 141924 199884
rect 141647 199856 141924 199858
rect 141463 199853 141529 199854
rect 141647 199853 141713 199856
rect 141918 199820 141924 199856
rect 141988 199820 141994 199884
rect 142102 199820 142108 199884
rect 142172 199882 142178 199884
rect 142659 199882 142664 199914
rect 142172 199858 142664 199882
rect 142720 199858 142725 199914
rect 142843 199914 142909 199919
rect 142843 199884 142848 199914
rect 142904 199884 142909 199914
rect 143027 199914 143093 199919
rect 143855 199916 143921 199919
rect 144407 199916 144473 199919
rect 142172 199853 142725 199858
rect 142172 199822 142722 199853
rect 142172 199820 142178 199822
rect 142838 199820 142844 199884
rect 142908 199882 142914 199884
rect 142908 199822 142966 199882
rect 143027 199858 143032 199914
rect 143088 199882 143093 199914
rect 143812 199914 143921 199916
rect 143206 199882 143212 199884
rect 143088 199858 143212 199882
rect 143027 199853 143212 199858
rect 143030 199822 143212 199853
rect 142908 199820 142914 199822
rect 143206 199820 143212 199822
rect 143276 199820 143282 199884
rect 143812 199858 143860 199914
rect 143916 199858 143921 199914
rect 144180 199914 144473 199916
rect 144180 199884 144412 199914
rect 143812 199853 143921 199858
rect 142061 199746 142127 199749
rect 141190 199744 142127 199746
rect 141190 199688 142066 199744
rect 142122 199688 142127 199744
rect 141190 199686 142127 199688
rect 140405 199683 140471 199686
rect 142061 199683 142127 199686
rect 142245 199746 142311 199749
rect 142654 199746 142660 199748
rect 142245 199744 142660 199746
rect 142245 199688 142250 199744
rect 142306 199688 142660 199744
rect 142245 199686 142660 199688
rect 142245 199683 142311 199686
rect 142654 199684 142660 199686
rect 142724 199684 142730 199748
rect 143812 199746 143872 199853
rect 144126 199820 144132 199884
rect 144196 199858 144412 199884
rect 144468 199858 144473 199914
rect 144196 199856 144473 199858
rect 144196 199822 144240 199856
rect 144407 199853 144473 199856
rect 144683 199914 144749 199919
rect 144683 199858 144688 199914
rect 144744 199858 144749 199914
rect 145419 199914 145485 199919
rect 145879 199916 145945 199919
rect 145419 199884 145424 199914
rect 145480 199884 145485 199914
rect 145744 199914 145945 199916
rect 144683 199853 144749 199858
rect 144196 199820 144202 199822
rect 142846 199686 143872 199746
rect 139393 199610 139459 199613
rect 142846 199610 142906 199686
rect 139393 199608 142906 199610
rect 139393 199552 139398 199608
rect 139454 199552 142906 199608
rect 139393 199550 142906 199552
rect 143349 199610 143415 199613
rect 144686 199610 144746 199853
rect 145414 199820 145420 199884
rect 145484 199882 145490 199884
rect 145484 199822 145542 199882
rect 145744 199858 145884 199914
rect 145940 199858 145945 199914
rect 145744 199856 145945 199858
rect 145484 199820 145490 199822
rect 145744 199749 145804 199856
rect 145879 199853 145945 199856
rect 146063 199916 146129 199919
rect 146063 199914 146402 199916
rect 146063 199858 146068 199914
rect 146124 199858 146402 199914
rect 146523 199914 146589 199919
rect 146523 199884 146528 199914
rect 146584 199884 146589 199914
rect 146891 199914 146957 199919
rect 146063 199856 146402 199858
rect 146063 199853 146129 199856
rect 145005 199748 145071 199749
rect 145005 199746 145052 199748
rect 144960 199744 145052 199746
rect 144960 199688 145010 199744
rect 144960 199686 145052 199688
rect 145005 199684 145052 199686
rect 145116 199684 145122 199748
rect 145741 199744 145807 199749
rect 145741 199688 145746 199744
rect 145802 199688 145807 199744
rect 145005 199683 145071 199684
rect 145741 199683 145807 199688
rect 143349 199608 144746 199610
rect 143349 199552 143354 199608
rect 143410 199552 144746 199608
rect 143349 199550 144746 199552
rect 146342 199610 146402 199856
rect 146518 199820 146524 199884
rect 146588 199882 146594 199884
rect 146588 199822 146646 199882
rect 146891 199858 146896 199914
rect 146952 199858 146957 199914
rect 147259 199914 147325 199919
rect 147259 199884 147264 199914
rect 147320 199884 147325 199914
rect 150571 199914 150637 199919
rect 146891 199853 146957 199858
rect 146588 199820 146594 199822
rect 146569 199748 146635 199749
rect 146518 199684 146524 199748
rect 146588 199746 146635 199748
rect 146588 199744 146680 199746
rect 146630 199688 146680 199744
rect 146588 199686 146680 199688
rect 146588 199684 146635 199686
rect 146569 199683 146635 199684
rect 146477 199610 146543 199613
rect 146342 199608 146543 199610
rect 146342 199552 146482 199608
rect 146538 199552 146543 199608
rect 146342 199550 146543 199552
rect 139393 199547 139459 199550
rect 143349 199547 143415 199550
rect 146477 199547 146543 199550
rect 139577 199474 139643 199477
rect 139258 199472 139643 199474
rect 139258 199416 139582 199472
rect 139638 199416 139643 199472
rect 139258 199414 139643 199416
rect 139577 199411 139643 199414
rect 141601 199474 141667 199477
rect 143717 199474 143783 199477
rect 141601 199472 143783 199474
rect 141601 199416 141606 199472
rect 141662 199416 143722 199472
rect 143778 199416 143783 199472
rect 141601 199414 143783 199416
rect 141601 199411 141667 199414
rect 143717 199411 143783 199414
rect 144177 199474 144243 199477
rect 146569 199474 146635 199477
rect 144177 199472 146635 199474
rect 144177 199416 144182 199472
rect 144238 199416 146574 199472
rect 146630 199416 146635 199472
rect 144177 199414 146635 199416
rect 146894 199474 146954 199853
rect 147254 199820 147260 199884
rect 147324 199882 147330 199884
rect 147324 199822 147382 199882
rect 147324 199820 147330 199822
rect 148174 199820 148180 199884
rect 148244 199882 148250 199884
rect 150571 199882 150576 199914
rect 148244 199858 150576 199882
rect 150632 199858 150637 199914
rect 148244 199853 150637 199858
rect 151491 199914 151557 199919
rect 151491 199858 151496 199914
rect 151552 199858 151557 199914
rect 151491 199853 151557 199858
rect 152595 199914 152661 199919
rect 153055 199916 153121 199919
rect 152595 199858 152600 199914
rect 152656 199858 152661 199914
rect 153012 199914 153121 199916
rect 152595 199853 152661 199858
rect 148244 199822 150634 199853
rect 148244 199820 148250 199822
rect 151494 199749 151554 199853
rect 152774 199820 152780 199884
rect 152844 199882 152850 199884
rect 153012 199882 153060 199914
rect 152844 199858 153060 199882
rect 153116 199858 153121 199914
rect 152844 199853 153121 199858
rect 153423 199916 153489 199919
rect 153423 199914 153624 199916
rect 153423 199858 153428 199914
rect 153484 199858 153624 199914
rect 153423 199856 153624 199858
rect 153423 199853 153489 199856
rect 152844 199822 153072 199853
rect 152844 199820 152850 199822
rect 147581 199748 147647 199749
rect 147581 199744 147628 199748
rect 147692 199746 147698 199748
rect 147581 199688 147586 199744
rect 147581 199684 147628 199688
rect 147692 199686 147738 199746
rect 147692 199684 147698 199686
rect 147806 199684 147812 199748
rect 147876 199746 147882 199748
rect 148639 199746 148705 199749
rect 148869 199748 148935 199749
rect 148869 199746 148916 199748
rect 147876 199744 148705 199746
rect 147876 199688 148644 199744
rect 148700 199688 148705 199744
rect 147876 199686 148705 199688
rect 148824 199744 148916 199746
rect 148824 199688 148874 199744
rect 148824 199686 148916 199688
rect 147876 199684 147882 199686
rect 147581 199683 147647 199684
rect 148639 199683 148705 199686
rect 148869 199684 148916 199686
rect 148980 199684 148986 199748
rect 150433 199746 150499 199749
rect 149286 199744 150499 199746
rect 149286 199688 150438 199744
rect 150494 199688 150499 199744
rect 149286 199686 150499 199688
rect 148869 199683 148935 199684
rect 147121 199474 147187 199477
rect 146894 199472 147187 199474
rect 146894 199416 147126 199472
rect 147182 199416 147187 199472
rect 146894 199414 147187 199416
rect 144177 199411 144243 199414
rect 146569 199411 146635 199414
rect 147121 199411 147187 199414
rect 147857 199474 147923 199477
rect 149286 199474 149346 199686
rect 150433 199683 150499 199686
rect 151445 199744 151554 199749
rect 151445 199688 151450 199744
rect 151506 199688 151554 199744
rect 151445 199686 151554 199688
rect 151445 199683 151511 199686
rect 147857 199472 149346 199474
rect 147857 199416 147862 199472
rect 147918 199416 149346 199472
rect 147857 199414 149346 199416
rect 153564 199474 153624 199856
rect 153883 199914 153949 199919
rect 153883 199858 153888 199914
rect 153944 199858 153949 199914
rect 153883 199853 153949 199858
rect 154343 199916 154409 199919
rect 154343 199914 154682 199916
rect 154343 199858 154348 199914
rect 154404 199858 154682 199914
rect 154343 199856 154682 199858
rect 154343 199853 154409 199856
rect 153886 199746 153946 199853
rect 154113 199746 154179 199749
rect 153886 199744 154179 199746
rect 153886 199688 154118 199744
rect 154174 199688 154179 199744
rect 153886 199686 154179 199688
rect 154113 199683 154179 199686
rect 154297 199746 154363 199749
rect 154622 199746 154682 199856
rect 154803 199914 154869 199919
rect 154803 199858 154808 199914
rect 154864 199858 154869 199914
rect 154803 199853 154869 199858
rect 155079 199914 155145 199919
rect 155079 199858 155084 199914
rect 155140 199858 155145 199914
rect 155079 199853 155145 199858
rect 156091 199914 156157 199919
rect 157103 199916 157169 199919
rect 156091 199858 156096 199914
rect 156152 199858 156157 199914
rect 156922 199914 157169 199916
rect 156922 199882 157108 199914
rect 156091 199853 156157 199858
rect 156876 199858 157108 199882
rect 157164 199858 157169 199914
rect 156876 199856 157169 199858
rect 154806 199749 154866 199853
rect 154297 199744 154682 199746
rect 154297 199688 154302 199744
rect 154358 199688 154682 199744
rect 154297 199686 154682 199688
rect 154757 199744 154866 199749
rect 154757 199688 154762 199744
rect 154818 199688 154866 199744
rect 154757 199686 154866 199688
rect 154297 199683 154363 199686
rect 154757 199683 154823 199686
rect 155082 199610 155142 199853
rect 156094 199749 156154 199853
rect 156045 199744 156154 199749
rect 156045 199688 156050 199744
rect 156106 199688 156154 199744
rect 156045 199686 156154 199688
rect 156876 199822 156982 199856
rect 157103 199853 157169 199856
rect 157747 199914 157813 199919
rect 157747 199858 157752 199914
rect 157808 199858 157813 199914
rect 157747 199853 157813 199858
rect 158023 199916 158089 199919
rect 158023 199914 158224 199916
rect 158023 199858 158028 199914
rect 158084 199858 158224 199914
rect 158299 199914 158365 199919
rect 158299 199884 158304 199914
rect 158360 199884 158365 199914
rect 158667 199914 158733 199919
rect 158667 199884 158672 199914
rect 158728 199884 158733 199914
rect 159311 199914 159377 199919
rect 158023 199856 158224 199858
rect 158023 199853 158089 199856
rect 156045 199683 156111 199686
rect 156321 199610 156387 199613
rect 155082 199608 156387 199610
rect 155082 199552 156326 199608
rect 156382 199552 156387 199608
rect 155082 199550 156387 199552
rect 156876 199610 156936 199822
rect 157011 199748 157077 199749
rect 157006 199684 157012 199748
rect 157076 199746 157082 199748
rect 157076 199686 157168 199746
rect 157076 199684 157082 199686
rect 157011 199683 157077 199684
rect 157750 199613 157810 199853
rect 157977 199746 158043 199749
rect 158164 199746 158224 199856
rect 158294 199820 158300 199884
rect 158364 199882 158370 199884
rect 158364 199822 158422 199882
rect 158364 199820 158370 199822
rect 158662 199820 158668 199884
rect 158732 199882 158738 199884
rect 158732 199822 158790 199882
rect 159311 199858 159316 199914
rect 159372 199858 159377 199914
rect 159311 199853 159377 199858
rect 160047 199914 160113 199919
rect 160047 199858 160052 199914
rect 160108 199858 160113 199914
rect 160047 199853 160113 199858
rect 160415 199916 160481 199919
rect 160415 199914 160616 199916
rect 160415 199858 160420 199914
rect 160476 199882 160616 199914
rect 161059 199914 161125 199919
rect 160870 199882 160876 199884
rect 160476 199858 160876 199882
rect 160415 199856 160876 199858
rect 160415 199853 160481 199856
rect 158732 199820 158738 199822
rect 157977 199744 158224 199746
rect 157977 199688 157982 199744
rect 158038 199688 158224 199744
rect 157977 199686 158224 199688
rect 158391 199746 158457 199749
rect 159081 199746 159147 199749
rect 159314 199746 159374 199853
rect 158391 199744 158730 199746
rect 158391 199688 158396 199744
rect 158452 199688 158730 199744
rect 158391 199686 158730 199688
rect 157977 199683 158043 199686
rect 158391 199683 158457 199686
rect 157057 199610 157123 199613
rect 156876 199608 157123 199610
rect 156876 199552 157062 199608
rect 157118 199552 157123 199608
rect 156876 199550 157123 199552
rect 157750 199608 157859 199613
rect 157750 199552 157798 199608
rect 157854 199552 157859 199608
rect 157750 199550 157859 199552
rect 158670 199610 158730 199686
rect 159081 199744 159374 199746
rect 159081 199688 159086 199744
rect 159142 199688 159374 199744
rect 159081 199686 159374 199688
rect 159081 199683 159147 199686
rect 158805 199610 158871 199613
rect 158670 199608 158871 199610
rect 158670 199552 158810 199608
rect 158866 199552 158871 199608
rect 158670 199550 158871 199552
rect 160050 199610 160110 199853
rect 160556 199822 160876 199856
rect 160870 199820 160876 199822
rect 160940 199820 160946 199884
rect 161059 199858 161064 199914
rect 161120 199858 161125 199914
rect 161243 199884 161309 199885
rect 161059 199853 161125 199858
rect 161238 199820 161244 199884
rect 161308 199882 161314 199884
rect 161308 199822 161400 199882
rect 162163 199880 162229 199885
rect 162163 199824 162168 199880
rect 162224 199824 162229 199880
rect 161308 199820 161314 199822
rect 161243 199819 161309 199820
rect 162163 199819 162229 199824
rect 162166 199749 162226 199819
rect 161238 199684 161244 199748
rect 161308 199746 161314 199748
rect 161565 199746 161631 199749
rect 161308 199744 161631 199746
rect 161308 199688 161570 199744
rect 161626 199688 161631 199744
rect 161308 199686 161631 199688
rect 162166 199744 162275 199749
rect 162166 199688 162214 199744
rect 162270 199688 162275 199744
rect 162166 199686 162275 199688
rect 162396 199746 162456 199958
rect 171182 199919 171242 200094
rect 162715 199914 162781 199919
rect 162526 199820 162532 199884
rect 162596 199882 162602 199884
rect 162715 199882 162720 199914
rect 162596 199858 162720 199882
rect 162776 199858 162781 199914
rect 162596 199853 162781 199858
rect 163175 199914 163241 199919
rect 163175 199858 163180 199914
rect 163236 199858 163241 199914
rect 164739 199914 164805 199919
rect 163175 199853 163241 199858
rect 164003 199880 164069 199885
rect 164739 199884 164744 199914
rect 164800 199884 164805 199914
rect 165291 199914 165357 199919
rect 162596 199822 162778 199853
rect 162596 199820 162602 199822
rect 163178 199749 163238 199853
rect 164003 199824 164008 199880
rect 164064 199824 164069 199880
rect 164003 199819 164069 199824
rect 164734 199820 164740 199884
rect 164804 199882 164810 199884
rect 164804 199822 164862 199882
rect 164804 199820 164810 199822
rect 165102 199820 165108 199884
rect 165172 199882 165178 199884
rect 165291 199882 165296 199914
rect 165172 199858 165296 199882
rect 165352 199858 165357 199914
rect 165475 199914 165541 199919
rect 165475 199884 165480 199914
rect 165536 199884 165541 199914
rect 168235 199914 168301 199919
rect 165843 199884 165909 199885
rect 165172 199853 165357 199858
rect 165172 199822 165354 199853
rect 165172 199820 165178 199822
rect 165470 199820 165476 199884
rect 165540 199882 165546 199884
rect 165838 199882 165844 199884
rect 165540 199822 165598 199882
rect 165752 199822 165844 199882
rect 165540 199820 165546 199822
rect 165838 199820 165844 199822
rect 165908 199820 165914 199884
rect 166574 199820 166580 199884
rect 166644 199882 166650 199884
rect 166855 199882 166921 199885
rect 167959 199882 168025 199885
rect 166644 199880 166921 199882
rect 166644 199824 166860 199880
rect 166916 199824 166921 199880
rect 166644 199822 166921 199824
rect 166644 199820 166650 199822
rect 165843 199819 165909 199820
rect 166855 199819 166921 199822
rect 167732 199880 168025 199882
rect 167732 199824 167964 199880
rect 168020 199824 168025 199880
rect 168235 199858 168240 199914
rect 168296 199858 168301 199914
rect 168603 199914 168669 199919
rect 168603 199884 168608 199914
rect 168664 199884 168669 199914
rect 168879 199916 168945 199919
rect 168879 199914 168988 199916
rect 168235 199853 168301 199858
rect 167732 199822 168025 199824
rect 162577 199746 162643 199749
rect 162396 199744 162643 199746
rect 162396 199688 162582 199744
rect 162638 199688 162643 199744
rect 162396 199686 162643 199688
rect 161308 199684 161314 199686
rect 161565 199683 161631 199686
rect 162209 199683 162275 199686
rect 162577 199683 162643 199686
rect 163129 199744 163238 199749
rect 163129 199688 163134 199744
rect 163190 199688 163238 199744
rect 163129 199686 163238 199688
rect 164006 199746 164066 199819
rect 164141 199746 164207 199749
rect 164006 199744 164207 199746
rect 164006 199688 164146 199744
rect 164202 199688 164207 199744
rect 164006 199686 164207 199688
rect 163129 199683 163195 199686
rect 164141 199683 164207 199686
rect 165337 199746 165403 199749
rect 165470 199746 165476 199748
rect 165337 199744 165476 199746
rect 165337 199688 165342 199744
rect 165398 199688 165476 199744
rect 165337 199686 165476 199688
rect 165337 199683 165403 199686
rect 165470 199684 165476 199686
rect 165540 199684 165546 199748
rect 167732 199746 167792 199822
rect 167959 199819 168025 199822
rect 167913 199746 167979 199749
rect 167732 199744 167979 199746
rect 167732 199688 167918 199744
rect 167974 199688 167979 199744
rect 167732 199686 167979 199688
rect 167913 199683 167979 199686
rect 168238 199613 168298 199853
rect 168598 199820 168604 199884
rect 168668 199882 168674 199884
rect 168668 199822 168726 199882
rect 168879 199858 168884 199914
rect 168940 199858 168988 199914
rect 169155 199914 169221 199919
rect 169155 199884 169160 199914
rect 169216 199884 169221 199914
rect 169431 199914 169497 199919
rect 168879 199853 168988 199858
rect 168668 199820 168674 199822
rect 168928 199749 168988 199853
rect 169150 199820 169156 199884
rect 169220 199882 169226 199884
rect 169220 199822 169278 199882
rect 169431 199858 169436 199914
rect 169492 199882 169497 199914
rect 170075 199914 170141 199919
rect 170535 199916 170601 199919
rect 169886 199882 169892 199884
rect 169492 199858 169892 199882
rect 169431 199853 169892 199858
rect 169434 199822 169892 199853
rect 169220 199820 169226 199822
rect 169886 199820 169892 199822
rect 169956 199820 169962 199884
rect 170075 199858 170080 199914
rect 170136 199858 170141 199914
rect 170075 199853 170141 199858
rect 170492 199914 170601 199916
rect 170492 199858 170540 199914
rect 170596 199858 170601 199914
rect 170995 199914 171061 199919
rect 170995 199884 171000 199914
rect 171056 199884 171061 199914
rect 171179 199914 171245 199919
rect 170492 199853 170601 199858
rect 168649 199744 168715 199749
rect 168649 199688 168654 199744
rect 168710 199688 168715 199744
rect 168649 199683 168715 199688
rect 168925 199744 168991 199749
rect 168925 199688 168930 199744
rect 168986 199688 168991 199744
rect 168925 199683 168991 199688
rect 162301 199610 162367 199613
rect 160050 199608 162367 199610
rect 160050 199552 162306 199608
rect 162362 199552 162367 199608
rect 160050 199550 162367 199552
rect 156321 199547 156387 199550
rect 157057 199547 157123 199550
rect 157793 199547 157859 199550
rect 158805 199547 158871 199550
rect 162301 199547 162367 199550
rect 163773 199612 163839 199613
rect 163773 199608 163820 199612
rect 163884 199610 163890 199612
rect 164417 199610 164483 199613
rect 165153 199610 165219 199613
rect 163773 199552 163778 199608
rect 163773 199548 163820 199552
rect 163884 199550 163930 199610
rect 164417 199608 165219 199610
rect 164417 199552 164422 199608
rect 164478 199552 165158 199608
rect 165214 199552 165219 199608
rect 164417 199550 165219 199552
rect 163884 199548 163890 199550
rect 163773 199547 163839 199548
rect 164417 199547 164483 199550
rect 165153 199547 165219 199550
rect 165889 199610 165955 199613
rect 166022 199610 166028 199612
rect 165889 199608 166028 199610
rect 165889 199552 165894 199608
rect 165950 199552 166028 199608
rect 165889 199550 166028 199552
rect 165889 199547 165955 199550
rect 166022 199548 166028 199550
rect 166092 199548 166098 199612
rect 166809 199610 166875 199613
rect 168046 199610 168052 199612
rect 166809 199608 168052 199610
rect 166809 199552 166814 199608
rect 166870 199552 168052 199608
rect 166809 199550 168052 199552
rect 166809 199547 166875 199550
rect 168046 199548 168052 199550
rect 168116 199548 168122 199612
rect 168189 199608 168298 199613
rect 168189 199552 168194 199608
rect 168250 199552 168298 199608
rect 168189 199550 168298 199552
rect 168652 199610 168712 199683
rect 169334 199610 169340 199612
rect 168652 199550 169340 199610
rect 168189 199547 168255 199550
rect 169334 199548 169340 199550
rect 169404 199548 169410 199612
rect 170078 199610 170138 199853
rect 170492 199746 170552 199853
rect 170990 199820 170996 199884
rect 171060 199882 171066 199884
rect 171060 199822 171118 199882
rect 171179 199858 171184 199914
rect 171240 199858 171245 199914
rect 171179 199853 171245 199858
rect 171639 199916 171705 199919
rect 172191 199916 172257 199919
rect 171639 199914 171748 199916
rect 171639 199858 171644 199914
rect 171700 199882 171748 199914
rect 172191 199914 172300 199916
rect 171910 199882 171916 199884
rect 171700 199858 171916 199882
rect 171639 199853 171916 199858
rect 171688 199822 171916 199853
rect 171060 199820 171066 199822
rect 171910 199820 171916 199822
rect 171980 199820 171986 199884
rect 172191 199858 172196 199914
rect 172252 199858 172300 199914
rect 172191 199853 172300 199858
rect 172375 199914 172441 199919
rect 172375 199858 172380 199914
rect 172436 199882 172441 199914
rect 173571 199914 173637 199919
rect 172646 199882 172652 199884
rect 172436 199858 172652 199882
rect 172375 199853 172652 199858
rect 172240 199746 172300 199853
rect 172378 199822 172652 199853
rect 172646 199820 172652 199822
rect 172716 199820 172722 199884
rect 172927 199882 172993 199885
rect 173571 199884 173576 199914
rect 173632 199884 173637 199914
rect 173755 199914 173821 199919
rect 172927 199880 173450 199882
rect 172927 199824 172932 199880
rect 172988 199824 173450 199880
rect 172927 199822 173450 199824
rect 172927 199819 172993 199822
rect 172421 199746 172487 199749
rect 170492 199686 171288 199746
rect 172240 199744 172487 199746
rect 172240 199688 172426 199744
rect 172482 199688 172487 199744
rect 172240 199686 172487 199688
rect 170949 199610 171015 199613
rect 170078 199608 171015 199610
rect 170078 199552 170954 199608
rect 171010 199552 171015 199608
rect 170078 199550 171015 199552
rect 171228 199610 171288 199686
rect 172421 199683 172487 199686
rect 172697 199746 172763 199749
rect 172697 199744 173036 199746
rect 172697 199688 172702 199744
rect 172758 199688 173036 199744
rect 172697 199686 173036 199688
rect 172697 199683 172763 199686
rect 172976 199613 173036 199686
rect 171542 199610 171548 199612
rect 171228 199550 171548 199610
rect 170949 199547 171015 199550
rect 171542 199548 171548 199550
rect 171612 199548 171618 199612
rect 172973 199608 173039 199613
rect 172973 199552 172978 199608
rect 173034 199552 173039 199608
rect 172973 199547 173039 199552
rect 173390 199610 173450 199822
rect 173566 199820 173572 199884
rect 173636 199882 173642 199884
rect 173636 199822 173694 199882
rect 173755 199858 173760 199914
rect 173816 199858 173821 199914
rect 173755 199853 173821 199858
rect 173636 199820 173642 199822
rect 173758 199748 173818 199853
rect 173988 199749 174048 200230
rect 207289 200227 207355 200230
rect 180517 200154 180583 200157
rect 174126 200152 180583 200154
rect 174126 200096 180522 200152
rect 180578 200096 180583 200152
rect 174126 200094 180583 200096
rect 174126 199919 174186 200094
rect 180517 200091 180583 200094
rect 187141 200154 187207 200157
rect 209957 200154 210023 200157
rect 187141 200152 210023 200154
rect 187141 200096 187146 200152
rect 187202 200096 209962 200152
rect 210018 200096 210023 200152
rect 187141 200094 210023 200096
rect 187141 200091 187207 200094
rect 209957 200091 210023 200094
rect 174123 199914 174189 199919
rect 174123 199858 174128 199914
rect 174184 199858 174189 199914
rect 174123 199853 174189 199858
rect 174307 199914 174373 199919
rect 174307 199858 174312 199914
rect 174368 199858 174373 199914
rect 174307 199853 174373 199858
rect 174675 199914 174741 199919
rect 175135 199916 175201 199919
rect 174675 199858 174680 199914
rect 174736 199858 174741 199914
rect 175092 199914 175201 199916
rect 174675 199853 174741 199858
rect 173750 199684 173756 199748
rect 173820 199684 173826 199748
rect 173985 199744 174051 199749
rect 173985 199688 173990 199744
rect 174046 199688 174051 199744
rect 173985 199683 174051 199688
rect 173801 199610 173867 199613
rect 173390 199608 173867 199610
rect 173390 199552 173806 199608
rect 173862 199552 173867 199608
rect 173390 199550 173867 199552
rect 174310 199610 174370 199853
rect 174678 199613 174738 199853
rect 174854 199820 174860 199884
rect 174924 199882 174930 199884
rect 175092 199882 175140 199914
rect 174924 199858 175140 199882
rect 175196 199858 175201 199914
rect 174924 199853 175201 199858
rect 175963 199914 176029 199919
rect 175963 199858 175968 199914
rect 176024 199858 176029 199914
rect 175963 199853 176029 199858
rect 176239 199916 176305 199919
rect 176239 199914 176348 199916
rect 176239 199858 176244 199914
rect 176300 199884 176348 199914
rect 176883 199914 176949 199919
rect 176300 199858 176332 199884
rect 176239 199853 176332 199858
rect 174924 199822 175152 199853
rect 174924 199820 174930 199822
rect 174445 199610 174511 199613
rect 174310 199608 174511 199610
rect 174310 199552 174450 199608
rect 174506 199552 174511 199608
rect 174310 199550 174511 199552
rect 173801 199547 173867 199550
rect 174445 199547 174511 199550
rect 174629 199608 174738 199613
rect 174629 199552 174634 199608
rect 174690 199552 174738 199608
rect 174629 199550 174738 199552
rect 175966 199610 176026 199853
rect 176288 199822 176332 199853
rect 176326 199820 176332 199822
rect 176396 199820 176402 199884
rect 176883 199858 176888 199914
rect 176944 199882 176949 199914
rect 179505 199882 179571 199885
rect 176944 199880 179571 199882
rect 176944 199858 179510 199880
rect 176883 199853 179510 199858
rect 176886 199824 179510 199853
rect 179566 199824 179571 199880
rect 176886 199822 179571 199824
rect 179505 199819 179571 199822
rect 180517 199610 180583 199613
rect 175966 199608 180583 199610
rect 175966 199552 180522 199608
rect 180578 199552 180583 199608
rect 175966 199550 180583 199552
rect 174629 199547 174695 199550
rect 180517 199547 180583 199550
rect 171358 199474 171364 199476
rect 153564 199414 171364 199474
rect 147857 199411 147923 199414
rect 171358 199412 171364 199414
rect 171428 199412 171434 199476
rect 171685 199474 171751 199477
rect 177849 199474 177915 199477
rect 171685 199472 177915 199474
rect 171685 199416 171690 199472
rect 171746 199416 177854 199472
rect 177910 199416 177915 199472
rect 171685 199414 177915 199416
rect 171685 199411 171751 199414
rect 177849 199411 177915 199414
rect 181345 199474 181411 199477
rect 181345 199472 186330 199474
rect 181345 199416 181350 199472
rect 181406 199416 186330 199472
rect 181345 199414 186330 199416
rect 181345 199411 181411 199414
rect 131849 199336 137202 199338
rect 131849 199280 131854 199336
rect 131910 199280 137202 199336
rect 131849 199278 137202 199280
rect 142153 199338 142219 199341
rect 147673 199338 147739 199341
rect 142153 199336 147739 199338
rect 142153 199280 142158 199336
rect 142214 199280 147678 199336
rect 147734 199280 147739 199336
rect 142153 199278 147739 199280
rect 103145 199275 103211 199278
rect 131849 199275 131915 199278
rect 142153 199275 142219 199278
rect 147673 199275 147739 199278
rect 155585 199338 155651 199341
rect 179597 199338 179663 199341
rect 155585 199336 179663 199338
rect 155585 199280 155590 199336
rect 155646 199280 179602 199336
rect 179658 199280 179663 199336
rect 155585 199278 179663 199280
rect 186270 199338 186330 199414
rect 203006 199338 203012 199340
rect 186270 199278 203012 199338
rect 155585 199275 155651 199278
rect 179597 199275 179663 199278
rect 203006 199276 203012 199278
rect 203076 199276 203082 199340
rect 99281 199202 99347 199205
rect 142153 199202 142219 199205
rect 99281 199200 142219 199202
rect 99281 199144 99286 199200
rect 99342 199144 142158 199200
rect 142214 199144 142219 199200
rect 99281 199142 142219 199144
rect 99281 199139 99347 199142
rect 142153 199139 142219 199142
rect 143625 199202 143691 199205
rect 144913 199202 144979 199205
rect 145373 199204 145439 199205
rect 145046 199202 145052 199204
rect 143625 199200 143826 199202
rect 143625 199144 143630 199200
rect 143686 199144 143826 199200
rect 143625 199142 143826 199144
rect 143625 199139 143691 199142
rect 122097 199066 122163 199069
rect 143625 199066 143691 199069
rect 122097 199064 143691 199066
rect 122097 199008 122102 199064
rect 122158 199008 143630 199064
rect 143686 199008 143691 199064
rect 122097 199006 143691 199008
rect 122097 199003 122163 199006
rect 143625 199003 143691 199006
rect 132217 198930 132283 198933
rect 136817 198930 136883 198933
rect 132217 198928 136883 198930
rect 132217 198872 132222 198928
rect 132278 198872 136822 198928
rect 136878 198872 136883 198928
rect 132217 198870 136883 198872
rect 132217 198867 132283 198870
rect 136817 198867 136883 198870
rect 138013 198930 138079 198933
rect 138422 198930 138428 198932
rect 138013 198928 138428 198930
rect 138013 198872 138018 198928
rect 138074 198872 138428 198928
rect 138013 198870 138428 198872
rect 138013 198867 138079 198870
rect 138422 198868 138428 198870
rect 138492 198868 138498 198932
rect 138841 198930 138907 198933
rect 143766 198930 143826 199142
rect 144913 199200 145052 199202
rect 144913 199144 144918 199200
rect 144974 199144 145052 199200
rect 144913 199142 145052 199144
rect 144913 199139 144979 199142
rect 145046 199140 145052 199142
rect 145116 199140 145122 199204
rect 145373 199202 145420 199204
rect 145328 199200 145420 199202
rect 145328 199144 145378 199200
rect 145328 199142 145420 199144
rect 145373 199140 145420 199142
rect 145484 199140 145490 199204
rect 146109 199202 146175 199205
rect 146334 199202 146340 199204
rect 146109 199200 146340 199202
rect 146109 199144 146114 199200
rect 146170 199144 146340 199200
rect 146109 199142 146340 199144
rect 145373 199139 145439 199140
rect 146109 199139 146175 199142
rect 146334 199140 146340 199142
rect 146404 199140 146410 199204
rect 164601 199202 164667 199205
rect 166809 199202 166875 199205
rect 164601 199200 166875 199202
rect 164601 199144 164606 199200
rect 164662 199144 166814 199200
rect 166870 199144 166875 199200
rect 164601 199142 166875 199144
rect 164601 199139 164667 199142
rect 166809 199139 166875 199142
rect 168598 199140 168604 199204
rect 168668 199202 168674 199204
rect 171685 199202 171751 199205
rect 173709 199204 173775 199205
rect 173709 199202 173756 199204
rect 168668 199200 171751 199202
rect 168668 199144 171690 199200
rect 171746 199144 171751 199200
rect 168668 199142 171751 199144
rect 173664 199200 173756 199202
rect 173664 199144 173714 199200
rect 173664 199142 173756 199144
rect 168668 199140 168674 199142
rect 171685 199139 171751 199142
rect 173709 199140 173756 199142
rect 173820 199140 173826 199204
rect 174353 199202 174419 199205
rect 200798 199202 200804 199204
rect 174353 199200 200804 199202
rect 174353 199144 174358 199200
rect 174414 199144 200804 199200
rect 174353 199142 200804 199144
rect 173709 199139 173775 199140
rect 174353 199139 174419 199142
rect 200798 199140 200804 199142
rect 200868 199140 200874 199204
rect 160093 199066 160159 199069
rect 167545 199066 167611 199069
rect 160093 199064 167611 199066
rect 160093 199008 160098 199064
rect 160154 199008 167550 199064
rect 167606 199008 167611 199064
rect 160093 199006 167611 199008
rect 160093 199003 160159 199006
rect 167545 199003 167611 199006
rect 175549 199066 175615 199069
rect 205030 199066 205036 199068
rect 175549 199064 205036 199066
rect 175549 199008 175554 199064
rect 175610 199008 205036 199064
rect 175549 199006 205036 199008
rect 175549 199003 175615 199006
rect 205030 199004 205036 199006
rect 205100 199004 205106 199068
rect 138841 198928 143826 198930
rect 138841 198872 138846 198928
rect 138902 198872 143826 198928
rect 138841 198870 143826 198872
rect 138841 198867 138907 198870
rect 144310 198868 144316 198932
rect 144380 198930 144386 198932
rect 144545 198930 144611 198933
rect 144380 198928 144611 198930
rect 144380 198872 144550 198928
rect 144606 198872 144611 198928
rect 144380 198870 144611 198872
rect 144380 198868 144386 198870
rect 144545 198867 144611 198870
rect 163313 198930 163379 198933
rect 169109 198930 169175 198933
rect 163313 198928 169175 198930
rect 163313 198872 163318 198928
rect 163374 198872 169114 198928
rect 169170 198872 169175 198928
rect 163313 198870 169175 198872
rect 163313 198867 163379 198870
rect 169109 198867 169175 198870
rect 175825 198930 175891 198933
rect 205214 198930 205220 198932
rect 175825 198928 205220 198930
rect 175825 198872 175830 198928
rect 175886 198872 205220 198928
rect 175825 198870 205220 198872
rect 175825 198867 175891 198870
rect 205214 198868 205220 198870
rect 205284 198868 205290 198932
rect 129181 198794 129247 198797
rect 152365 198794 152431 198797
rect 129181 198792 152431 198794
rect 129181 198736 129186 198792
rect 129242 198736 152370 198792
rect 152426 198736 152431 198792
rect 129181 198734 152431 198736
rect 129181 198731 129247 198734
rect 152365 198731 152431 198734
rect 160921 198794 160987 198797
rect 176009 198794 176075 198797
rect 217317 198794 217383 198797
rect 160921 198792 173266 198794
rect 160921 198736 160926 198792
rect 160982 198736 173266 198792
rect 160921 198734 173266 198736
rect 160921 198731 160987 198734
rect 138473 198658 138539 198661
rect 139158 198658 139164 198660
rect 138473 198656 139164 198658
rect 138473 198600 138478 198656
rect 138534 198600 139164 198656
rect 138473 198598 139164 198600
rect 138473 198595 138539 198598
rect 139158 198596 139164 198598
rect 139228 198596 139234 198660
rect 145741 198658 145807 198661
rect 146518 198658 146524 198660
rect 145741 198656 146524 198658
rect 145741 198600 145746 198656
rect 145802 198600 146524 198656
rect 145741 198598 146524 198600
rect 145741 198595 145807 198598
rect 146518 198596 146524 198598
rect 146588 198596 146594 198660
rect 160686 198596 160692 198660
rect 160756 198658 160762 198660
rect 166993 198658 167059 198661
rect 160756 198656 167059 198658
rect 160756 198600 166998 198656
rect 167054 198600 167059 198656
rect 160756 198598 167059 198600
rect 160756 198596 160762 198598
rect 166993 198595 167059 198598
rect 167729 198658 167795 198661
rect 169201 198660 169267 198661
rect 167862 198658 167868 198660
rect 167729 198656 167868 198658
rect 167729 198600 167734 198656
rect 167790 198600 167868 198656
rect 167729 198598 167868 198600
rect 167729 198595 167795 198598
rect 167862 198596 167868 198598
rect 167932 198596 167938 198660
rect 169150 198596 169156 198660
rect 169220 198658 169267 198660
rect 169385 198658 169451 198661
rect 169518 198658 169524 198660
rect 169220 198656 169312 198658
rect 169262 198600 169312 198656
rect 169220 198598 169312 198600
rect 169385 198656 169524 198658
rect 169385 198600 169390 198656
rect 169446 198600 169524 198656
rect 169385 198598 169524 198600
rect 169220 198596 169267 198598
rect 169201 198595 169267 198596
rect 169385 198595 169451 198598
rect 169518 198596 169524 198598
rect 169588 198596 169594 198660
rect 173206 198658 173266 198734
rect 176009 198792 217383 198794
rect 176009 198736 176014 198792
rect 176070 198736 217322 198792
rect 217378 198736 217383 198792
rect 176009 198734 217383 198736
rect 176009 198731 176075 198734
rect 217317 198731 217383 198734
rect 177665 198658 177731 198661
rect 173206 198656 177731 198658
rect 173206 198600 177670 198656
rect 177726 198600 177731 198656
rect 173206 198598 177731 198600
rect 177665 198595 177731 198598
rect 124070 198460 124076 198524
rect 124140 198522 124146 198524
rect 148133 198522 148199 198525
rect 124140 198520 148199 198522
rect 124140 198464 148138 198520
rect 148194 198464 148199 198520
rect 124140 198462 148199 198464
rect 124140 198460 124146 198462
rect 148133 198459 148199 198462
rect 150014 198460 150020 198524
rect 150084 198522 150090 198524
rect 162025 198522 162091 198525
rect 150084 198520 162091 198522
rect 150084 198464 162030 198520
rect 162086 198464 162091 198520
rect 150084 198462 162091 198464
rect 150084 198460 150090 198462
rect 162025 198459 162091 198462
rect 171910 198460 171916 198524
rect 171980 198522 171986 198524
rect 174997 198522 175063 198525
rect 171980 198520 175063 198522
rect 171980 198464 175002 198520
rect 175058 198464 175063 198520
rect 171980 198462 175063 198464
rect 171980 198460 171986 198462
rect 174997 198459 175063 198462
rect 176837 198522 176903 198525
rect 201534 198522 201540 198524
rect 176837 198520 201540 198522
rect 176837 198464 176842 198520
rect 176898 198464 201540 198520
rect 176837 198462 201540 198464
rect 176837 198459 176903 198462
rect 201534 198460 201540 198462
rect 201604 198460 201610 198524
rect 106038 198324 106044 198388
rect 106108 198386 106114 198388
rect 132401 198386 132467 198389
rect 136449 198388 136515 198389
rect 106108 198384 132467 198386
rect 106108 198328 132406 198384
rect 132462 198328 132467 198384
rect 106108 198326 132467 198328
rect 106108 198324 106114 198326
rect 132401 198323 132467 198326
rect 136398 198324 136404 198388
rect 136468 198386 136515 198388
rect 138565 198386 138631 198389
rect 149329 198386 149395 198389
rect 136468 198384 136560 198386
rect 136510 198328 136560 198384
rect 136468 198326 136560 198328
rect 138565 198384 149395 198386
rect 138565 198328 138570 198384
rect 138626 198328 149334 198384
rect 149390 198328 149395 198384
rect 138565 198326 149395 198328
rect 136468 198324 136515 198326
rect 136449 198323 136515 198324
rect 138565 198323 138631 198326
rect 149329 198323 149395 198326
rect 151486 198324 151492 198388
rect 151556 198386 151562 198388
rect 159081 198386 159147 198389
rect 151556 198384 159147 198386
rect 151556 198328 159086 198384
rect 159142 198328 159147 198384
rect 151556 198326 159147 198328
rect 151556 198324 151562 198326
rect 159081 198323 159147 198326
rect 173566 198324 173572 198388
rect 173636 198386 173642 198388
rect 212533 198386 212599 198389
rect 173636 198384 212599 198386
rect 173636 198328 212538 198384
rect 212594 198328 212599 198384
rect 173636 198326 212599 198328
rect 173636 198324 173642 198326
rect 212533 198323 212599 198326
rect 107510 198188 107516 198252
rect 107580 198250 107586 198252
rect 127157 198250 127223 198253
rect 107580 198248 127223 198250
rect 107580 198192 127162 198248
rect 127218 198192 127223 198248
rect 107580 198190 127223 198192
rect 107580 198188 107586 198190
rect 127157 198187 127223 198190
rect 141693 198250 141759 198253
rect 141918 198250 141924 198252
rect 141693 198248 141924 198250
rect 141693 198192 141698 198248
rect 141754 198192 141924 198248
rect 141693 198190 141924 198192
rect 141693 198187 141759 198190
rect 141918 198188 141924 198190
rect 141988 198188 141994 198252
rect 172053 198250 172119 198253
rect 213913 198250 213979 198253
rect 172053 198248 213979 198250
rect 172053 198192 172058 198248
rect 172114 198192 213918 198248
rect 213974 198192 213979 198248
rect 172053 198190 213979 198192
rect 172053 198187 172119 198190
rect 213913 198187 213979 198190
rect 107326 198052 107332 198116
rect 107396 198114 107402 198116
rect 129273 198114 129339 198117
rect 107396 198112 129339 198114
rect 107396 198056 129278 198112
rect 129334 198056 129339 198112
rect 107396 198054 129339 198056
rect 107396 198052 107402 198054
rect 129273 198051 129339 198054
rect 148174 198052 148180 198116
rect 148244 198114 148250 198116
rect 150893 198114 150959 198117
rect 148244 198112 150959 198114
rect 148244 198056 150898 198112
rect 150954 198056 150959 198112
rect 148244 198054 150959 198056
rect 148244 198052 148250 198054
rect 150893 198051 150959 198054
rect 156873 198114 156939 198117
rect 157190 198114 157196 198116
rect 156873 198112 157196 198114
rect 156873 198056 156878 198112
rect 156934 198056 157196 198112
rect 156873 198054 157196 198056
rect 156873 198051 156939 198054
rect 157190 198052 157196 198054
rect 157260 198052 157266 198116
rect 171133 198114 171199 198117
rect 214005 198114 214071 198117
rect 171133 198112 214071 198114
rect 171133 198056 171138 198112
rect 171194 198056 214010 198112
rect 214066 198056 214071 198112
rect 171133 198054 214071 198056
rect 171133 198051 171199 198054
rect 214005 198051 214071 198054
rect 102910 197916 102916 197980
rect 102980 197978 102986 197980
rect 102980 197918 118710 197978
rect 102980 197916 102986 197918
rect 118650 197842 118710 197918
rect 147438 197916 147444 197980
rect 147508 197978 147514 197980
rect 160001 197978 160067 197981
rect 147508 197976 160067 197978
rect 147508 197920 160006 197976
rect 160062 197920 160067 197976
rect 147508 197918 160067 197920
rect 147508 197916 147514 197918
rect 160001 197915 160067 197918
rect 171542 197916 171548 197980
rect 171612 197978 171618 197980
rect 214189 197978 214255 197981
rect 171612 197976 214255 197978
rect 171612 197920 214194 197976
rect 214250 197920 214255 197976
rect 171612 197918 214255 197920
rect 171612 197916 171618 197918
rect 214189 197915 214255 197918
rect 134190 197842 134196 197844
rect 118650 197782 134196 197842
rect 134190 197780 134196 197782
rect 134260 197780 134266 197844
rect 178401 197842 178467 197845
rect 202822 197842 202828 197844
rect 178401 197840 202828 197842
rect 178401 197784 178406 197840
rect 178462 197784 202828 197840
rect 178401 197782 202828 197784
rect 178401 197779 178467 197782
rect 202822 197780 202828 197782
rect 202892 197780 202898 197844
rect 164734 197644 164740 197708
rect 164804 197706 164810 197708
rect 168741 197706 168807 197709
rect 164804 197704 168807 197706
rect 164804 197648 168746 197704
rect 168802 197648 168807 197704
rect 164804 197646 168807 197648
rect 164804 197644 164810 197646
rect 168741 197643 168807 197646
rect 172421 197570 172487 197573
rect 172421 197568 178050 197570
rect 172421 197512 172426 197568
rect 172482 197512 178050 197568
rect 172421 197510 178050 197512
rect 172421 197507 172487 197510
rect 142797 197436 142863 197437
rect 142797 197434 142844 197436
rect 142752 197432 142844 197434
rect 142752 197376 142802 197432
rect 142752 197374 142844 197376
rect 142797 197372 142844 197374
rect 142908 197372 142914 197436
rect 142981 197434 143047 197437
rect 143206 197434 143212 197436
rect 142981 197432 143212 197434
rect 142981 197376 142986 197432
rect 143042 197376 143212 197432
rect 142981 197374 143212 197376
rect 142797 197371 142863 197372
rect 142981 197371 143047 197374
rect 143206 197372 143212 197374
rect 143276 197372 143282 197436
rect 177990 197434 178050 197510
rect 200614 197434 200620 197436
rect 177990 197374 200620 197434
rect 200614 197372 200620 197374
rect 200684 197372 200690 197436
rect 165102 197236 165108 197300
rect 165172 197298 165178 197300
rect 198733 197298 198799 197301
rect 165172 197296 198799 197298
rect 165172 197240 198738 197296
rect 198794 197240 198799 197296
rect 165172 197238 198799 197240
rect 165172 197236 165178 197238
rect 198733 197235 198799 197238
rect 160829 197162 160895 197165
rect 194593 197162 194659 197165
rect 160829 197160 194659 197162
rect 160829 197104 160834 197160
rect 160890 197104 194598 197160
rect 194654 197104 194659 197160
rect 160829 197102 194659 197104
rect 160829 197099 160895 197102
rect 194593 197099 194659 197102
rect 135529 197028 135595 197029
rect 135478 196964 135484 197028
rect 135548 197026 135595 197028
rect 140037 197026 140103 197029
rect 142102 197026 142108 197028
rect 135548 197024 135640 197026
rect 135590 196968 135640 197024
rect 135548 196966 135640 196968
rect 140037 197024 142108 197026
rect 140037 196968 140042 197024
rect 140098 196968 142108 197024
rect 140037 196966 142108 196968
rect 135548 196964 135595 196966
rect 135529 196963 135595 196964
rect 140037 196963 140103 196966
rect 142102 196964 142108 196966
rect 142172 196964 142178 197028
rect 147254 196964 147260 197028
rect 147324 197026 147330 197028
rect 151813 197026 151879 197029
rect 161054 197026 161060 197028
rect 147324 197024 151879 197026
rect 147324 196968 151818 197024
rect 151874 196968 151879 197024
rect 147324 196966 151879 196968
rect 147324 196964 147330 196966
rect 151813 196963 151879 196966
rect 160326 196966 161060 197026
rect 160326 196893 160386 196966
rect 161054 196964 161060 196966
rect 161124 196964 161130 197028
rect 163681 197026 163747 197029
rect 197445 197026 197511 197029
rect 163681 197024 197511 197026
rect 163681 196968 163686 197024
rect 163742 196968 197450 197024
rect 197506 196968 197511 197024
rect 163681 196966 197511 196968
rect 163681 196963 163747 196966
rect 197445 196963 197511 196966
rect 135437 196892 135503 196893
rect 134006 196828 134012 196892
rect 134076 196890 134082 196892
rect 134742 196890 134748 196892
rect 134076 196830 134748 196890
rect 134076 196828 134082 196830
rect 134742 196828 134748 196830
rect 134812 196828 134818 196892
rect 135437 196888 135484 196892
rect 135548 196890 135554 196892
rect 135437 196832 135442 196888
rect 135437 196828 135484 196832
rect 135548 196830 135594 196890
rect 135548 196828 135554 196830
rect 139526 196828 139532 196892
rect 139596 196890 139602 196892
rect 140405 196890 140471 196893
rect 139596 196888 140471 196890
rect 139596 196832 140410 196888
rect 140466 196832 140471 196888
rect 139596 196830 140471 196832
rect 139596 196828 139602 196830
rect 135437 196827 135503 196828
rect 140405 196827 140471 196830
rect 140589 196892 140655 196893
rect 140589 196888 140636 196892
rect 140700 196890 140706 196892
rect 141509 196890 141575 196893
rect 142286 196890 142292 196892
rect 140589 196832 140594 196888
rect 140589 196828 140636 196832
rect 140700 196830 140746 196890
rect 141509 196888 142292 196890
rect 141509 196832 141514 196888
rect 141570 196832 142292 196888
rect 141509 196830 142292 196832
rect 140700 196828 140706 196830
rect 140589 196827 140655 196828
rect 141509 196827 141575 196830
rect 142286 196828 142292 196830
rect 142356 196828 142362 196892
rect 160277 196888 160386 196893
rect 161105 196892 161171 196893
rect 161054 196890 161060 196892
rect 160277 196832 160282 196888
rect 160338 196832 160386 196888
rect 160277 196830 160386 196832
rect 161014 196830 161060 196890
rect 161124 196888 161171 196892
rect 161166 196832 161171 196888
rect 160277 196827 160343 196830
rect 161054 196828 161060 196830
rect 161124 196828 161171 196832
rect 161105 196827 161171 196828
rect 162853 196890 162919 196893
rect 196014 196890 196020 196892
rect 162853 196888 196020 196890
rect 162853 196832 162858 196888
rect 162914 196832 196020 196888
rect 162853 196830 196020 196832
rect 162853 196827 162919 196830
rect 196014 196828 196020 196830
rect 196084 196828 196090 196892
rect 106774 196692 106780 196756
rect 106844 196754 106850 196756
rect 136357 196754 136423 196757
rect 106844 196752 136423 196754
rect 106844 196696 136362 196752
rect 136418 196696 136423 196752
rect 106844 196694 136423 196696
rect 106844 196692 106850 196694
rect 136357 196691 136423 196694
rect 136582 196692 136588 196756
rect 136652 196754 136658 196756
rect 137369 196754 137435 196757
rect 136652 196752 137435 196754
rect 136652 196696 137374 196752
rect 137430 196696 137435 196752
rect 136652 196694 137435 196696
rect 136652 196692 136658 196694
rect 137369 196691 137435 196694
rect 139669 196754 139735 196757
rect 160921 196756 160987 196757
rect 143758 196754 143764 196756
rect 139669 196752 143764 196754
rect 139669 196696 139674 196752
rect 139730 196696 143764 196752
rect 139669 196694 143764 196696
rect 139669 196691 139735 196694
rect 143758 196692 143764 196694
rect 143828 196692 143834 196756
rect 160870 196692 160876 196756
rect 160940 196754 160987 196756
rect 160940 196752 161032 196754
rect 160982 196696 161032 196752
rect 160940 196694 161032 196696
rect 160940 196692 160987 196694
rect 165838 196692 165844 196756
rect 165908 196754 165914 196756
rect 200389 196754 200455 196757
rect 165908 196752 200455 196754
rect 165908 196696 200394 196752
rect 200450 196696 200455 196752
rect 165908 196694 200455 196696
rect 165908 196692 165914 196694
rect 160921 196691 160987 196692
rect 200389 196691 200455 196694
rect 109953 196618 110019 196621
rect 142705 196618 142771 196621
rect 109953 196616 142771 196618
rect 109953 196560 109958 196616
rect 110014 196560 142710 196616
rect 142766 196560 142771 196616
rect 109953 196558 142771 196560
rect 109953 196555 110019 196558
rect 142705 196555 142771 196558
rect 153929 196618 153995 196621
rect 218145 196618 218211 196621
rect 153929 196616 218211 196618
rect 153929 196560 153934 196616
rect 153990 196560 218150 196616
rect 218206 196560 218211 196616
rect 153929 196558 218211 196560
rect 153929 196555 153995 196558
rect 218145 196555 218211 196558
rect 134149 196484 134215 196485
rect 134149 196480 134196 196484
rect 134260 196482 134266 196484
rect 140773 196482 140839 196485
rect 142470 196482 142476 196484
rect 134149 196424 134154 196480
rect 134149 196420 134196 196424
rect 134260 196422 134306 196482
rect 140773 196480 142476 196482
rect 140773 196424 140778 196480
rect 140834 196424 142476 196480
rect 140773 196422 142476 196424
rect 134260 196420 134266 196422
rect 134149 196419 134215 196420
rect 140773 196419 140839 196422
rect 142470 196420 142476 196422
rect 142540 196420 142546 196484
rect 147489 196482 147555 196485
rect 147622 196482 147628 196484
rect 147489 196480 147628 196482
rect 147489 196424 147494 196480
rect 147550 196424 147628 196480
rect 147489 196422 147628 196424
rect 147489 196419 147555 196422
rect 147622 196420 147628 196422
rect 147692 196420 147698 196484
rect 169886 196420 169892 196484
rect 169956 196482 169962 196484
rect 171133 196482 171199 196485
rect 169956 196480 171199 196482
rect 169956 196424 171138 196480
rect 171194 196424 171199 196480
rect 169956 196422 171199 196424
rect 169956 196420 169962 196422
rect 171133 196419 171199 196422
rect 165981 196348 166047 196349
rect 165981 196346 166028 196348
rect 165936 196344 166028 196346
rect 165936 196288 165986 196344
rect 165936 196286 166028 196288
rect 165981 196284 166028 196286
rect 166092 196284 166098 196348
rect 165981 196283 166047 196284
rect 135662 196012 135668 196076
rect 135732 196074 135738 196076
rect 135897 196074 135963 196077
rect 135732 196072 135963 196074
rect 135732 196016 135902 196072
rect 135958 196016 135963 196072
rect 135732 196014 135963 196016
rect 135732 196012 135738 196014
rect 135897 196011 135963 196014
rect 140221 196074 140287 196077
rect 144269 196076 144335 196077
rect 143574 196074 143580 196076
rect 140221 196072 143580 196074
rect 140221 196016 140226 196072
rect 140282 196016 143580 196072
rect 140221 196014 143580 196016
rect 140221 196011 140287 196014
rect 143574 196012 143580 196014
rect 143644 196012 143650 196076
rect 144269 196074 144316 196076
rect 144224 196072 144316 196074
rect 144224 196016 144274 196072
rect 144224 196014 144316 196016
rect 144269 196012 144316 196014
rect 144380 196012 144386 196076
rect 157793 196074 157859 196077
rect 158294 196074 158300 196076
rect 157793 196072 158300 196074
rect 157793 196016 157798 196072
rect 157854 196016 158300 196072
rect 157793 196014 158300 196016
rect 144269 196011 144335 196012
rect 157793 196011 157859 196014
rect 158294 196012 158300 196014
rect 158364 196012 158370 196076
rect 170990 196012 170996 196076
rect 171060 196074 171066 196076
rect 171777 196074 171843 196077
rect 171060 196072 171843 196074
rect 171060 196016 171782 196072
rect 171838 196016 171843 196072
rect 171060 196014 171843 196016
rect 171060 196012 171066 196014
rect 171777 196011 171843 196014
rect 135294 195876 135300 195940
rect 135364 195938 135370 195940
rect 136173 195938 136239 195941
rect 135364 195936 136239 195938
rect 135364 195880 136178 195936
rect 136234 195880 136239 195936
rect 135364 195878 136239 195880
rect 135364 195876 135370 195878
rect 136173 195875 136239 195878
rect 154062 195876 154068 195940
rect 154132 195938 154138 195940
rect 158989 195938 159055 195941
rect 154132 195936 159055 195938
rect 154132 195880 158994 195936
rect 159050 195880 159055 195936
rect 154132 195878 159055 195880
rect 154132 195876 154138 195878
rect 158989 195875 159055 195878
rect 161422 195876 161428 195940
rect 161492 195938 161498 195940
rect 161565 195938 161631 195941
rect 161492 195936 161631 195938
rect 161492 195880 161570 195936
rect 161626 195880 161631 195936
rect 161492 195878 161631 195880
rect 161492 195876 161498 195878
rect 161565 195875 161631 195878
rect 167269 195938 167335 195941
rect 170949 195940 171015 195941
rect 168046 195938 168052 195940
rect 167269 195936 168052 195938
rect 167269 195880 167274 195936
rect 167330 195880 168052 195936
rect 167269 195878 168052 195880
rect 167269 195875 167335 195878
rect 168046 195876 168052 195878
rect 168116 195876 168122 195940
rect 170949 195936 170996 195940
rect 171060 195938 171066 195940
rect 174905 195938 174971 195941
rect 201718 195938 201724 195940
rect 170949 195880 170954 195936
rect 170949 195876 170996 195880
rect 171060 195878 171106 195938
rect 174905 195936 201724 195938
rect 174905 195880 174910 195936
rect 174966 195880 201724 195936
rect 174905 195878 201724 195880
rect 171060 195876 171066 195878
rect 170949 195875 171015 195876
rect 174905 195875 174971 195878
rect 201718 195876 201724 195878
rect 201788 195876 201794 195940
rect 122373 195802 122439 195805
rect 145189 195802 145255 195805
rect 122373 195800 145255 195802
rect 122373 195744 122378 195800
rect 122434 195744 145194 195800
rect 145250 195744 145255 195800
rect 122373 195742 145255 195744
rect 122373 195739 122439 195742
rect 145189 195739 145255 195742
rect 163773 195802 163839 195805
rect 195973 195802 196039 195805
rect 163773 195800 196039 195802
rect 163773 195744 163778 195800
rect 163834 195744 195978 195800
rect 196034 195744 196039 195800
rect 163773 195742 196039 195744
rect 163773 195739 163839 195742
rect 195973 195739 196039 195742
rect 122189 195666 122255 195669
rect 143349 195666 143415 195669
rect 122189 195664 143415 195666
rect 122189 195608 122194 195664
rect 122250 195608 143354 195664
rect 143410 195608 143415 195664
rect 122189 195606 143415 195608
rect 122189 195603 122255 195606
rect 143349 195603 143415 195606
rect 147581 195666 147647 195669
rect 148910 195666 148916 195668
rect 147581 195664 148916 195666
rect 147581 195608 147586 195664
rect 147642 195608 148916 195664
rect 147581 195606 148916 195608
rect 147581 195603 147647 195606
rect 148910 195604 148916 195606
rect 148980 195604 148986 195668
rect 158662 195604 158668 195668
rect 158732 195666 158738 195668
rect 162301 195666 162367 195669
rect 158732 195664 162367 195666
rect 158732 195608 162306 195664
rect 162362 195608 162367 195664
rect 158732 195606 162367 195608
rect 158732 195604 158738 195606
rect 162301 195603 162367 195606
rect 176285 195666 176351 195669
rect 217133 195666 217199 195669
rect 176285 195664 217199 195666
rect 176285 195608 176290 195664
rect 176346 195608 217138 195664
rect 217194 195608 217199 195664
rect 176285 195606 217199 195608
rect 176285 195603 176351 195606
rect 217133 195603 217199 195606
rect 126421 195530 126487 195533
rect 153101 195530 153167 195533
rect 126421 195528 153167 195530
rect 126421 195472 126426 195528
rect 126482 195472 153106 195528
rect 153162 195472 153167 195528
rect 126421 195470 153167 195472
rect 126421 195467 126487 195470
rect 153101 195467 153167 195470
rect 175181 195530 175247 195533
rect 217225 195530 217291 195533
rect 175181 195528 217291 195530
rect 175181 195472 175186 195528
rect 175242 195472 217230 195528
rect 217286 195472 217291 195528
rect 175181 195470 217291 195472
rect 175181 195467 175247 195470
rect 217225 195467 217291 195470
rect 104617 195394 104683 195397
rect 129641 195394 129707 195397
rect 104617 195392 129707 195394
rect 104617 195336 104622 195392
rect 104678 195336 129646 195392
rect 129702 195336 129707 195392
rect 104617 195334 129707 195336
rect 104617 195331 104683 195334
rect 129641 195331 129707 195334
rect 151721 195394 151787 195397
rect 215753 195394 215819 195397
rect 151721 195392 215819 195394
rect 151721 195336 151726 195392
rect 151782 195336 215758 195392
rect 215814 195336 215819 195392
rect 151721 195334 215819 195336
rect 151721 195331 151787 195334
rect 215753 195331 215819 195334
rect 100569 195258 100635 195261
rect 134609 195258 134675 195261
rect 100569 195256 134675 195258
rect 100569 195200 100574 195256
rect 100630 195200 134614 195256
rect 134670 195200 134675 195256
rect 100569 195198 134675 195200
rect 100569 195195 100635 195198
rect 134609 195195 134675 195198
rect 152549 195258 152615 195261
rect 220905 195258 220971 195261
rect 152549 195256 220971 195258
rect 152549 195200 152554 195256
rect 152610 195200 220910 195256
rect 220966 195200 220971 195256
rect 152549 195198 220971 195200
rect 152549 195195 152615 195198
rect 220905 195195 220971 195198
rect 118182 194516 118188 194580
rect 118252 194578 118258 194580
rect 120717 194578 120783 194581
rect 118252 194576 120783 194578
rect 118252 194520 120722 194576
rect 120778 194520 120783 194576
rect 118252 194518 120783 194520
rect 118252 194516 118258 194518
rect 120717 194515 120783 194518
rect 122966 194380 122972 194444
rect 123036 194442 123042 194444
rect 144126 194442 144132 194444
rect 123036 194382 144132 194442
rect 123036 194380 123042 194382
rect 144126 194380 144132 194382
rect 144196 194380 144202 194444
rect 173525 194442 173591 194445
rect 207054 194442 207060 194444
rect 173525 194440 207060 194442
rect 173525 194384 173530 194440
rect 173586 194384 207060 194440
rect 173525 194382 207060 194384
rect 173525 194379 173591 194382
rect 207054 194380 207060 194382
rect 207124 194380 207130 194444
rect 122414 194244 122420 194308
rect 122484 194306 122490 194308
rect 152774 194306 152780 194308
rect 122484 194246 152780 194306
rect 122484 194244 122490 194246
rect 152774 194244 152780 194246
rect 152844 194244 152850 194308
rect 172646 194244 172652 194308
rect 172716 194306 172722 194308
rect 205582 194306 205588 194308
rect 172716 194246 205588 194306
rect 172716 194244 172722 194246
rect 205582 194244 205588 194246
rect 205652 194244 205658 194308
rect 101990 194108 101996 194172
rect 102060 194170 102066 194172
rect 126605 194170 126671 194173
rect 102060 194168 126671 194170
rect 102060 194112 126610 194168
rect 126666 194112 126671 194168
rect 102060 194110 126671 194112
rect 102060 194108 102066 194110
rect 126605 194107 126671 194110
rect 171961 194170 172027 194173
rect 205766 194170 205772 194172
rect 171961 194168 205772 194170
rect 171961 194112 171966 194168
rect 172022 194112 205772 194168
rect 171961 194110 205772 194112
rect 171961 194107 172027 194110
rect 205766 194108 205772 194110
rect 205836 194108 205842 194172
rect 122598 193972 122604 194036
rect 122668 194034 122674 194036
rect 154849 194034 154915 194037
rect 122668 194032 154915 194034
rect 122668 193976 154854 194032
rect 154910 193976 154915 194032
rect 122668 193974 154915 193976
rect 122668 193972 122674 193974
rect 154849 193971 154915 193974
rect 180609 194034 180675 194037
rect 208485 194034 208551 194037
rect 180609 194032 208551 194034
rect 180609 193976 180614 194032
rect 180670 193976 208490 194032
rect 208546 193976 208551 194032
rect 180609 193974 208551 193976
rect 180609 193971 180675 193974
rect 208485 193971 208551 193974
rect 97206 193836 97212 193900
rect 97276 193898 97282 193900
rect 132033 193898 132099 193901
rect 97276 193896 132099 193898
rect 97276 193840 132038 193896
rect 132094 193840 132099 193896
rect 97276 193838 132099 193840
rect 97276 193836 97282 193838
rect 132033 193835 132099 193838
rect 173893 193898 173959 193901
rect 212625 193898 212691 193901
rect 173893 193896 212691 193898
rect 173893 193840 173898 193896
rect 173954 193840 212630 193896
rect 212686 193840 212691 193896
rect 173893 193838 212691 193840
rect 173893 193835 173959 193838
rect 212625 193835 212691 193838
rect 154246 193292 154252 193356
rect 154316 193354 154322 193356
rect 154389 193354 154455 193357
rect 154316 193352 154455 193354
rect 154316 193296 154394 193352
rect 154450 193296 154455 193352
rect 154316 193294 154455 193296
rect 154316 193292 154322 193294
rect 154389 193291 154455 193294
rect 130561 193218 130627 193221
rect 147806 193218 147812 193220
rect 130561 193216 147812 193218
rect 130561 193160 130566 193216
rect 130622 193160 147812 193216
rect 130561 193158 147812 193160
rect 130561 193155 130627 193158
rect 147806 193156 147812 193158
rect 147876 193156 147882 193220
rect 159030 193156 159036 193220
rect 159100 193218 159106 193220
rect 159449 193218 159515 193221
rect 159100 193216 159515 193218
rect 159100 193160 159454 193216
rect 159510 193160 159515 193216
rect 159100 193158 159515 193160
rect 159100 193156 159106 193158
rect 159449 193155 159515 193158
rect 104014 193020 104020 193084
rect 104084 193082 104090 193084
rect 129733 193082 129799 193085
rect 104084 193080 129799 193082
rect 104084 193024 129738 193080
rect 129794 193024 129799 193080
rect 104084 193022 129799 193024
rect 104084 193020 104090 193022
rect 129733 193019 129799 193022
rect 171133 193082 171199 193085
rect 196198 193082 196204 193084
rect 171133 193080 196204 193082
rect 171133 193024 171138 193080
rect 171194 193024 196204 193080
rect 171133 193022 196204 193024
rect 171133 193019 171199 193022
rect 196198 193020 196204 193022
rect 196268 193020 196274 193084
rect 103421 192946 103487 192949
rect 133873 192946 133939 192949
rect 103421 192944 133939 192946
rect 103421 192888 103426 192944
rect 103482 192888 133878 192944
rect 133934 192888 133939 192944
rect 103421 192886 133939 192888
rect 103421 192883 103487 192886
rect 133873 192883 133939 192886
rect 154113 192946 154179 192949
rect 187734 192946 187740 192948
rect 154113 192944 187740 192946
rect 154113 192888 154118 192944
rect 154174 192888 187740 192944
rect 154113 192886 187740 192888
rect 154113 192883 154179 192886
rect 187734 192884 187740 192886
rect 187804 192884 187810 192948
rect 119838 192748 119844 192812
rect 119908 192810 119914 192812
rect 153561 192810 153627 192813
rect 119908 192808 153627 192810
rect 119908 192752 153566 192808
rect 153622 192752 153627 192808
rect 119908 192750 153627 192752
rect 119908 192748 119914 192750
rect 153561 192747 153627 192750
rect 168925 192810 168991 192813
rect 202965 192810 203031 192813
rect 168925 192808 203031 192810
rect 168925 192752 168930 192808
rect 168986 192752 202970 192808
rect 203026 192752 203031 192808
rect 168925 192750 203031 192752
rect 168925 192747 168991 192750
rect 202965 192747 203031 192750
rect 97717 192674 97783 192677
rect 147990 192674 147996 192676
rect 97717 192672 147996 192674
rect 97717 192616 97722 192672
rect 97778 192616 147996 192672
rect 97717 192614 147996 192616
rect 97717 192611 97783 192614
rect 147990 192612 147996 192614
rect 148060 192612 148066 192676
rect 171409 192674 171475 192677
rect 205909 192674 205975 192677
rect 171409 192672 205975 192674
rect 171409 192616 171414 192672
rect 171470 192616 205914 192672
rect 205970 192616 205975 192672
rect 171409 192614 205975 192616
rect 171409 192611 171475 192614
rect 205909 192611 205975 192614
rect 97533 192538 97599 192541
rect 148174 192538 148180 192540
rect 97533 192536 148180 192538
rect 97533 192480 97538 192536
rect 97594 192480 148180 192536
rect 97533 192478 148180 192480
rect 97533 192475 97599 192478
rect 148174 192476 148180 192478
rect 148244 192476 148250 192540
rect 158621 192538 158687 192541
rect 216673 192538 216739 192541
rect 158621 192536 216739 192538
rect 158621 192480 158626 192536
rect 158682 192480 216678 192536
rect 216734 192480 216739 192536
rect 158621 192478 216739 192480
rect 158621 192475 158687 192478
rect 216673 192475 216739 192478
rect 580349 192538 580415 192541
rect 583520 192538 584960 192628
rect 580349 192536 584960 192538
rect 580349 192480 580354 192536
rect 580410 192480 584960 192536
rect 580349 192478 584960 192480
rect 580349 192475 580415 192478
rect 583520 192388 584960 192478
rect 108798 191524 108804 191588
rect 108868 191586 108874 191588
rect 139393 191586 139459 191589
rect 108868 191584 139459 191586
rect 108868 191528 139398 191584
rect 139454 191528 139459 191584
rect 108868 191526 139459 191528
rect 108868 191524 108874 191526
rect 139393 191523 139459 191526
rect 100518 191388 100524 191452
rect 100588 191450 100594 191452
rect 133689 191450 133755 191453
rect 100588 191448 133755 191450
rect 100588 191392 133694 191448
rect 133750 191392 133755 191448
rect 100588 191390 133755 191392
rect 100588 191388 100594 191390
rect 133689 191387 133755 191390
rect 105997 191314 106063 191317
rect 138422 191314 138428 191316
rect 105997 191312 138428 191314
rect 105997 191256 106002 191312
rect 106058 191256 138428 191312
rect 105997 191254 138428 191256
rect 105997 191251 106063 191254
rect 138422 191252 138428 191254
rect 138492 191252 138498 191316
rect 100334 191116 100340 191180
rect 100404 191178 100410 191180
rect 133321 191178 133387 191181
rect 100404 191176 133387 191178
rect 100404 191120 133326 191176
rect 133382 191120 133387 191176
rect 100404 191118 133387 191120
rect 100404 191116 100410 191118
rect 133321 191115 133387 191118
rect 162342 191116 162348 191180
rect 162412 191178 162418 191180
rect 209865 191178 209931 191181
rect 162412 191176 209931 191178
rect 162412 191120 209870 191176
rect 209926 191120 209931 191176
rect 162412 191118 209931 191120
rect 162412 191116 162418 191118
rect 209865 191115 209931 191118
rect 100661 191042 100727 191045
rect 134006 191042 134012 191044
rect 100661 191040 134012 191042
rect 100661 190984 100666 191040
rect 100722 190984 134012 191040
rect 100661 190982 134012 190984
rect 100661 190979 100727 190982
rect 134006 190980 134012 190982
rect 134076 190980 134082 191044
rect 165286 190980 165292 191044
rect 165356 191042 165362 191044
rect 219433 191042 219499 191045
rect 165356 191040 219499 191042
rect 165356 190984 219438 191040
rect 219494 190984 219499 191040
rect 165356 190982 219499 190984
rect 165356 190980 165362 190982
rect 219433 190979 219499 190982
rect 104382 190300 104388 190364
rect 104452 190362 104458 190364
rect 137001 190362 137067 190365
rect 104452 190360 137067 190362
rect 104452 190304 137006 190360
rect 137062 190304 137067 190360
rect 104452 190302 137067 190304
rect 104452 190300 104458 190302
rect 137001 190299 137067 190302
rect 104198 190164 104204 190228
rect 104268 190226 104274 190228
rect 136817 190226 136883 190229
rect 104268 190224 136883 190226
rect 104268 190168 136822 190224
rect 136878 190168 136883 190224
rect 104268 190166 136883 190168
rect 104268 190164 104274 190166
rect 136817 190163 136883 190166
rect 176326 190164 176332 190228
rect 176396 190226 176402 190228
rect 209814 190226 209820 190228
rect 176396 190166 209820 190226
rect 176396 190164 176402 190166
rect 209814 190164 209820 190166
rect 209884 190164 209890 190228
rect 107193 190090 107259 190093
rect 142286 190090 142292 190092
rect 107193 190088 142292 190090
rect 107193 190032 107198 190088
rect 107254 190032 142292 190088
rect 107193 190030 142292 190032
rect 107193 190027 107259 190030
rect 142286 190028 142292 190030
rect 142356 190028 142362 190092
rect 174670 190028 174676 190092
rect 174740 190090 174746 190092
rect 208393 190090 208459 190093
rect 174740 190088 208459 190090
rect 174740 190032 208398 190088
rect 208454 190032 208459 190088
rect 174740 190030 208459 190032
rect 174740 190028 174746 190030
rect 208393 190027 208459 190030
rect 107009 189954 107075 189957
rect 142470 189954 142476 189956
rect 107009 189952 142476 189954
rect 107009 189896 107014 189952
rect 107070 189896 142476 189952
rect 107009 189894 142476 189896
rect 107009 189891 107075 189894
rect 142470 189892 142476 189894
rect 142540 189892 142546 189956
rect 159030 189892 159036 189956
rect 159100 189954 159106 189956
rect 209773 189954 209839 189957
rect 159100 189952 209839 189954
rect 159100 189896 209778 189952
rect 209834 189896 209839 189952
rect 159100 189894 209839 189896
rect 159100 189892 159106 189894
rect 209773 189891 209839 189894
rect 107101 189818 107167 189821
rect 143758 189818 143764 189820
rect 107101 189816 143764 189818
rect 107101 189760 107106 189816
rect 107162 189760 143764 189816
rect 107101 189758 143764 189760
rect 107101 189755 107167 189758
rect 143758 189756 143764 189758
rect 143828 189756 143834 189820
rect 157006 189756 157012 189820
rect 157076 189818 157082 189820
rect 211153 189818 211219 189821
rect 157076 189816 211219 189818
rect 157076 189760 211158 189816
rect 211214 189760 211219 189816
rect 157076 189758 211219 189760
rect 157076 189756 157082 189758
rect 211153 189755 211219 189758
rect 105537 189682 105603 189685
rect 143574 189682 143580 189684
rect 105537 189680 143580 189682
rect 105537 189624 105542 189680
rect 105598 189624 143580 189680
rect 105537 189622 143580 189624
rect 105537 189619 105603 189622
rect 143574 189620 143580 189622
rect 143644 189620 143650 189684
rect 154246 189620 154252 189684
rect 154316 189682 154322 189684
rect 221273 189682 221339 189685
rect 154316 189680 221339 189682
rect 154316 189624 221278 189680
rect 221334 189624 221339 189680
rect 154316 189622 221339 189624
rect 154316 189620 154322 189622
rect 221273 189619 221339 189622
rect 124806 189484 124812 189548
rect 124876 189546 124882 189548
rect 151629 189546 151695 189549
rect 124876 189544 151695 189546
rect 124876 189488 151634 189544
rect 151690 189488 151695 189544
rect 124876 189486 151695 189488
rect 124876 189484 124882 189486
rect 151629 189483 151695 189486
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 106181 187642 106247 187645
rect 138238 187642 138244 187644
rect 106181 187640 138244 187642
rect 106181 187584 106186 187640
rect 106242 187584 138244 187640
rect 106181 187582 138244 187584
rect 106181 187579 106247 187582
rect 138238 187580 138244 187582
rect 138308 187580 138314 187644
rect 103278 187444 103284 187508
rect 103348 187506 103354 187508
rect 135662 187506 135668 187508
rect 103348 187446 135668 187506
rect 103348 187444 103354 187446
rect 135662 187444 135668 187446
rect 135732 187444 135738 187508
rect 120574 187308 120580 187372
rect 120644 187370 120650 187372
rect 153745 187370 153811 187373
rect 120644 187368 153811 187370
rect 120644 187312 153750 187368
rect 153806 187312 153811 187368
rect 120644 187310 153811 187312
rect 120644 187308 120650 187310
rect 153745 187307 153811 187310
rect 99230 187172 99236 187236
rect 99300 187234 99306 187236
rect 132861 187234 132927 187237
rect 99300 187232 132927 187234
rect 99300 187176 132866 187232
rect 132922 187176 132927 187232
rect 99300 187174 132927 187176
rect 99300 187172 99306 187174
rect 132861 187171 132927 187174
rect 102041 187098 102107 187101
rect 135478 187098 135484 187100
rect 102041 187096 135484 187098
rect 102041 187040 102046 187096
rect 102102 187040 135484 187096
rect 102041 187038 135484 187040
rect 102041 187035 102107 187038
rect 135478 187036 135484 187038
rect 135548 187036 135554 187100
rect 169385 187098 169451 187101
rect 187182 187098 187188 187100
rect 169385 187096 187188 187098
rect 169385 187040 169390 187096
rect 169446 187040 187188 187096
rect 169385 187038 187188 187040
rect 169385 187035 169451 187038
rect 187182 187036 187188 187038
rect 187252 187036 187258 187100
rect 115606 186900 115612 186964
rect 115676 186962 115682 186964
rect 152825 186962 152891 186965
rect 115676 186960 152891 186962
rect 115676 186904 152830 186960
rect 152886 186904 152891 186960
rect 115676 186902 152891 186904
rect 115676 186900 115682 186902
rect 152825 186899 152891 186902
rect 167862 186900 167868 186964
rect 167932 186962 167938 186964
rect 214097 186962 214163 186965
rect 167932 186960 214163 186962
rect 167932 186904 214102 186960
rect 214158 186904 214163 186960
rect 167932 186902 214163 186904
rect 167932 186900 167938 186902
rect 214097 186899 214163 186902
rect 147581 186420 147647 186421
rect 147581 186418 147628 186420
rect 147536 186416 147628 186418
rect 147536 186360 147586 186416
rect 147536 186358 147628 186360
rect 147581 186356 147628 186358
rect 147692 186356 147698 186420
rect 147581 186355 147647 186356
rect 580349 179210 580415 179213
rect 583520 179210 584960 179300
rect 580349 179208 584960 179210
rect 580349 179152 580354 179208
rect 580410 179152 584960 179208
rect 580349 179150 584960 179152
rect 580349 179147 580415 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3509 162890 3575 162893
rect -960 162888 3575 162890
rect -960 162832 3514 162888
rect 3570 162832 3575 162888
rect -960 162830 3575 162832
rect -960 162740 480 162830
rect 3509 162827 3575 162830
rect 168046 158068 168052 158132
rect 168116 158130 168122 158132
rect 201861 158130 201927 158133
rect 168116 158128 201927 158130
rect 168116 158072 201866 158128
rect 201922 158072 201927 158128
rect 168116 158070 201927 158072
rect 168116 158068 168122 158070
rect 201861 158067 201927 158070
rect 177021 157994 177087 157997
rect 211102 157994 211108 157996
rect 177021 157992 211108 157994
rect 177021 157936 177026 157992
rect 177082 157936 211108 157992
rect 177021 157934 211108 157936
rect 177021 157931 177087 157934
rect 211102 157932 211108 157934
rect 211172 157932 211178 157996
rect 165470 155756 165476 155820
rect 165540 155818 165546 155820
rect 185945 155818 186011 155821
rect 165540 155816 186011 155818
rect 165540 155760 185950 155816
rect 186006 155760 186011 155816
rect 165540 155758 186011 155760
rect 165540 155756 165546 155758
rect 185945 155755 186011 155758
rect 154062 155620 154068 155684
rect 154132 155682 154138 155684
rect 187049 155682 187115 155685
rect 154132 155680 187115 155682
rect 154132 155624 187054 155680
rect 187110 155624 187115 155680
rect 154132 155622 187115 155624
rect 154132 155620 154138 155622
rect 187049 155619 187115 155622
rect 169334 155484 169340 155548
rect 169404 155546 169410 155548
rect 203333 155546 203399 155549
rect 169404 155544 203399 155546
rect 169404 155488 203338 155544
rect 203394 155488 203399 155544
rect 169404 155486 203399 155488
rect 169404 155484 169410 155486
rect 203333 155483 203399 155486
rect 176929 155410 176995 155413
rect 211286 155410 211292 155412
rect 176929 155408 211292 155410
rect 176929 155352 176934 155408
rect 176990 155352 211292 155408
rect 176929 155350 211292 155352
rect 176929 155347 176995 155350
rect 211286 155348 211292 155350
rect 211356 155348 211362 155412
rect 168230 155212 168236 155276
rect 168300 155274 168306 155276
rect 215569 155274 215635 155277
rect 168300 155272 215635 155274
rect 168300 155216 215574 155272
rect 215630 155216 215635 155272
rect 168300 155214 215635 155216
rect 168300 155212 168306 155214
rect 215569 155211 215635 155214
rect 96521 153778 96587 153781
rect 139526 153778 139532 153780
rect 96521 153776 139532 153778
rect 96521 153720 96526 153776
rect 96582 153720 139532 153776
rect 96521 153718 139532 153720
rect 96521 153715 96587 153718
rect 139526 153716 139532 153718
rect 139596 153716 139602 153780
rect 175641 152826 175707 152829
rect 203190 152826 203196 152828
rect 175641 152824 203196 152826
rect 175641 152768 175646 152824
rect 175702 152768 203196 152824
rect 175641 152766 203196 152768
rect 175641 152763 175707 152766
rect 203190 152764 203196 152766
rect 203260 152764 203266 152828
rect 157190 152628 157196 152692
rect 157260 152690 157266 152692
rect 195421 152690 195487 152693
rect 157260 152688 195487 152690
rect 157260 152632 195426 152688
rect 195482 152632 195487 152688
rect 157260 152630 195487 152632
rect 157260 152628 157266 152630
rect 195421 152627 195487 152630
rect 580073 152690 580139 152693
rect 583520 152690 584960 152780
rect 580073 152688 584960 152690
rect 580073 152632 580078 152688
rect 580134 152632 584960 152688
rect 580073 152630 584960 152632
rect 580073 152627 580139 152630
rect 161054 152492 161060 152556
rect 161124 152554 161130 152556
rect 218513 152554 218579 152557
rect 161124 152552 218579 152554
rect 161124 152496 218518 152552
rect 218574 152496 218579 152552
rect 583520 152540 584960 152630
rect 161124 152494 218579 152496
rect 161124 152492 161130 152494
rect 218513 152491 218579 152494
rect 112846 152356 112852 152420
rect 112916 152418 112922 152420
rect 171685 152418 171751 152421
rect 112916 152416 171751 152418
rect 112916 152360 171690 152416
rect 171746 152360 171751 152416
rect 112916 152358 171751 152360
rect 112916 152356 112922 152358
rect 171685 152355 171751 152358
rect 176837 152418 176903 152421
rect 209998 152418 210004 152420
rect 176837 152416 210004 152418
rect 176837 152360 176842 152416
rect 176898 152360 210004 152416
rect 176837 152358 210004 152360
rect 176837 152355 176903 152358
rect 209998 152356 210004 152358
rect 210068 152356 210074 152420
rect 166574 151268 166580 151332
rect 166644 151330 166650 151332
rect 196382 151330 196388 151332
rect 166644 151270 196388 151330
rect 166644 151268 166650 151270
rect 196382 151268 196388 151270
rect 196452 151268 196458 151332
rect 104750 151132 104756 151196
rect 104820 151194 104826 151196
rect 136766 151194 136772 151196
rect 104820 151134 136772 151194
rect 104820 151132 104826 151134
rect 136766 151132 136772 151134
rect 136836 151132 136842 151196
rect 167177 151194 167243 151197
rect 197302 151194 197308 151196
rect 167177 151192 197308 151194
rect 167177 151136 167182 151192
rect 167238 151136 197308 151192
rect 167177 151134 197308 151136
rect 167177 151131 167243 151134
rect 197302 151132 197308 151134
rect 197372 151132 197378 151196
rect 100201 151058 100267 151061
rect 134190 151058 134196 151060
rect 100201 151056 134196 151058
rect 100201 151000 100206 151056
rect 100262 151000 134196 151056
rect 100201 150998 134196 151000
rect 100201 150995 100267 150998
rect 134190 150996 134196 150998
rect 134260 150996 134266 151060
rect 160686 150996 160692 151060
rect 160756 151058 160762 151060
rect 201953 151058 202019 151061
rect 160756 151056 202019 151058
rect 160756 151000 201958 151056
rect 202014 151000 202019 151056
rect 160756 150998 202019 151000
rect 160756 150996 160762 150998
rect 201953 150995 202019 150998
rect 117865 150514 117931 150517
rect 580257 150514 580323 150517
rect 117865 150512 580323 150514
rect 117865 150456 117870 150512
rect 117926 150456 580262 150512
rect 580318 150456 580323 150512
rect 117865 150454 580323 150456
rect 117865 150451 117931 150454
rect 580257 150451 580323 150454
rect 175457 150106 175523 150109
rect 200982 150106 200988 150108
rect 175457 150104 200988 150106
rect 175457 150048 175462 150104
rect 175518 150048 200988 150104
rect 175457 150046 200988 150048
rect 175457 150043 175523 150046
rect 200982 150044 200988 150046
rect 201052 150044 201058 150108
rect 175273 149970 175339 149973
rect 206134 149970 206140 149972
rect 175273 149968 206140 149970
rect -960 149834 480 149924
rect 175273 149912 175278 149968
rect 175334 149912 206140 149968
rect 175273 149910 206140 149912
rect 175273 149907 175339 149910
rect 206134 149908 206140 149910
rect 206204 149908 206210 149972
rect 3141 149834 3207 149837
rect -960 149832 3207 149834
rect -960 149776 3146 149832
rect 3202 149776 3207 149832
rect -960 149774 3207 149776
rect -960 149684 480 149774
rect 3141 149771 3207 149774
rect 172789 149834 172855 149837
rect 205950 149834 205956 149836
rect 172789 149832 205956 149834
rect 172789 149776 172794 149832
rect 172850 149776 205956 149832
rect 172789 149774 205956 149776
rect 172789 149771 172855 149774
rect 205950 149772 205956 149774
rect 206020 149772 206026 149836
rect 172605 149698 172671 149701
rect 207238 149698 207244 149700
rect 172605 149696 207244 149698
rect 172605 149640 172610 149696
rect 172666 149640 207244 149696
rect 172605 149638 207244 149640
rect 172605 149635 172671 149638
rect 207238 149636 207244 149638
rect 207308 149636 207314 149700
rect 123569 148882 123635 148885
rect 140814 148882 140820 148884
rect 123569 148880 140820 148882
rect 123569 148824 123574 148880
rect 123630 148824 140820 148880
rect 123569 148822 140820 148824
rect 123569 148819 123635 148822
rect 140814 148820 140820 148822
rect 140884 148820 140890 148884
rect 108430 148684 108436 148748
rect 108500 148746 108506 148748
rect 132125 148746 132191 148749
rect 108500 148744 132191 148746
rect 108500 148688 132130 148744
rect 132186 148688 132191 148744
rect 108500 148686 132191 148688
rect 108500 148684 108506 148686
rect 132125 148683 132191 148686
rect 121310 148548 121316 148612
rect 121380 148610 121386 148612
rect 150801 148610 150867 148613
rect 121380 148608 150867 148610
rect 121380 148552 150806 148608
rect 150862 148552 150867 148608
rect 121380 148550 150867 148552
rect 121380 148548 121386 148550
rect 150801 148547 150867 148550
rect 167085 148610 167151 148613
rect 193622 148610 193628 148612
rect 167085 148608 193628 148610
rect 167085 148552 167090 148608
rect 167146 148552 193628 148608
rect 167085 148550 193628 148552
rect 167085 148547 167151 148550
rect 193622 148548 193628 148550
rect 193692 148548 193698 148612
rect 122046 148412 122052 148476
rect 122116 148474 122122 148476
rect 153377 148474 153443 148477
rect 122116 148472 153443 148474
rect 122116 148416 153382 148472
rect 153438 148416 153443 148472
rect 122116 148414 153443 148416
rect 122116 148412 122122 148414
rect 153377 148411 153443 148414
rect 163814 148412 163820 148476
rect 163884 148474 163890 148476
rect 191598 148474 191604 148476
rect 163884 148414 191604 148474
rect 163884 148412 163890 148414
rect 191598 148412 191604 148414
rect 191668 148412 191674 148476
rect 101581 148338 101647 148341
rect 135294 148338 135300 148340
rect 101581 148336 135300 148338
rect 101581 148280 101586 148336
rect 101642 148280 135300 148336
rect 101581 148278 135300 148280
rect 101581 148275 101647 148278
rect 135294 148276 135300 148278
rect 135364 148276 135370 148340
rect 169518 148276 169524 148340
rect 169588 148338 169594 148340
rect 203241 148338 203307 148341
rect 169588 148336 203307 148338
rect 169588 148280 203246 148336
rect 203302 148280 203307 148336
rect 169588 148278 203307 148280
rect 169588 148276 169594 148278
rect 203241 148275 203307 148278
rect 112662 147596 112668 147660
rect 112732 147658 112738 147660
rect 138657 147658 138723 147661
rect 112732 147656 138723 147658
rect 112732 147600 138662 147656
rect 138718 147600 138723 147656
rect 112732 147598 138723 147600
rect 112732 147596 112738 147598
rect 138657 147595 138723 147598
rect 183185 147658 183251 147661
rect 187918 147658 187924 147660
rect 183185 147656 187924 147658
rect 183185 147600 183190 147656
rect 183246 147600 187924 147656
rect 183185 147598 187924 147600
rect 183185 147595 183251 147598
rect 187918 147596 187924 147598
rect 187988 147596 187994 147660
rect 113541 147522 113607 147525
rect 142654 147522 142660 147524
rect 113541 147520 142660 147522
rect 113541 147464 113546 147520
rect 113602 147464 142660 147520
rect 113541 147462 142660 147464
rect 113541 147459 113607 147462
rect 142654 147460 142660 147462
rect 142724 147460 142730 147524
rect 171225 147522 171291 147525
rect 197670 147522 197676 147524
rect 171225 147520 197676 147522
rect 171225 147464 171230 147520
rect 171286 147464 197676 147520
rect 171225 147462 197676 147464
rect 171225 147459 171291 147462
rect 197670 147460 197676 147462
rect 197740 147460 197746 147524
rect 112478 147324 112484 147388
rect 112548 147386 112554 147388
rect 143533 147386 143599 147389
rect 112548 147384 143599 147386
rect 112548 147328 143538 147384
rect 143594 147328 143599 147384
rect 112548 147326 143599 147328
rect 112548 147324 112554 147326
rect 143533 147323 143599 147326
rect 169937 147386 170003 147389
rect 197486 147386 197492 147388
rect 169937 147384 197492 147386
rect 169937 147328 169942 147384
rect 169998 147328 197492 147384
rect 169937 147326 197492 147328
rect 169937 147323 170003 147326
rect 197486 147324 197492 147326
rect 197556 147324 197562 147388
rect 108614 147188 108620 147252
rect 108684 147250 108690 147252
rect 139342 147250 139348 147252
rect 108684 147190 139348 147250
rect 108684 147188 108690 147190
rect 139342 147188 139348 147190
rect 139412 147188 139418 147252
rect 166206 147188 166212 147252
rect 166276 147250 166282 147252
rect 199142 147250 199148 147252
rect 166276 147190 199148 147250
rect 166276 147188 166282 147190
rect 199142 147188 199148 147190
rect 199212 147188 199218 147252
rect 110822 147052 110828 147116
rect 110892 147114 110898 147116
rect 142153 147114 142219 147117
rect 110892 147112 142219 147114
rect 110892 147056 142158 147112
rect 142214 147056 142219 147112
rect 110892 147054 142219 147056
rect 110892 147052 110898 147054
rect 142153 147051 142219 147054
rect 170990 147052 170996 147116
rect 171060 147114 171066 147116
rect 204713 147114 204779 147117
rect 171060 147112 204779 147114
rect 171060 147056 204718 147112
rect 204774 147056 204779 147112
rect 171060 147054 204779 147056
rect 171060 147052 171066 147054
rect 204713 147051 204779 147054
rect 107142 146916 107148 146980
rect 107212 146978 107218 146980
rect 138054 146978 138060 146980
rect 107212 146918 138060 146978
rect 107212 146916 107218 146918
rect 138054 146916 138060 146918
rect 138124 146916 138130 146980
rect 150014 146916 150020 146980
rect 150084 146978 150090 146980
rect 196709 146978 196775 146981
rect 150084 146976 196775 146978
rect 150084 146920 196714 146976
rect 196770 146920 196775 146976
rect 150084 146918 196775 146920
rect 150084 146916 150090 146918
rect 196709 146915 196775 146918
rect 119654 146780 119660 146844
rect 119724 146842 119730 146844
rect 136582 146842 136588 146844
rect 119724 146782 136588 146842
rect 119724 146780 119730 146782
rect 136582 146780 136588 146782
rect 136652 146780 136658 146844
rect 109534 146236 109540 146300
rect 109604 146298 109610 146300
rect 131849 146298 131915 146301
rect 109604 146296 131915 146298
rect 109604 146240 131854 146296
rect 131910 146240 131915 146296
rect 109604 146238 131915 146240
rect 109604 146236 109610 146238
rect 131849 146235 131915 146238
rect 115790 146100 115796 146164
rect 115860 146162 115866 146164
rect 142245 146162 142311 146165
rect 115860 146160 142311 146162
rect 115860 146104 142250 146160
rect 142306 146104 142311 146160
rect 115860 146102 142311 146104
rect 115860 146100 115866 146102
rect 142245 146099 142311 146102
rect 180333 146162 180399 146165
rect 191782 146162 191788 146164
rect 180333 146160 191788 146162
rect 180333 146104 180338 146160
rect 180394 146104 191788 146160
rect 180333 146102 191788 146104
rect 180333 146099 180399 146102
rect 191782 146100 191788 146102
rect 191852 146100 191858 146164
rect 111558 145964 111564 146028
rect 111628 146026 111634 146028
rect 144361 146026 144427 146029
rect 111628 146024 144427 146026
rect 111628 145968 144366 146024
rect 144422 145968 144427 146024
rect 111628 145966 144427 145968
rect 111628 145964 111634 145966
rect 144361 145963 144427 145966
rect 171777 146026 171843 146029
rect 189206 146026 189212 146028
rect 171777 146024 189212 146026
rect 171777 145968 171782 146024
rect 171838 145968 189212 146024
rect 171777 145966 189212 145968
rect 171777 145963 171843 145966
rect 189206 145964 189212 145966
rect 189276 145964 189282 146028
rect 113950 145828 113956 145892
rect 114020 145890 114026 145892
rect 146753 145890 146819 145893
rect 114020 145888 146819 145890
rect 114020 145832 146758 145888
rect 146814 145832 146819 145888
rect 114020 145830 146819 145832
rect 114020 145828 114026 145830
rect 146753 145827 146819 145830
rect 163957 145890 164023 145893
rect 191966 145890 191972 145892
rect 163957 145888 191972 145890
rect 163957 145832 163962 145888
rect 164018 145832 191972 145888
rect 163957 145830 191972 145832
rect 163957 145827 164023 145830
rect 191966 145828 191972 145830
rect 192036 145828 192042 145892
rect 116342 145692 116348 145756
rect 116412 145754 116418 145756
rect 153285 145754 153351 145757
rect 116412 145752 153351 145754
rect 116412 145696 153290 145752
rect 153346 145696 153351 145752
rect 116412 145694 153351 145696
rect 116412 145692 116418 145694
rect 153285 145691 153351 145694
rect 166993 145754 167059 145757
rect 198774 145754 198780 145756
rect 166993 145752 198780 145754
rect 166993 145696 166998 145752
rect 167054 145696 198780 145752
rect 166993 145694 198780 145696
rect 166993 145691 167059 145694
rect 198774 145692 198780 145694
rect 198844 145692 198850 145756
rect 111374 145556 111380 145620
rect 111444 145618 111450 145620
rect 146293 145618 146359 145621
rect 111444 145616 146359 145618
rect 111444 145560 146298 145616
rect 146354 145560 146359 145616
rect 111444 145558 146359 145560
rect 111444 145556 111450 145558
rect 146293 145555 146359 145558
rect 147438 145556 147444 145620
rect 147508 145618 147514 145620
rect 195513 145618 195579 145621
rect 147508 145616 195579 145618
rect 147508 145560 195518 145616
rect 195574 145560 195579 145616
rect 147508 145558 195579 145560
rect 147508 145556 147514 145558
rect 195513 145555 195579 145558
rect 113030 144740 113036 144804
rect 113100 144802 113106 144804
rect 145557 144802 145623 144805
rect 113100 144800 145623 144802
rect 113100 144744 145562 144800
rect 145618 144744 145623 144800
rect 113100 144742 145623 144744
rect 113100 144740 113106 144742
rect 145557 144739 145623 144742
rect 180425 144802 180491 144805
rect 189758 144802 189764 144804
rect 180425 144800 189764 144802
rect 180425 144744 180430 144800
rect 180486 144744 189764 144800
rect 180425 144742 189764 144744
rect 180425 144739 180491 144742
rect 189758 144740 189764 144742
rect 189828 144740 189834 144804
rect 118182 144604 118188 144668
rect 118252 144666 118258 144668
rect 151077 144666 151143 144669
rect 118252 144664 151143 144666
rect 118252 144608 151082 144664
rect 151138 144608 151143 144664
rect 118252 144606 151143 144608
rect 118252 144604 118258 144606
rect 151077 144603 151143 144606
rect 164141 144666 164207 144669
rect 193254 144666 193260 144668
rect 164141 144664 193260 144666
rect 164141 144608 164146 144664
rect 164202 144608 193260 144664
rect 164141 144606 193260 144608
rect 164141 144603 164207 144606
rect 193254 144604 193260 144606
rect 193324 144604 193330 144668
rect 115013 144530 115079 144533
rect 147622 144530 147628 144532
rect 115013 144528 147628 144530
rect 115013 144472 115018 144528
rect 115074 144472 147628 144528
rect 115013 144470 147628 144472
rect 115013 144467 115079 144470
rect 147622 144468 147628 144470
rect 147692 144468 147698 144532
rect 162761 144530 162827 144533
rect 193438 144530 193444 144532
rect 162761 144528 193444 144530
rect 162761 144472 162766 144528
rect 162822 144472 193444 144528
rect 162761 144470 193444 144472
rect 162761 144467 162827 144470
rect 193438 144468 193444 144470
rect 193508 144468 193514 144532
rect 118182 144332 118188 144396
rect 118252 144394 118258 144396
rect 151905 144394 151971 144397
rect 118252 144392 151971 144394
rect 118252 144336 151910 144392
rect 151966 144336 151971 144392
rect 118252 144334 151971 144336
rect 118252 144332 118258 144334
rect 151905 144331 151971 144334
rect 154573 144394 154639 144397
rect 189022 144394 189028 144396
rect 154573 144392 189028 144394
rect 154573 144336 154578 144392
rect 154634 144336 189028 144392
rect 154573 144334 189028 144336
rect 154573 144331 154639 144334
rect 189022 144332 189028 144334
rect 189092 144332 189098 144396
rect 115238 144196 115244 144260
rect 115308 144258 115314 144260
rect 152457 144258 152523 144261
rect 115308 144256 152523 144258
rect 115308 144200 152462 144256
rect 152518 144200 152523 144256
rect 115308 144198 152523 144200
rect 115308 144196 115314 144198
rect 152457 144195 152523 144198
rect 154297 144258 154363 144261
rect 187693 144258 187759 144261
rect 154297 144256 187759 144258
rect 154297 144200 154302 144256
rect 154358 144200 187698 144256
rect 187754 144200 187759 144256
rect 154297 144198 187759 144200
rect 154297 144195 154363 144198
rect 187693 144195 187759 144198
rect 113950 144060 113956 144124
rect 114020 144122 114026 144124
rect 151997 144122 152063 144125
rect 114020 144120 152063 144122
rect 114020 144064 152002 144120
rect 152058 144064 152063 144120
rect 114020 144062 152063 144064
rect 114020 144060 114026 144062
rect 151997 144059 152063 144062
rect 152641 144122 152707 144125
rect 186998 144122 187004 144124
rect 152641 144120 187004 144122
rect 152641 144064 152646 144120
rect 152702 144064 187004 144120
rect 152641 144062 187004 144064
rect 152641 144059 152707 144062
rect 186998 144060 187004 144062
rect 187068 144060 187074 144124
rect 118366 143380 118372 143444
rect 118436 143442 118442 143444
rect 145097 143442 145163 143445
rect 118436 143440 145163 143442
rect 118436 143384 145102 143440
rect 145158 143384 145163 143440
rect 118436 143382 145163 143384
rect 118436 143380 118442 143382
rect 145097 143379 145163 143382
rect 118366 143244 118372 143308
rect 118436 143306 118442 143308
rect 146937 143306 147003 143309
rect 118436 143304 147003 143306
rect 118436 143248 146942 143304
rect 146998 143248 147003 143304
rect 118436 143246 147003 143248
rect 118436 143244 118442 143246
rect 146937 143243 147003 143246
rect 118550 143108 118556 143172
rect 118620 143170 118626 143172
rect 148317 143170 148383 143173
rect 118620 143168 148383 143170
rect 118620 143112 148322 143168
rect 148378 143112 148383 143168
rect 118620 143110 148383 143112
rect 118620 143108 118626 143110
rect 148317 143107 148383 143110
rect 162209 143170 162275 143173
rect 189441 143170 189507 143173
rect 162209 143168 189507 143170
rect 162209 143112 162214 143168
rect 162270 143112 189446 143168
rect 189502 143112 189507 143168
rect 162209 143110 189507 143112
rect 162209 143107 162275 143110
rect 189441 143107 189507 143110
rect 117078 142972 117084 143036
rect 117148 143034 117154 143036
rect 146661 143034 146727 143037
rect 117148 143032 146727 143034
rect 117148 142976 146666 143032
rect 146722 142976 146727 143032
rect 117148 142974 146727 142976
rect 117148 142972 117154 142974
rect 146661 142971 146727 142974
rect 163865 143034 163931 143037
rect 191005 143034 191071 143037
rect 163865 143032 191071 143034
rect 163865 142976 163870 143032
rect 163926 142976 191010 143032
rect 191066 142976 191071 143032
rect 163865 142974 191071 142976
rect 163865 142971 163931 142974
rect 191005 142971 191071 142974
rect 116894 142836 116900 142900
rect 116964 142898 116970 142900
rect 149973 142898 150039 142901
rect 116964 142896 150039 142898
rect 116964 142840 149978 142896
rect 150034 142840 150039 142896
rect 116964 142838 150039 142840
rect 116964 142836 116970 142838
rect 149973 142835 150039 142838
rect 157241 142898 157307 142901
rect 189165 142898 189231 142901
rect 157241 142896 189231 142898
rect 157241 142840 157246 142896
rect 157302 142840 189170 142896
rect 189226 142840 189231 142896
rect 157241 142838 189231 142840
rect 157241 142835 157307 142838
rect 189165 142835 189231 142838
rect 111006 142700 111012 142764
rect 111076 142762 111082 142764
rect 183461 142762 183527 142765
rect 111076 142760 183527 142762
rect 111076 142704 183466 142760
rect 183522 142704 183527 142760
rect 111076 142702 183527 142704
rect 111076 142700 111082 142702
rect 183461 142699 183527 142702
rect 111190 142564 111196 142628
rect 111260 142626 111266 142628
rect 124857 142626 124923 142629
rect 111260 142624 124923 142626
rect 111260 142568 124862 142624
rect 124918 142568 124923 142624
rect 111260 142566 124923 142568
rect 111260 142564 111266 142566
rect 124857 142563 124923 142566
rect 124857 142218 124923 142221
rect 580349 142218 580415 142221
rect 124857 142216 580415 142218
rect 124857 142160 124862 142216
rect 124918 142160 580354 142216
rect 580410 142160 580415 142216
rect 124857 142158 580415 142160
rect 124857 142155 124923 142158
rect 580349 142155 580415 142158
rect 117865 142082 117931 142085
rect 123661 142082 123727 142085
rect 117865 142080 123727 142082
rect 117865 142024 117870 142080
rect 117926 142024 123666 142080
rect 123722 142024 123727 142080
rect 117865 142022 123727 142024
rect 117865 142019 117931 142022
rect 123661 142019 123727 142022
rect 118325 141538 118391 141541
rect 139485 141538 139551 141541
rect 118325 141536 139551 141538
rect 118325 141480 118330 141536
rect 118386 141480 139490 141536
rect 139546 141480 139551 141536
rect 118325 141478 139551 141480
rect 118325 141475 118391 141478
rect 139485 141475 139551 141478
rect 162669 141538 162735 141541
rect 189574 141538 189580 141540
rect 162669 141536 189580 141538
rect 162669 141480 162674 141536
rect 162730 141480 189580 141536
rect 162669 141478 189580 141480
rect 162669 141475 162735 141478
rect 189574 141476 189580 141478
rect 189644 141476 189650 141540
rect 114134 141340 114140 141404
rect 114204 141402 114210 141404
rect 136725 141402 136791 141405
rect 114204 141400 136791 141402
rect 114204 141344 136730 141400
rect 136786 141344 136791 141400
rect 114204 141342 136791 141344
rect 114204 141340 114210 141342
rect 136725 141339 136791 141342
rect 161105 141402 161171 141405
rect 194041 141402 194107 141405
rect 161105 141400 194107 141402
rect 161105 141344 161110 141400
rect 161166 141344 194046 141400
rect 194102 141344 194107 141400
rect 161105 141342 194107 141344
rect 161105 141339 161171 141342
rect 194041 141339 194107 141342
rect 116526 141204 116532 141268
rect 116596 141266 116602 141268
rect 183645 141266 183711 141269
rect 184841 141266 184907 141269
rect 116596 141264 184907 141266
rect 116596 141208 183650 141264
rect 183706 141208 184846 141264
rect 184902 141208 184907 141264
rect 116596 141206 184907 141208
rect 116596 141204 116602 141206
rect 183645 141203 183711 141206
rect 184841 141203 184907 141206
rect 127433 141130 127499 141133
rect 482277 141130 482343 141133
rect 127433 141128 482343 141130
rect 127433 141072 127438 141128
rect 127494 141072 482282 141128
rect 482338 141072 482343 141128
rect 127433 141070 482343 141072
rect 127433 141067 127499 141070
rect 482277 141067 482343 141070
rect 127525 140994 127591 140997
rect 580717 140994 580783 140997
rect 127525 140992 580783 140994
rect 127525 140936 127530 140992
rect 127586 140936 580722 140992
rect 580778 140936 580783 140992
rect 127525 140934 580783 140936
rect 127525 140931 127591 140934
rect 580717 140931 580783 140934
rect 118550 140796 118556 140860
rect 118620 140858 118626 140860
rect 122465 140858 122531 140861
rect 118620 140856 122531 140858
rect 118620 140800 122470 140856
rect 122526 140800 122531 140856
rect 118620 140798 122531 140800
rect 118620 140796 118626 140798
rect 122465 140795 122531 140798
rect 124213 140858 124279 140861
rect 124673 140858 124739 140861
rect 580441 140858 580507 140861
rect 124213 140856 580507 140858
rect 124213 140800 124218 140856
rect 124274 140800 124678 140856
rect 124734 140800 580446 140856
rect 580502 140800 580507 140856
rect 124213 140798 580507 140800
rect 124213 140795 124279 140798
rect 124673 140795 124739 140798
rect 580441 140795 580507 140798
rect 193438 140660 193444 140724
rect 193508 140722 193514 140724
rect 193673 140722 193739 140725
rect 193508 140720 193739 140722
rect 193508 140664 193678 140720
rect 193734 140664 193739 140720
rect 193508 140662 193739 140664
rect 193508 140660 193514 140662
rect 193673 140659 193739 140662
rect 120022 140524 120028 140588
rect 120092 140586 120098 140588
rect 126329 140586 126395 140589
rect 120092 140584 126395 140586
rect 120092 140528 126334 140584
rect 126390 140528 126395 140584
rect 120092 140526 126395 140528
rect 120092 140524 120098 140526
rect 126329 140523 126395 140526
rect 181437 140450 181503 140453
rect 188286 140450 188292 140452
rect 181437 140448 188292 140450
rect 181437 140392 181442 140448
rect 181498 140392 188292 140448
rect 181437 140390 188292 140392
rect 181437 140387 181503 140390
rect 188286 140388 188292 140390
rect 188356 140388 188362 140452
rect 117998 140252 118004 140316
rect 118068 140314 118074 140316
rect 127617 140314 127683 140317
rect 118068 140312 127683 140314
rect 118068 140256 127622 140312
rect 127678 140256 127683 140312
rect 118068 140254 127683 140256
rect 118068 140252 118074 140254
rect 127617 140251 127683 140254
rect 130326 140252 130332 140316
rect 130396 140314 130402 140316
rect 130469 140314 130535 140317
rect 130396 140312 130535 140314
rect 130396 140256 130474 140312
rect 130530 140256 130535 140312
rect 130396 140254 130535 140256
rect 130396 140252 130402 140254
rect 130469 140251 130535 140254
rect 182817 140314 182883 140317
rect 190678 140314 190684 140316
rect 182817 140312 190684 140314
rect 182817 140256 182822 140312
rect 182878 140256 190684 140312
rect 182817 140254 190684 140256
rect 182817 140251 182883 140254
rect 190678 140252 190684 140254
rect 190748 140252 190754 140316
rect 120758 140116 120764 140180
rect 120828 140178 120834 140180
rect 154021 140178 154087 140181
rect 120828 140176 154087 140178
rect 120828 140120 154026 140176
rect 154082 140120 154087 140176
rect 120828 140118 154087 140120
rect 120828 140116 120834 140118
rect 154021 140115 154087 140118
rect 178769 140178 178835 140181
rect 194542 140178 194548 140180
rect 178769 140176 194548 140178
rect 178769 140120 178774 140176
rect 178830 140120 194548 140176
rect 178769 140118 194548 140120
rect 178769 140115 178835 140118
rect 194542 140116 194548 140118
rect 194612 140116 194618 140180
rect 109534 139980 109540 140044
rect 109604 140042 109610 140044
rect 131665 140042 131731 140045
rect 109604 140040 131731 140042
rect 109604 139984 131670 140040
rect 131726 139984 131731 140040
rect 109604 139982 131731 139984
rect 109604 139980 109610 139982
rect 131665 139979 131731 139982
rect 151486 139980 151492 140044
rect 151556 140042 151562 140044
rect 194041 140042 194107 140045
rect 151556 140040 194107 140042
rect 151556 139984 194046 140040
rect 194102 139984 194107 140040
rect 151556 139982 194107 139984
rect 151556 139980 151562 139982
rect 194041 139979 194107 139982
rect 185485 139906 185551 139909
rect 190494 139906 190500 139908
rect 185485 139904 190500 139906
rect 185485 139848 185490 139904
rect 185546 139848 190500 139904
rect 185485 139846 190500 139848
rect 185485 139843 185551 139846
rect 190494 139844 190500 139846
rect 190564 139844 190570 139908
rect 113766 139708 113772 139772
rect 113836 139770 113842 139772
rect 122373 139770 122439 139773
rect 113836 139768 122439 139770
rect 113836 139712 122378 139768
rect 122434 139712 122439 139768
rect 113836 139710 122439 139712
rect 113836 139708 113842 139710
rect 122373 139707 122439 139710
rect 185761 139770 185827 139773
rect 192150 139770 192156 139772
rect 185761 139768 192156 139770
rect 185761 139712 185766 139768
rect 185822 139712 192156 139768
rect 185761 139710 192156 139712
rect 185761 139707 185827 139710
rect 192150 139708 192156 139710
rect 192220 139708 192226 139772
rect 116710 139572 116716 139636
rect 116780 139634 116786 139636
rect 182633 139634 182699 139637
rect 185393 139634 185459 139637
rect 116780 139632 182699 139634
rect 116780 139576 182638 139632
rect 182694 139576 182699 139632
rect 116780 139574 182699 139576
rect 116780 139572 116786 139574
rect 182633 139571 182699 139574
rect 182774 139632 185459 139634
rect 182774 139576 185398 139632
rect 185454 139576 185459 139632
rect 182774 139574 185459 139576
rect 17217 139498 17283 139501
rect 182774 139498 182834 139574
rect 185393 139571 185459 139574
rect 17217 139496 182834 139498
rect 17217 139440 17222 139496
rect 17278 139440 182834 139496
rect 17217 139438 182834 139440
rect 183001 139498 183067 139501
rect 189390 139498 189396 139500
rect 183001 139496 189396 139498
rect 183001 139440 183006 139496
rect 183062 139440 189396 139496
rect 183001 139438 189396 139440
rect 17217 139435 17283 139438
rect 183001 139435 183067 139438
rect 189390 139436 189396 139438
rect 189460 139436 189466 139500
rect 112345 139362 112411 139365
rect 126237 139362 126303 139365
rect 130561 139362 130627 139365
rect 149421 139362 149487 139365
rect 112345 139360 126303 139362
rect 112345 139304 112350 139360
rect 112406 139304 126242 139360
rect 126298 139304 126303 139360
rect 112345 139302 126303 139304
rect 112345 139299 112411 139302
rect 126237 139299 126303 139302
rect 126838 139360 130627 139362
rect 126838 139304 130566 139360
rect 130622 139304 130627 139360
rect 126838 139302 130627 139304
rect 115197 139226 115263 139229
rect 126838 139226 126898 139302
rect 130561 139299 130627 139302
rect 142110 139360 149487 139362
rect 142110 139304 149426 139360
rect 149482 139304 149487 139360
rect 142110 139302 149487 139304
rect 115197 139224 126898 139226
rect 115197 139168 115202 139224
rect 115258 139168 126898 139224
rect 115197 139166 126898 139168
rect 115197 139163 115263 139166
rect 114134 139028 114140 139092
rect 114204 139090 114210 139092
rect 130326 139090 130332 139092
rect 114204 139030 130332 139090
rect 114204 139028 114210 139030
rect 130326 139028 130332 139030
rect 130396 139028 130402 139092
rect 106825 138954 106891 138957
rect 113173 138954 113239 138957
rect 106825 138952 113239 138954
rect 106825 138896 106830 138952
rect 106886 138896 113178 138952
rect 113234 138896 113239 138952
rect 106825 138894 113239 138896
rect 106825 138891 106891 138894
rect 113173 138891 113239 138894
rect 102593 138818 102659 138821
rect 122097 138818 122163 138821
rect 102593 138816 122163 138818
rect 102593 138760 102598 138816
rect 102654 138760 122102 138816
rect 122158 138760 122163 138816
rect 102593 138758 122163 138760
rect 102593 138755 102659 138758
rect 122097 138755 122163 138758
rect 122741 138818 122807 138821
rect 123937 138818 124003 138821
rect 122741 138816 124003 138818
rect 122741 138760 122746 138816
rect 122802 138760 123942 138816
rect 123998 138760 124003 138816
rect 122741 138758 124003 138760
rect 122741 138755 122807 138758
rect 123937 138755 124003 138758
rect 101213 138682 101279 138685
rect 142110 138682 142170 139302
rect 149421 139299 149487 139302
rect 174997 139362 175063 139365
rect 184105 139362 184171 139365
rect 184381 139362 184447 139365
rect 185945 139362 186011 139365
rect 174997 139360 180810 139362
rect 174997 139304 175002 139360
rect 175058 139304 180810 139360
rect 174997 139302 180810 139304
rect 174997 139299 175063 139302
rect 101213 138680 142170 138682
rect 101213 138624 101218 138680
rect 101274 138624 142170 138680
rect 101213 138622 142170 138624
rect 180750 138682 180810 139302
rect 184105 139360 184306 139362
rect 184105 139304 184110 139360
rect 184166 139304 184306 139360
rect 184105 139302 184306 139304
rect 184105 139299 184171 139302
rect 184246 138818 184306 139302
rect 184381 139360 184490 139362
rect 184381 139304 184386 139360
rect 184442 139304 184490 139360
rect 184381 139299 184490 139304
rect 184430 139226 184490 139299
rect 185902 139360 186011 139362
rect 185902 139304 185950 139360
rect 186006 139304 186011 139360
rect 185902 139299 186011 139304
rect 186497 139362 186563 139365
rect 187049 139362 187115 139365
rect 193857 139362 193923 139365
rect 186497 139360 186698 139362
rect 186497 139304 186502 139360
rect 186558 139304 186698 139360
rect 186497 139302 186698 139304
rect 186497 139299 186563 139302
rect 184430 139166 184674 139226
rect 184614 138954 184674 139166
rect 185902 139090 185962 139299
rect 186638 139226 186698 139302
rect 187049 139360 193923 139362
rect 187049 139304 187054 139360
rect 187110 139304 193862 139360
rect 193918 139304 193923 139360
rect 187049 139302 193923 139304
rect 187049 139299 187115 139302
rect 193857 139299 193923 139302
rect 579797 139362 579863 139365
rect 583520 139362 584960 139452
rect 579797 139360 584960 139362
rect 579797 139304 579802 139360
rect 579858 139304 584960 139360
rect 579797 139302 584960 139304
rect 579797 139299 579863 139302
rect 195237 139226 195303 139229
rect 186638 139224 195303 139226
rect 186638 139168 195242 139224
rect 195298 139168 195303 139224
rect 583520 139212 584960 139302
rect 186638 139166 195303 139168
rect 195237 139163 195303 139166
rect 199101 139090 199167 139093
rect 185902 139088 199167 139090
rect 185902 139032 199106 139088
rect 199162 139032 199167 139088
rect 185902 139030 199167 139032
rect 199101 139027 199167 139030
rect 197813 138954 197879 138957
rect 184614 138952 197879 138954
rect 184614 138896 197818 138952
rect 197874 138896 197879 138952
rect 184614 138894 197879 138896
rect 197813 138891 197879 138894
rect 199561 138818 199627 138821
rect 184246 138816 199627 138818
rect 184246 138760 199566 138816
rect 199622 138760 199627 138816
rect 184246 138758 199627 138760
rect 199561 138755 199627 138758
rect 196617 138682 196683 138685
rect 180750 138680 196683 138682
rect 180750 138624 196622 138680
rect 196678 138624 196683 138680
rect 180750 138622 196683 138624
rect 101213 138619 101279 138622
rect 196617 138619 196683 138622
rect 112529 138546 112595 138549
rect 122281 138546 122347 138549
rect 112529 138544 122347 138546
rect 112529 138488 112534 138544
rect 112590 138488 122286 138544
rect 122342 138488 122347 138544
rect 112529 138486 122347 138488
rect 112529 138483 112595 138486
rect 122281 138483 122347 138486
rect 113173 138410 113239 138413
rect 123569 138410 123635 138413
rect 113173 138408 123635 138410
rect 113173 138352 113178 138408
rect 113234 138352 123574 138408
rect 123630 138352 123635 138408
rect 113173 138350 123635 138352
rect 113173 138347 113239 138350
rect 123569 138347 123635 138350
rect 120809 138138 120875 138141
rect 121126 138138 121132 138140
rect 120809 138136 121132 138138
rect 120809 138080 120814 138136
rect 120870 138080 121132 138136
rect 120809 138078 121132 138080
rect 120809 138075 120875 138078
rect 121126 138076 121132 138078
rect 121196 138076 121202 138140
rect 123150 138076 123156 138140
rect 123220 138138 123226 138140
rect 124029 138138 124095 138141
rect 123220 138136 124095 138138
rect 123220 138080 124034 138136
rect 124090 138080 124095 138136
rect 123220 138078 124095 138080
rect 123220 138076 123226 138078
rect 124029 138075 124095 138078
rect 194501 138138 194567 138141
rect 198958 138138 198964 138140
rect 194501 138136 198964 138138
rect 194501 138080 194506 138136
rect 194562 138080 198964 138136
rect 194501 138078 198964 138080
rect 194501 138075 194567 138078
rect 198958 138076 198964 138078
rect 199028 138076 199034 138140
rect 122741 138004 122807 138005
rect 122741 138000 122788 138004
rect 122852 138002 122858 138004
rect 122741 137944 122746 138000
rect 122741 137940 122788 137944
rect 122852 137942 122898 138002
rect 122852 137940 122858 137942
rect 187918 137940 187924 138004
rect 187988 138002 187994 138004
rect 188889 138002 188955 138005
rect 187988 138000 188955 138002
rect 187988 137944 188894 138000
rect 188950 137944 188955 138000
rect 187988 137942 188955 137944
rect 187988 137940 187994 137942
rect 122741 137939 122807 137940
rect 188889 137939 188955 137942
rect 119153 137866 119219 137869
rect 124806 137866 124812 137868
rect 119153 137864 124812 137866
rect 119153 137808 119158 137864
rect 119214 137808 124812 137864
rect 119153 137806 124812 137808
rect 119153 137803 119219 137806
rect 124806 137804 124812 137806
rect 124876 137804 124882 137868
rect 187182 137804 187188 137868
rect 187252 137866 187258 137868
rect 188153 137866 188219 137869
rect 187252 137864 188219 137866
rect 187252 137808 188158 137864
rect 188214 137808 188219 137864
rect 187252 137806 188219 137808
rect 187252 137804 187258 137806
rect 188153 137803 188219 137806
rect 188286 137804 188292 137868
rect 188356 137866 188362 137868
rect 200941 137866 201007 137869
rect 188356 137864 201007 137866
rect 188356 137808 200946 137864
rect 201002 137808 201007 137864
rect 188356 137806 201007 137808
rect 188356 137804 188362 137806
rect 200941 137803 201007 137806
rect 105118 137260 105124 137324
rect 105188 137322 105194 137324
rect 120574 137322 120580 137324
rect 105188 137262 120580 137322
rect 105188 137260 105194 137262
rect 120574 137260 120580 137262
rect 120644 137260 120650 137324
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 119654 130324 119660 130388
rect 119724 130386 119730 130388
rect 120022 130386 120028 130388
rect 119724 130326 120028 130386
rect 119724 130324 119730 130326
rect 120022 130324 120028 130326
rect 120092 130324 120098 130388
rect 122741 128484 122807 128485
rect 122741 128482 122788 128484
rect 122696 128480 122788 128482
rect 122696 128424 122746 128480
rect 122696 128422 122788 128424
rect 122741 128420 122788 128422
rect 122852 128420 122858 128484
rect 122741 128419 122807 128420
rect 580809 126034 580875 126037
rect 583520 126034 584960 126124
rect 580809 126032 584960 126034
rect 580809 125976 580814 126032
rect 580870 125976 584960 126032
rect 580809 125974 584960 125976
rect 580809 125971 580875 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 109493 123450 109559 123453
rect 123150 123450 123156 123452
rect 109493 123448 123156 123450
rect 109493 123392 109498 123448
rect 109554 123392 123156 123448
rect 109493 123390 123156 123392
rect 109493 123387 109559 123390
rect 123150 123388 123156 123390
rect 123220 123388 123226 123452
rect 122782 122980 122788 123044
rect 122852 122980 122858 123044
rect 122790 122909 122850 122980
rect 122741 122906 122850 122909
rect 122696 122904 122850 122906
rect 122696 122848 122746 122904
rect 122802 122848 122850 122904
rect 122696 122846 122850 122848
rect 122741 122843 122807 122846
rect 122230 122164 122236 122228
rect 122300 122226 122306 122228
rect 122598 122226 122604 122228
rect 122300 122166 122604 122226
rect 122300 122164 122306 122166
rect 122598 122164 122604 122166
rect 122668 122164 122674 122228
rect 191598 114412 191604 114476
rect 191668 114474 191674 114476
rect 198089 114474 198155 114477
rect 191668 114472 198155 114474
rect 191668 114416 198094 114472
rect 198150 114416 198155 114472
rect 191668 114414 198155 114416
rect 191668 114412 191674 114414
rect 198089 114411 198155 114414
rect 189574 113868 189580 113932
rect 189644 113930 189650 113932
rect 196801 113930 196867 113933
rect 189644 113928 196867 113930
rect 189644 113872 196806 113928
rect 196862 113872 196867 113928
rect 189644 113870 196867 113872
rect 189644 113868 189650 113870
rect 196801 113867 196867 113870
rect 103973 113794 104039 113797
rect 115238 113794 115244 113796
rect 103973 113792 115244 113794
rect 103973 113736 103978 113792
rect 104034 113736 115244 113792
rect 103973 113734 115244 113736
rect 103973 113731 104039 113734
rect 115238 113732 115244 113734
rect 115308 113732 115314 113796
rect 122230 113732 122236 113796
rect 122300 113794 122306 113796
rect 122598 113794 122604 113796
rect 122300 113734 122604 113794
rect 122300 113732 122306 113734
rect 122598 113732 122604 113734
rect 122668 113732 122674 113796
rect 189390 113324 189396 113388
rect 189460 113386 189466 113388
rect 189574 113386 189580 113388
rect 189460 113326 189580 113386
rect 189460 113324 189466 113326
rect 189574 113324 189580 113326
rect 189644 113324 189650 113388
rect 580717 112842 580783 112845
rect 583520 112842 584960 112932
rect 580717 112840 584960 112842
rect 580717 112784 580722 112840
rect 580778 112784 584960 112840
rect 580717 112782 584960 112784
rect 580717 112779 580783 112782
rect 122230 112644 122236 112708
rect 122300 112706 122306 112708
rect 122598 112706 122604 112708
rect 122300 112646 122604 112706
rect 122300 112644 122306 112646
rect 122598 112644 122604 112646
rect 122668 112644 122674 112708
rect 583520 112692 584960 112782
rect 102685 112434 102751 112437
rect 119470 112434 119476 112436
rect 102685 112432 119476 112434
rect 102685 112376 102690 112432
rect 102746 112376 119476 112432
rect 102685 112374 119476 112376
rect 102685 112371 102751 112374
rect 119470 112372 119476 112374
rect 119540 112372 119546 112436
rect 119470 111828 119476 111892
rect 119540 111890 119546 111892
rect 122046 111890 122052 111892
rect 119540 111830 122052 111890
rect 119540 111828 119546 111830
rect 122046 111828 122052 111830
rect 122116 111828 122122 111892
rect -960 110666 480 110756
rect 2773 110666 2839 110669
rect -960 110664 2839 110666
rect -960 110608 2778 110664
rect 2834 110608 2839 110664
rect -960 110606 2839 110608
rect -960 110516 480 110606
rect 2773 110603 2839 110606
rect 115013 110666 115079 110669
rect 122046 110666 122052 110668
rect 115013 110664 122052 110666
rect 115013 110608 115018 110664
rect 115074 110608 122052 110664
rect 115013 110606 122052 110608
rect 115013 110603 115079 110606
rect 122046 110604 122052 110606
rect 122116 110604 122122 110668
rect 189390 110604 189396 110668
rect 189460 110666 189466 110668
rect 189533 110666 189599 110669
rect 189460 110664 189599 110666
rect 189460 110608 189538 110664
rect 189594 110608 189599 110664
rect 189460 110606 189599 110608
rect 189460 110604 189466 110606
rect 189533 110603 189599 110606
rect 113582 110468 113588 110532
rect 113652 110530 113658 110532
rect 120758 110530 120764 110532
rect 113652 110470 120764 110530
rect 113652 110468 113658 110470
rect 120758 110468 120764 110470
rect 120828 110468 120834 110532
rect 189390 109244 189396 109308
rect 189460 109306 189466 109308
rect 189460 109246 190470 109306
rect 189460 109244 189466 109246
rect 190410 109170 190470 109246
rect 191281 109170 191347 109173
rect 190410 109168 191347 109170
rect 190410 109112 191286 109168
rect 191342 109112 191347 109168
rect 190410 109110 191347 109112
rect 191281 109107 191347 109110
rect 189390 107068 189396 107132
rect 189460 107130 189466 107132
rect 189533 107130 189599 107133
rect 189460 107128 189599 107130
rect 189460 107072 189538 107128
rect 189594 107072 189599 107128
rect 189460 107070 189599 107072
rect 189460 107068 189466 107070
rect 189533 107067 189599 107070
rect 122230 103532 122236 103596
rect 122300 103594 122306 103596
rect 122598 103594 122604 103596
rect 122300 103534 122604 103594
rect 122300 103532 122306 103534
rect 122598 103532 122604 103534
rect 122668 103532 122674 103596
rect 122230 103124 122236 103188
rect 122300 103186 122306 103188
rect 122598 103186 122604 103188
rect 122300 103126 122604 103186
rect 122300 103124 122306 103126
rect 122598 103124 122604 103126
rect 122668 103124 122674 103188
rect 579613 99514 579679 99517
rect 583520 99514 584960 99604
rect 579613 99512 584960 99514
rect 579613 99456 579618 99512
rect 579674 99456 584960 99512
rect 579613 99454 584960 99456
rect 579613 99451 579679 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect -960 97550 674 97610
rect -960 97474 480 97550
rect 614 97474 674 97550
rect -960 97460 674 97474
rect 246 97414 674 97460
rect 246 96930 306 97414
rect 246 96870 6930 96930
rect 6870 96658 6930 96870
rect 116710 96658 116716 96660
rect 6870 96598 116716 96658
rect 116710 96596 116716 96598
rect 116780 96596 116786 96660
rect 122230 94012 122236 94076
rect 122300 94074 122306 94076
rect 122598 94074 122604 94076
rect 122300 94014 122604 94074
rect 122300 94012 122306 94014
rect 122598 94012 122604 94014
rect 122668 94012 122674 94076
rect 122230 93604 122236 93668
rect 122300 93666 122306 93668
rect 122598 93666 122604 93668
rect 122300 93606 122604 93666
rect 122300 93604 122306 93606
rect 122598 93604 122604 93606
rect 122668 93604 122674 93668
rect 579613 86186 579679 86189
rect 583520 86186 584960 86276
rect 579613 86184 584960 86186
rect 579613 86128 579618 86184
rect 579674 86128 584960 86184
rect 579613 86126 584960 86128
rect 579613 86123 579679 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 122230 84492 122236 84556
rect 122300 84554 122306 84556
rect 122598 84554 122604 84556
rect 122300 84494 122604 84554
rect 122300 84492 122306 84494
rect 122598 84492 122604 84494
rect 122668 84492 122674 84556
rect 122741 84146 122807 84149
rect 122696 84144 122850 84146
rect 122696 84088 122746 84144
rect 122802 84088 122850 84144
rect 122696 84086 122850 84088
rect 122741 84083 122850 84086
rect 122790 84012 122850 84083
rect 122782 83948 122788 84012
rect 122852 83948 122858 84012
rect 196157 82242 196223 82245
rect 196382 82242 196388 82244
rect 196157 82240 196388 82242
rect 196157 82184 196162 82240
rect 196218 82184 196388 82240
rect 196157 82182 196388 82184
rect 196157 82179 196223 82182
rect 196382 82180 196388 82182
rect 196452 82180 196458 82244
rect 191598 81500 191604 81564
rect 191668 81562 191674 81564
rect 199469 81562 199535 81565
rect 191668 81560 199535 81562
rect 191668 81504 199474 81560
rect 199530 81504 199535 81560
rect 191668 81502 199535 81504
rect 191668 81500 191674 81502
rect 199469 81499 199535 81502
rect 105169 81428 105235 81429
rect 105118 81426 105124 81428
rect 105078 81366 105124 81426
rect 105188 81424 105235 81428
rect 105230 81368 105235 81424
rect 105118 81364 105124 81366
rect 105188 81364 105235 81368
rect 105169 81363 105235 81364
rect 124070 81228 124076 81292
rect 124140 81290 124146 81292
rect 147806 81290 147812 81292
rect 124140 81230 147812 81290
rect 124140 81228 124146 81230
rect 147806 81228 147812 81230
rect 147876 81228 147882 81292
rect 163998 81228 164004 81292
rect 164068 81290 164074 81292
rect 191966 81290 191972 81292
rect 164068 81230 191972 81290
rect 164068 81228 164074 81230
rect 191966 81228 191972 81230
rect 192036 81228 192042 81292
rect 103973 81154 104039 81157
rect 124029 81154 124095 81157
rect 103973 81152 124095 81154
rect 103973 81096 103978 81152
rect 104034 81096 124034 81152
rect 124090 81096 124095 81152
rect 103973 81094 124095 81096
rect 103973 81091 104039 81094
rect 124029 81091 124095 81094
rect 175406 81092 175412 81156
rect 175476 81154 175482 81156
rect 207841 81154 207907 81157
rect 175476 81152 207907 81154
rect 175476 81096 207846 81152
rect 207902 81096 207907 81152
rect 175476 81094 207907 81096
rect 175476 81092 175482 81094
rect 207841 81091 207907 81094
rect 117773 81018 117839 81021
rect 151302 81018 151308 81020
rect 117773 81016 151308 81018
rect 117773 80960 117778 81016
rect 117834 80960 151308 81016
rect 117773 80958 151308 80960
rect 117773 80955 117839 80958
rect 151302 80956 151308 80958
rect 151372 80956 151378 81020
rect 174302 80956 174308 81020
rect 174372 81018 174378 81020
rect 207749 81018 207815 81021
rect 174372 81016 207815 81018
rect 174372 80960 207754 81016
rect 207810 80960 207815 81016
rect 174372 80958 207815 80960
rect 174372 80956 174378 80958
rect 207749 80955 207815 80958
rect 113817 80882 113883 80885
rect 148910 80882 148916 80884
rect 113817 80880 148916 80882
rect 113817 80824 113822 80880
rect 113878 80824 148916 80880
rect 113817 80822 148916 80824
rect 113817 80819 113883 80822
rect 148910 80820 148916 80822
rect 148980 80820 148986 80884
rect 172278 80820 172284 80884
rect 172348 80882 172354 80884
rect 204989 80882 205055 80885
rect 172348 80880 205055 80882
rect 172348 80824 204994 80880
rect 205050 80824 205055 80880
rect 172348 80822 205055 80824
rect 172348 80820 172354 80822
rect 204989 80819 205055 80822
rect 112253 80746 112319 80749
rect 146334 80746 146340 80748
rect 112253 80744 146340 80746
rect 112253 80688 112258 80744
rect 112314 80688 146340 80744
rect 112253 80686 146340 80688
rect 112253 80683 112319 80686
rect 146334 80684 146340 80686
rect 146404 80684 146410 80748
rect 181662 80684 181668 80748
rect 181732 80746 181738 80748
rect 206369 80746 206435 80749
rect 181732 80744 206435 80746
rect 181732 80688 206374 80744
rect 206430 80688 206435 80744
rect 181732 80686 206435 80688
rect 181732 80684 181738 80686
rect 206369 80683 206435 80686
rect 120073 80610 120139 80613
rect 122189 80610 122255 80613
rect 120073 80608 122255 80610
rect 120073 80552 120078 80608
rect 120134 80552 122194 80608
rect 122250 80552 122255 80608
rect 120073 80550 122255 80552
rect 120073 80547 120139 80550
rect 122189 80547 122255 80550
rect 124029 80610 124095 80613
rect 128997 80610 129063 80613
rect 124029 80608 129063 80610
rect 124029 80552 124034 80608
rect 124090 80552 129002 80608
rect 129058 80552 129063 80608
rect 124029 80550 129063 80552
rect 124029 80547 124095 80550
rect 128997 80547 129063 80550
rect 181621 80610 181687 80613
rect 197670 80610 197676 80612
rect 181621 80608 197676 80610
rect 181621 80552 181626 80608
rect 181682 80552 197676 80608
rect 181621 80550 197676 80552
rect 181621 80547 181687 80550
rect 197670 80548 197676 80550
rect 197740 80548 197746 80612
rect 113950 80412 113956 80476
rect 114020 80474 114026 80476
rect 120625 80474 120691 80477
rect 114020 80472 120691 80474
rect 114020 80416 120630 80472
rect 120686 80416 120691 80472
rect 114020 80414 120691 80416
rect 114020 80412 114026 80414
rect 120625 80411 120691 80414
rect 173014 80412 173020 80476
rect 173084 80474 173090 80476
rect 178217 80474 178283 80477
rect 173084 80472 178283 80474
rect 173084 80416 178222 80472
rect 178278 80416 178283 80472
rect 173084 80414 178283 80416
rect 173084 80412 173090 80414
rect 178217 80411 178283 80414
rect 178401 80474 178467 80477
rect 193438 80474 193444 80476
rect 178401 80472 193444 80474
rect 178401 80416 178406 80472
rect 178462 80416 193444 80472
rect 178401 80414 193444 80416
rect 178401 80411 178467 80414
rect 193438 80412 193444 80414
rect 193508 80412 193514 80476
rect 108246 80276 108252 80340
rect 108316 80338 108322 80340
rect 181621 80338 181687 80341
rect 108316 80278 136466 80338
rect 108316 80276 108322 80278
rect 119153 80202 119219 80205
rect 122373 80202 122439 80205
rect 119153 80200 122439 80202
rect 119153 80144 119158 80200
rect 119214 80144 122378 80200
rect 122434 80144 122439 80200
rect 119153 80142 122439 80144
rect 119153 80139 119219 80142
rect 122373 80139 122439 80142
rect 130285 80202 130351 80205
rect 130285 80200 135086 80202
rect 130285 80144 130290 80200
rect 130346 80144 135086 80200
rect 130285 80142 135086 80144
rect 130285 80139 130351 80142
rect 135026 79967 135086 80142
rect 135302 80142 136282 80202
rect 135302 80068 135362 80142
rect 135294 80004 135300 80068
rect 135364 80004 135370 80068
rect 132907 79962 132973 79967
rect 128261 79930 128327 79933
rect 132539 79930 132605 79933
rect 128261 79928 132605 79930
rect 128261 79872 128266 79928
rect 128322 79872 132544 79928
rect 132600 79872 132605 79928
rect 132907 79906 132912 79962
rect 132968 79906 132973 79962
rect 132907 79901 132973 79906
rect 133551 79962 133617 79967
rect 133551 79906 133556 79962
rect 133612 79906 133617 79962
rect 133551 79901 133617 79906
rect 133735 79964 133801 79967
rect 133735 79962 133844 79964
rect 133735 79906 133740 79962
rect 133796 79906 133844 79962
rect 133735 79901 133844 79906
rect 134011 79962 134077 79967
rect 134011 79906 134016 79962
rect 134072 79906 134077 79962
rect 134195 79962 134261 79967
rect 134195 79932 134200 79962
rect 134256 79932 134261 79962
rect 134563 79962 134629 79967
rect 134563 79932 134568 79962
rect 134624 79932 134629 79962
rect 135023 79962 135089 79967
rect 134011 79901 134077 79906
rect 128261 79870 132605 79872
rect 128261 79867 128327 79870
rect 132539 79867 132605 79870
rect 132910 79797 132970 79901
rect 132309 79794 132375 79797
rect 132309 79792 132510 79794
rect 132309 79736 132314 79792
rect 132370 79736 132510 79792
rect 132309 79734 132510 79736
rect 132910 79792 133019 79797
rect 132910 79736 132958 79792
rect 133014 79736 133019 79792
rect 132910 79734 133019 79736
rect 132309 79731 132375 79734
rect 132450 79658 132510 79734
rect 132953 79731 133019 79734
rect 133321 79794 133387 79797
rect 133554 79794 133614 79901
rect 133784 79797 133844 79901
rect 133321 79792 133614 79794
rect 133321 79736 133326 79792
rect 133382 79736 133614 79792
rect 133321 79734 133614 79736
rect 133735 79792 133844 79797
rect 133735 79736 133740 79792
rect 133796 79736 133844 79792
rect 133735 79734 133844 79736
rect 134014 79794 134074 79901
rect 134190 79868 134196 79932
rect 134260 79930 134266 79932
rect 134260 79870 134318 79930
rect 134260 79868 134266 79870
rect 134558 79868 134564 79932
rect 134628 79930 134634 79932
rect 134628 79870 134686 79930
rect 135023 79906 135028 79962
rect 135084 79906 135089 79962
rect 135023 79901 135089 79906
rect 135299 79928 135365 79933
rect 135299 79872 135304 79928
rect 135360 79872 135365 79928
rect 134628 79868 134634 79870
rect 135299 79867 135365 79872
rect 135575 79930 135641 79933
rect 135846 79930 135852 79932
rect 135575 79928 135852 79930
rect 135575 79872 135580 79928
rect 135636 79872 135852 79928
rect 135575 79870 135852 79872
rect 135575 79867 135641 79870
rect 135846 79868 135852 79870
rect 135916 79868 135922 79932
rect 136222 79899 136282 80142
rect 136219 79894 136285 79899
rect 134149 79794 134215 79797
rect 134014 79792 134215 79794
rect 134014 79736 134154 79792
rect 134210 79736 134215 79792
rect 134014 79734 134215 79736
rect 135302 79794 135362 79867
rect 136219 79838 136224 79894
rect 136280 79838 136285 79894
rect 136219 79833 136285 79838
rect 135662 79794 135668 79796
rect 135302 79734 135668 79794
rect 133321 79731 133387 79734
rect 133735 79731 133801 79734
rect 134149 79731 134215 79734
rect 135662 79732 135668 79734
rect 135732 79732 135738 79796
rect 136406 79794 136466 80278
rect 174080 80336 181687 80338
rect 174080 80280 181626 80336
rect 181682 80280 181687 80336
rect 174080 80278 181687 80280
rect 139342 80140 139348 80204
rect 139412 80202 139418 80204
rect 139412 80142 140422 80202
rect 139412 80140 139418 80142
rect 136955 79962 137021 79967
rect 139071 79964 139137 79967
rect 136955 79932 136960 79962
rect 137016 79932 137021 79962
rect 139028 79962 139137 79964
rect 136950 79868 136956 79932
rect 137020 79930 137026 79932
rect 137020 79870 137078 79930
rect 137139 79928 137205 79933
rect 137139 79872 137144 79928
rect 137200 79872 137205 79928
rect 137020 79868 137026 79870
rect 137139 79867 137205 79872
rect 137507 79928 137573 79933
rect 137875 79932 137941 79933
rect 138611 79932 138677 79933
rect 139028 79932 139076 79962
rect 137870 79930 137876 79932
rect 137507 79872 137512 79928
rect 137568 79872 137573 79928
rect 137507 79867 137573 79872
rect 137784 79870 137876 79930
rect 137870 79868 137876 79870
rect 137940 79868 137946 79932
rect 138606 79930 138612 79932
rect 138520 79870 138612 79930
rect 138606 79868 138612 79870
rect 138676 79868 138682 79932
rect 138974 79868 138980 79932
rect 139044 79906 139076 79932
rect 139132 79906 139137 79962
rect 140362 79933 140422 80142
rect 143390 80140 143396 80204
rect 143460 80202 143466 80204
rect 143460 80142 144056 80202
rect 143460 80140 143466 80142
rect 143996 79967 144056 80142
rect 147070 80140 147076 80204
rect 147140 80202 147146 80204
rect 158110 80202 158116 80204
rect 147140 80142 147506 80202
rect 147140 80140 147146 80142
rect 147446 79967 147506 80142
rect 157566 80142 158116 80202
rect 151670 80066 151676 80068
rect 151632 80004 151676 80066
rect 151740 80004 151746 80068
rect 141463 79962 141529 79967
rect 139044 79901 139137 79906
rect 139531 79930 139597 79933
rect 139899 79932 139965 79933
rect 139710 79930 139716 79932
rect 139531 79928 139716 79930
rect 139044 79870 139088 79901
rect 139531 79872 139536 79928
rect 139592 79872 139716 79928
rect 139531 79870 139716 79872
rect 139044 79868 139050 79870
rect 137875 79867 137941 79868
rect 138611 79867 138677 79868
rect 139531 79867 139597 79870
rect 139710 79868 139716 79870
rect 139780 79868 139786 79932
rect 139894 79868 139900 79932
rect 139964 79930 139970 79932
rect 139964 79870 140056 79930
rect 140359 79928 140425 79933
rect 140359 79872 140364 79928
rect 140420 79872 140425 79928
rect 139964 79868 139970 79870
rect 139899 79867 139965 79868
rect 140359 79867 140425 79872
rect 140630 79868 140636 79932
rect 140700 79930 140706 79932
rect 140911 79930 140977 79933
rect 140700 79928 140977 79930
rect 140700 79872 140916 79928
rect 140972 79872 140977 79928
rect 140700 79870 140977 79872
rect 140700 79868 140706 79870
rect 140911 79867 140977 79870
rect 141182 79868 141188 79932
rect 141252 79930 141258 79932
rect 141463 79930 141468 79962
rect 141252 79906 141468 79930
rect 141524 79906 141529 79962
rect 142291 79962 142357 79967
rect 142291 79932 142296 79962
rect 142352 79932 142357 79962
rect 142659 79962 142725 79967
rect 142659 79932 142664 79962
rect 142720 79932 142725 79962
rect 142843 79962 142909 79967
rect 143303 79964 143369 79967
rect 141252 79901 141529 79906
rect 141252 79870 141526 79901
rect 141252 79868 141258 79870
rect 142286 79868 142292 79932
rect 142356 79930 142362 79932
rect 142356 79870 142414 79930
rect 142356 79868 142362 79870
rect 142654 79868 142660 79932
rect 142724 79930 142730 79932
rect 142724 79870 142782 79930
rect 142843 79906 142848 79962
rect 142904 79930 142909 79962
rect 143260 79962 143369 79964
rect 143260 79932 143308 79962
rect 143022 79930 143028 79932
rect 142904 79906 143028 79930
rect 142843 79901 143028 79906
rect 142846 79870 143028 79901
rect 142724 79868 142730 79870
rect 143022 79868 143028 79870
rect 143092 79868 143098 79932
rect 143206 79868 143212 79932
rect 143276 79906 143308 79932
rect 143364 79906 143369 79962
rect 143763 79964 143829 79967
rect 143763 79962 143886 79964
rect 143763 79932 143768 79962
rect 143824 79932 143886 79962
rect 143276 79901 143369 79906
rect 143276 79870 143320 79901
rect 143276 79868 143282 79870
rect 143758 79868 143764 79932
rect 143828 79904 143886 79932
rect 143996 79962 144105 79967
rect 143996 79906 144044 79962
rect 144100 79906 144105 79962
rect 143996 79904 144105 79906
rect 143828 79868 143834 79904
rect 144039 79901 144105 79904
rect 144223 79964 144289 79967
rect 144223 79962 144332 79964
rect 144223 79906 144228 79962
rect 144284 79932 144332 79962
rect 145051 79962 145117 79967
rect 145695 79964 145761 79967
rect 144683 79932 144749 79933
rect 145051 79932 145056 79962
rect 145112 79932 145117 79962
rect 145652 79962 145761 79964
rect 145419 79932 145485 79933
rect 145652 79932 145700 79962
rect 144284 79906 144316 79932
rect 144223 79901 144316 79906
rect 144272 79870 144316 79901
rect 144310 79868 144316 79870
rect 144380 79868 144386 79932
rect 144678 79930 144684 79932
rect 144592 79870 144684 79930
rect 144678 79868 144684 79870
rect 144748 79868 144754 79932
rect 145046 79868 145052 79932
rect 145116 79930 145122 79932
rect 145414 79930 145420 79932
rect 145116 79870 145174 79930
rect 145328 79870 145420 79930
rect 145116 79868 145122 79870
rect 145414 79868 145420 79870
rect 145484 79868 145490 79932
rect 145598 79868 145604 79932
rect 145668 79906 145700 79932
rect 145756 79906 145761 79962
rect 147259 79962 147325 79967
rect 145668 79901 145761 79906
rect 145668 79870 145712 79901
rect 145668 79868 145674 79870
rect 146518 79868 146524 79932
rect 146588 79930 146594 79932
rect 147259 79930 147264 79962
rect 146588 79906 147264 79930
rect 147320 79906 147325 79962
rect 146588 79901 147325 79906
rect 147443 79962 147509 79967
rect 147719 79964 147785 79967
rect 147443 79906 147448 79962
rect 147504 79906 147509 79962
rect 147676 79962 147785 79964
rect 147676 79932 147724 79962
rect 147443 79901 147509 79906
rect 146588 79870 147322 79901
rect 146588 79868 146594 79870
rect 147622 79868 147628 79932
rect 147692 79906 147724 79932
rect 147780 79906 147785 79962
rect 147692 79901 147785 79906
rect 147903 79964 147969 79967
rect 149007 79964 149073 79967
rect 147903 79962 148012 79964
rect 147903 79906 147908 79962
rect 147964 79932 148012 79962
rect 148964 79962 149073 79964
rect 147964 79906 147996 79932
rect 147903 79901 147996 79906
rect 147692 79870 147736 79901
rect 147952 79870 147996 79901
rect 147692 79868 147698 79870
rect 147990 79868 147996 79870
rect 148060 79868 148066 79932
rect 148358 79868 148364 79932
rect 148428 79930 148434 79932
rect 148964 79930 149012 79962
rect 148428 79906 149012 79930
rect 149068 79906 149073 79962
rect 148428 79901 149073 79906
rect 149375 79964 149441 79967
rect 151307 79964 151373 79967
rect 149375 79962 149484 79964
rect 149375 79906 149380 79962
rect 149436 79932 149484 79962
rect 151307 79962 151430 79964
rect 149436 79906 149468 79932
rect 149375 79901 149468 79906
rect 148428 79870 149024 79901
rect 149424 79870 149468 79901
rect 148428 79868 148434 79870
rect 149462 79868 149468 79870
rect 149532 79868 149538 79932
rect 149646 79868 149652 79932
rect 149716 79930 149722 79932
rect 150203 79930 150269 79933
rect 149716 79928 150269 79930
rect 149716 79872 150208 79928
rect 150264 79872 150269 79928
rect 149716 79870 150269 79872
rect 149716 79868 149722 79870
rect 144683 79867 144749 79868
rect 145419 79867 145485 79868
rect 150203 79867 150269 79870
rect 150847 79930 150913 79933
rect 151307 79932 151312 79962
rect 151368 79932 151430 79962
rect 151118 79930 151124 79932
rect 150847 79928 151124 79930
rect 150847 79872 150852 79928
rect 150908 79872 151124 79928
rect 150847 79870 151124 79872
rect 150847 79867 150913 79870
rect 151118 79868 151124 79870
rect 151188 79868 151194 79932
rect 151302 79868 151308 79932
rect 151372 79904 151430 79932
rect 151632 79930 151692 80004
rect 157566 79967 157626 80142
rect 158110 80140 158116 80142
rect 158180 80140 158186 80204
rect 165102 80202 165108 80204
rect 164512 80142 165108 80202
rect 158846 80004 158852 80068
rect 158916 80066 158922 80068
rect 158916 80006 159788 80066
rect 158916 80004 158922 80006
rect 152779 79962 152845 79967
rect 153607 79964 153673 79967
rect 151767 79930 151833 79933
rect 152319 79930 152385 79933
rect 151632 79928 151833 79930
rect 151372 79868 151378 79904
rect 151632 79872 151772 79928
rect 151828 79872 151833 79928
rect 151632 79870 151833 79872
rect 151767 79867 151833 79870
rect 152276 79928 152385 79930
rect 152276 79872 152324 79928
rect 152380 79872 152385 79928
rect 152276 79867 152385 79872
rect 152595 79928 152661 79933
rect 152595 79872 152600 79928
rect 152656 79872 152661 79928
rect 152779 79906 152784 79962
rect 152840 79906 152845 79962
rect 153564 79962 153673 79964
rect 153055 79930 153121 79933
rect 152779 79901 152845 79906
rect 152920 79928 153121 79930
rect 152595 79867 152661 79872
rect 136909 79794 136975 79797
rect 136406 79792 136975 79794
rect 136406 79736 136914 79792
rect 136970 79736 136975 79792
rect 136406 79734 136975 79736
rect 136909 79731 136975 79734
rect 137142 79661 137202 79867
rect 137510 79797 137570 79867
rect 152276 79797 152336 79867
rect 152598 79797 152658 79867
rect 137461 79792 137570 79797
rect 151491 79796 151557 79797
rect 137461 79736 137466 79792
rect 137522 79736 137570 79792
rect 137461 79734 137570 79736
rect 137970 79734 149346 79794
rect 137461 79731 137527 79734
rect 136909 79658 136975 79661
rect 132450 79656 136975 79658
rect 132450 79600 136914 79656
rect 136970 79600 136975 79656
rect 132450 79598 136975 79600
rect 137142 79656 137251 79661
rect 137142 79600 137190 79656
rect 137246 79600 137251 79656
rect 137142 79598 137251 79600
rect 136909 79595 136975 79598
rect 137185 79595 137251 79598
rect 116301 79522 116367 79525
rect 137970 79522 138030 79734
rect 139117 79656 139183 79661
rect 139117 79600 139122 79656
rect 139178 79600 139183 79656
rect 139117 79595 139183 79600
rect 140037 79658 140103 79661
rect 142797 79658 142863 79661
rect 140037 79656 142863 79658
rect 140037 79600 140042 79656
rect 140098 79600 142802 79656
rect 142858 79600 142863 79656
rect 140037 79598 142863 79600
rect 140037 79595 140103 79598
rect 142797 79595 142863 79598
rect 143022 79596 143028 79660
rect 143092 79658 143098 79660
rect 143165 79658 143231 79661
rect 143092 79656 143231 79658
rect 143092 79600 143170 79656
rect 143226 79600 143231 79656
rect 143092 79598 143231 79600
rect 143092 79596 143098 79598
rect 143165 79595 143231 79598
rect 146334 79596 146340 79660
rect 146404 79658 146410 79660
rect 146661 79658 146727 79661
rect 146404 79656 146727 79658
rect 146404 79600 146666 79656
rect 146722 79600 146727 79656
rect 146404 79598 146727 79600
rect 146404 79596 146410 79598
rect 146661 79595 146727 79598
rect 147254 79596 147260 79660
rect 147324 79658 147330 79660
rect 147673 79658 147739 79661
rect 147324 79656 147739 79658
rect 147324 79600 147678 79656
rect 147734 79600 147739 79656
rect 147324 79598 147739 79600
rect 147324 79596 147330 79598
rect 147673 79595 147739 79598
rect 147806 79596 147812 79660
rect 147876 79658 147882 79660
rect 148041 79658 148107 79661
rect 148961 79660 149027 79661
rect 147876 79656 148107 79658
rect 147876 79600 148046 79656
rect 148102 79600 148107 79656
rect 147876 79598 148107 79600
rect 147876 79596 147882 79598
rect 148041 79595 148107 79598
rect 148910 79596 148916 79660
rect 148980 79658 149027 79660
rect 148980 79656 149072 79658
rect 149022 79600 149072 79656
rect 148980 79598 149072 79600
rect 148980 79596 149027 79598
rect 148961 79595 149027 79596
rect 116301 79520 138030 79522
rect 116301 79464 116306 79520
rect 116362 79464 138030 79520
rect 116301 79462 138030 79464
rect 138841 79522 138907 79525
rect 139120 79522 139180 79595
rect 138841 79520 139180 79522
rect 138841 79464 138846 79520
rect 138902 79464 139180 79520
rect 138841 79462 139180 79464
rect 140681 79522 140747 79525
rect 140814 79522 140820 79524
rect 140681 79520 140820 79522
rect 140681 79464 140686 79520
rect 140742 79464 140820 79520
rect 140681 79462 140820 79464
rect 116301 79459 116367 79462
rect 138841 79459 138907 79462
rect 140681 79459 140747 79462
rect 140814 79460 140820 79462
rect 140884 79460 140890 79524
rect 142521 79522 142587 79525
rect 142654 79522 142660 79524
rect 142521 79520 142660 79522
rect 142521 79464 142526 79520
rect 142582 79464 142660 79520
rect 142521 79462 142660 79464
rect 142521 79459 142587 79462
rect 142654 79460 142660 79462
rect 142724 79460 142730 79524
rect 143165 79522 143231 79525
rect 143390 79522 143396 79524
rect 143165 79520 143396 79522
rect 143165 79464 143170 79520
rect 143226 79464 143396 79520
rect 143165 79462 143396 79464
rect 143165 79459 143231 79462
rect 143390 79460 143396 79462
rect 143460 79460 143466 79524
rect 143717 79522 143783 79525
rect 145005 79524 145071 79525
rect 144678 79522 144684 79524
rect 143717 79520 144684 79522
rect 143717 79464 143722 79520
rect 143778 79464 144684 79520
rect 143717 79462 144684 79464
rect 143717 79459 143783 79462
rect 144678 79460 144684 79462
rect 144748 79460 144754 79524
rect 145005 79522 145052 79524
rect 144960 79520 145052 79522
rect 144960 79464 145010 79520
rect 144960 79462 145052 79464
rect 145005 79460 145052 79462
rect 145116 79460 145122 79524
rect 147806 79460 147812 79524
rect 147876 79522 147882 79524
rect 148869 79522 148935 79525
rect 147876 79520 148935 79522
rect 147876 79464 148874 79520
rect 148930 79464 148935 79520
rect 147876 79462 148935 79464
rect 149286 79522 149346 79734
rect 151486 79732 151492 79796
rect 151556 79794 151562 79796
rect 151556 79734 151648 79794
rect 152273 79792 152339 79797
rect 152273 79736 152278 79792
rect 152334 79736 152339 79792
rect 151556 79732 151562 79734
rect 151491 79731 151557 79732
rect 152273 79731 152339 79736
rect 152549 79792 152658 79797
rect 152549 79736 152554 79792
rect 152610 79736 152658 79792
rect 152549 79734 152658 79736
rect 152549 79731 152615 79734
rect 152782 79661 152842 79901
rect 152733 79656 152842 79661
rect 152733 79600 152738 79656
rect 152794 79600 152842 79656
rect 152733 79598 152842 79600
rect 152920 79872 153060 79928
rect 153116 79872 153121 79928
rect 152920 79870 153121 79872
rect 152733 79595 152799 79598
rect 151445 79522 151511 79525
rect 149286 79520 151511 79522
rect 149286 79464 151450 79520
rect 151506 79464 151511 79520
rect 149286 79462 151511 79464
rect 147876 79460 147882 79462
rect 145005 79459 145071 79460
rect 148869 79459 148935 79462
rect 151445 79459 151511 79462
rect 152406 79460 152412 79524
rect 152476 79522 152482 79524
rect 152920 79522 152980 79870
rect 153055 79867 153121 79870
rect 153564 79906 153612 79962
rect 153668 79906 153673 79962
rect 154251 79962 154317 79967
rect 153883 79932 153949 79933
rect 154251 79932 154256 79962
rect 154312 79932 154317 79962
rect 155263 79964 155329 79967
rect 155263 79962 155372 79964
rect 153878 79930 153884 79932
rect 153564 79901 153673 79906
rect 153285 79794 153351 79797
rect 153564 79794 153624 79901
rect 153792 79870 153884 79930
rect 153878 79868 153884 79870
rect 153948 79868 153954 79932
rect 154246 79868 154252 79932
rect 154316 79930 154322 79932
rect 154711 79930 154777 79933
rect 154316 79870 154374 79930
rect 154711 79928 154820 79930
rect 154711 79872 154716 79928
rect 154772 79872 154820 79928
rect 155263 79906 155268 79962
rect 155324 79930 155372 79962
rect 157563 79962 157629 79967
rect 158391 79964 158457 79967
rect 155718 79930 155724 79932
rect 155324 79906 155724 79930
rect 155263 79901 155724 79906
rect 154316 79868 154322 79870
rect 153883 79867 153949 79868
rect 154711 79867 154820 79872
rect 155312 79870 155724 79901
rect 155718 79868 155724 79870
rect 155788 79868 155794 79932
rect 156459 79928 156525 79933
rect 156459 79872 156464 79928
rect 156520 79872 156525 79928
rect 156459 79867 156525 79872
rect 156822 79868 156828 79932
rect 156892 79930 156898 79932
rect 157011 79930 157077 79933
rect 157195 79932 157261 79933
rect 156892 79928 157077 79930
rect 156892 79872 157016 79928
rect 157072 79872 157077 79928
rect 156892 79870 157077 79872
rect 156892 79868 156898 79870
rect 157011 79867 157077 79870
rect 157190 79868 157196 79932
rect 157260 79930 157266 79932
rect 157260 79870 157352 79930
rect 157563 79906 157568 79962
rect 157624 79906 157629 79962
rect 158348 79962 158457 79964
rect 157563 79901 157629 79906
rect 157747 79928 157813 79933
rect 158348 79932 158396 79962
rect 157747 79872 157752 79928
rect 157808 79872 157813 79928
rect 157260 79868 157266 79870
rect 157195 79867 157261 79868
rect 157747 79867 157813 79872
rect 158294 79868 158300 79932
rect 158364 79906 158396 79932
rect 158452 79906 158457 79962
rect 159587 79930 159653 79933
rect 158364 79901 158457 79906
rect 159222 79928 159653 79930
rect 158364 79870 158408 79901
rect 159222 79872 159592 79928
rect 159648 79872 159653 79928
rect 159222 79870 159653 79872
rect 159728 79930 159788 80006
rect 164512 79967 164572 80142
rect 165102 80140 165108 80142
rect 165172 80140 165178 80204
rect 174080 80202 174140 80278
rect 181621 80275 181687 80278
rect 187734 80276 187740 80340
rect 187804 80338 187810 80340
rect 188889 80338 188955 80341
rect 187804 80336 188955 80338
rect 187804 80280 188894 80336
rect 188950 80280 188955 80336
rect 187804 80278 188955 80280
rect 187804 80276 187810 80278
rect 188889 80275 188955 80278
rect 181662 80202 181668 80204
rect 173942 80142 174140 80202
rect 174264 80142 181668 80202
rect 173758 80066 173864 80070
rect 171688 80006 173864 80066
rect 162255 79962 162321 79967
rect 160047 79930 160113 79933
rect 159728 79928 160113 79930
rect 159728 79872 160052 79928
rect 160108 79872 160113 79928
rect 159728 79870 160113 79872
rect 158364 79868 158370 79870
rect 153285 79792 153624 79794
rect 153285 79736 153290 79792
rect 153346 79736 153624 79792
rect 153285 79734 153624 79736
rect 154021 79792 154087 79797
rect 154021 79736 154026 79792
rect 154082 79736 154087 79792
rect 153285 79731 153351 79734
rect 154021 79731 154087 79736
rect 154389 79796 154455 79797
rect 154389 79792 154436 79796
rect 154500 79794 154506 79796
rect 154389 79736 154394 79792
rect 154389 79732 154436 79736
rect 154500 79734 154546 79794
rect 154500 79732 154506 79734
rect 154389 79731 154455 79732
rect 154024 79525 154084 79731
rect 154760 79661 154820 79867
rect 155309 79794 155375 79797
rect 155534 79794 155540 79796
rect 155309 79792 155540 79794
rect 155309 79736 155314 79792
rect 155370 79736 155540 79792
rect 155309 79734 155540 79736
rect 155309 79731 155375 79734
rect 155534 79732 155540 79734
rect 155604 79732 155610 79796
rect 154757 79656 154823 79661
rect 154757 79600 154762 79656
rect 154818 79600 154823 79656
rect 154757 79595 154823 79600
rect 152476 79462 152980 79522
rect 154021 79520 154087 79525
rect 154021 79464 154026 79520
rect 154082 79464 154087 79520
rect 152476 79460 152482 79462
rect 154021 79459 154087 79464
rect 156137 79522 156203 79525
rect 156462 79522 156522 79867
rect 156137 79520 156522 79522
rect 156137 79464 156142 79520
rect 156198 79464 156522 79520
rect 156137 79462 156522 79464
rect 157750 79525 157810 79867
rect 158115 79826 158181 79831
rect 158115 79770 158120 79826
rect 158176 79770 158181 79826
rect 158115 79765 158181 79770
rect 158299 79794 158365 79797
rect 158478 79794 158484 79796
rect 158299 79792 158484 79794
rect 157885 79658 157951 79661
rect 158118 79658 158178 79765
rect 158299 79736 158304 79792
rect 158360 79736 158484 79792
rect 158299 79734 158484 79736
rect 158299 79731 158365 79734
rect 158478 79732 158484 79734
rect 158548 79732 158554 79796
rect 158851 79792 158917 79797
rect 158851 79736 158856 79792
rect 158912 79736 158917 79792
rect 158851 79731 158917 79736
rect 157885 79656 158178 79658
rect 157885 79600 157890 79656
rect 157946 79600 158178 79656
rect 157885 79598 158178 79600
rect 158854 79658 158914 79731
rect 159081 79658 159147 79661
rect 158854 79656 159147 79658
rect 158854 79600 159086 79656
rect 159142 79600 159147 79656
rect 158854 79598 159147 79600
rect 157885 79595 157951 79598
rect 159081 79595 159147 79598
rect 157750 79520 157859 79525
rect 157750 79464 157798 79520
rect 157854 79464 157859 79520
rect 157750 79462 157859 79464
rect 156137 79459 156203 79462
rect 157793 79459 157859 79462
rect 158713 79522 158779 79525
rect 159222 79522 159282 79870
rect 159587 79867 159653 79870
rect 160047 79867 160113 79870
rect 160415 79928 160481 79933
rect 160875 79932 160941 79933
rect 160870 79930 160876 79932
rect 160415 79872 160420 79928
rect 160476 79872 160481 79928
rect 160415 79867 160481 79872
rect 160784 79870 160876 79930
rect 160870 79868 160876 79870
rect 160940 79868 160946 79932
rect 162255 79906 162260 79962
rect 162316 79906 162321 79962
rect 162255 79901 162321 79906
rect 162623 79962 162689 79967
rect 162623 79906 162628 79962
rect 162684 79906 162689 79962
rect 163635 79962 163701 79967
rect 164279 79964 164345 79967
rect 162623 79901 162689 79906
rect 160875 79867 160941 79868
rect 160418 79794 160478 79867
rect 160829 79794 160895 79797
rect 160418 79792 160895 79794
rect 160418 79736 160834 79792
rect 160890 79736 160895 79792
rect 160418 79734 160895 79736
rect 160829 79731 160895 79734
rect 160967 79794 161033 79797
rect 162258 79794 162318 79901
rect 160967 79792 161168 79794
rect 160967 79736 160972 79792
rect 161028 79736 161168 79792
rect 160967 79734 161168 79736
rect 160967 79731 161033 79734
rect 159449 79658 159515 79661
rect 158713 79520 159282 79522
rect 158713 79464 158718 79520
rect 158774 79464 159282 79520
rect 158713 79462 159282 79464
rect 159406 79656 159515 79658
rect 159406 79600 159454 79656
rect 159510 79600 159515 79656
rect 159406 79595 159515 79600
rect 158713 79459 158779 79462
rect 113766 79324 113772 79388
rect 113836 79386 113842 79388
rect 127801 79386 127867 79389
rect 113836 79384 127867 79386
rect 113836 79328 127806 79384
rect 127862 79328 127867 79384
rect 113836 79326 127867 79328
rect 113836 79324 113842 79326
rect 127801 79323 127867 79326
rect 136582 79324 136588 79388
rect 136652 79386 136658 79388
rect 137001 79386 137067 79389
rect 136652 79384 137067 79386
rect 136652 79328 137006 79384
rect 137062 79328 137067 79384
rect 136652 79326 137067 79328
rect 136652 79324 136658 79326
rect 137001 79323 137067 79326
rect 139117 79386 139183 79389
rect 139894 79386 139900 79388
rect 139117 79384 139900 79386
rect 139117 79328 139122 79384
rect 139178 79328 139900 79384
rect 139117 79326 139900 79328
rect 139117 79323 139183 79326
rect 139894 79324 139900 79326
rect 139964 79324 139970 79388
rect 142705 79386 142771 79389
rect 147765 79386 147831 79389
rect 147949 79386 148015 79389
rect 142705 79384 148015 79386
rect 142705 79328 142710 79384
rect 142766 79328 147770 79384
rect 147826 79328 147954 79384
rect 148010 79328 148015 79384
rect 142705 79326 148015 79328
rect 142705 79323 142771 79326
rect 147765 79323 147831 79326
rect 147949 79323 148015 79326
rect 151302 79324 151308 79388
rect 151372 79386 151378 79388
rect 151629 79386 151695 79389
rect 151372 79384 151695 79386
rect 151372 79328 151634 79384
rect 151690 79328 151695 79384
rect 151372 79326 151695 79328
rect 159406 79386 159466 79595
rect 160829 79522 160895 79525
rect 161108 79522 161168 79734
rect 162212 79734 162318 79794
rect 162212 79660 162272 79734
rect 162158 79596 162164 79660
rect 162228 79598 162272 79660
rect 162228 79596 162234 79598
rect 162342 79596 162348 79660
rect 162412 79658 162418 79660
rect 162485 79658 162551 79661
rect 162412 79656 162551 79658
rect 162412 79600 162490 79656
rect 162546 79600 162551 79656
rect 162412 79598 162551 79600
rect 162412 79596 162418 79598
rect 162485 79595 162551 79598
rect 160829 79520 161168 79522
rect 160829 79464 160834 79520
rect 160890 79464 161168 79520
rect 160829 79462 161168 79464
rect 162626 79522 162686 79901
rect 163262 79868 163268 79932
rect 163332 79930 163338 79932
rect 163635 79930 163640 79962
rect 163332 79906 163640 79930
rect 163696 79906 163701 79962
rect 164236 79962 164345 79964
rect 164003 79932 164069 79933
rect 164236 79932 164284 79962
rect 163998 79930 164004 79932
rect 163332 79901 163701 79906
rect 163332 79870 163698 79901
rect 163912 79870 164004 79930
rect 163332 79868 163338 79870
rect 163998 79868 164004 79870
rect 164068 79868 164074 79932
rect 164182 79868 164188 79932
rect 164252 79906 164284 79932
rect 164340 79906 164345 79962
rect 164252 79901 164345 79906
rect 164463 79962 164572 79967
rect 164463 79906 164468 79962
rect 164524 79906 164572 79962
rect 166119 79962 166185 79967
rect 164463 79904 164572 79906
rect 164923 79930 164989 79933
rect 165659 79932 165725 79933
rect 165843 79932 165909 79933
rect 165286 79930 165292 79932
rect 164923 79928 165292 79930
rect 164463 79901 164529 79904
rect 164252 79870 164296 79901
rect 164923 79872 164928 79928
rect 164984 79872 165292 79928
rect 164923 79870 165292 79872
rect 164252 79868 164258 79870
rect 164003 79867 164069 79868
rect 164923 79867 164989 79870
rect 165286 79868 165292 79870
rect 165356 79868 165362 79932
rect 165654 79930 165660 79932
rect 165568 79870 165660 79930
rect 165654 79868 165660 79870
rect 165724 79868 165730 79932
rect 165838 79868 165844 79932
rect 165908 79930 165914 79932
rect 165908 79870 166000 79930
rect 166119 79906 166124 79962
rect 166180 79930 166185 79962
rect 167683 79962 167749 79967
rect 166390 79930 166396 79932
rect 166180 79906 166396 79930
rect 166119 79901 166396 79906
rect 166122 79870 166396 79901
rect 165908 79868 165914 79870
rect 166390 79868 166396 79870
rect 166460 79868 166466 79932
rect 167683 79906 167688 79962
rect 167744 79930 167749 79962
rect 168787 79962 168853 79967
rect 167862 79930 167868 79932
rect 167744 79906 167868 79930
rect 167683 79901 167868 79906
rect 167223 79896 167289 79899
rect 167223 79894 167332 79896
rect 165659 79867 165725 79868
rect 165843 79867 165909 79868
rect 167223 79838 167228 79894
rect 167284 79838 167332 79894
rect 167686 79870 167868 79901
rect 167862 79868 167868 79870
rect 167932 79868 167938 79932
rect 168051 79930 168117 79933
rect 168603 79930 168669 79933
rect 168051 79928 168298 79930
rect 168051 79872 168056 79928
rect 168112 79872 168298 79928
rect 168051 79870 168298 79872
rect 168051 79867 168117 79870
rect 167223 79833 167332 79838
rect 166579 79792 166645 79797
rect 166579 79736 166584 79792
rect 166640 79736 166645 79792
rect 166579 79731 166645 79736
rect 166758 79732 166764 79796
rect 166828 79794 166834 79796
rect 166947 79794 167013 79797
rect 166828 79792 167013 79794
rect 166828 79736 166952 79792
rect 167008 79736 167013 79792
rect 166828 79734 167013 79736
rect 166828 79732 166834 79734
rect 166947 79731 167013 79734
rect 166582 79661 166642 79731
rect 167272 79661 167332 79833
rect 167867 79794 167933 79797
rect 168046 79794 168052 79796
rect 167867 79792 168052 79794
rect 167867 79736 167872 79792
rect 167928 79736 168052 79792
rect 167867 79734 168052 79736
rect 167867 79731 167933 79734
rect 168046 79732 168052 79734
rect 168116 79732 168122 79796
rect 162853 79658 162919 79661
rect 163497 79658 163563 79661
rect 162853 79656 163563 79658
rect 162853 79600 162858 79656
rect 162914 79600 163502 79656
rect 163558 79600 163563 79656
rect 162853 79598 163563 79600
rect 162853 79595 162919 79598
rect 163497 79595 163563 79598
rect 166533 79656 166642 79661
rect 166533 79600 166538 79656
rect 166594 79600 166642 79656
rect 166533 79598 166642 79600
rect 167269 79656 167335 79661
rect 167269 79600 167274 79656
rect 167330 79600 167335 79656
rect 166533 79595 166599 79598
rect 167269 79595 167335 79600
rect 163681 79522 163747 79525
rect 162626 79520 163747 79522
rect 162626 79464 163686 79520
rect 163742 79464 163747 79520
rect 162626 79462 163747 79464
rect 160829 79459 160895 79462
rect 163681 79459 163747 79462
rect 163446 79386 163452 79388
rect 159406 79326 163452 79386
rect 151372 79324 151378 79326
rect 151629 79323 151695 79326
rect 163446 79324 163452 79326
rect 163516 79324 163522 79388
rect 167269 79386 167335 79389
rect 168238 79386 168298 79870
rect 168376 79928 168669 79930
rect 168376 79872 168608 79928
rect 168664 79872 168669 79928
rect 168787 79906 168792 79962
rect 168848 79906 168853 79962
rect 170443 79962 170509 79967
rect 168787 79901 168853 79906
rect 168376 79870 168669 79872
rect 168376 79797 168436 79870
rect 168603 79867 168669 79870
rect 168373 79792 168439 79797
rect 168373 79736 168378 79792
rect 168434 79736 168439 79792
rect 168373 79731 168439 79736
rect 168557 79794 168623 79797
rect 168790 79794 168850 79901
rect 168966 79868 168972 79932
rect 169036 79930 169042 79932
rect 169431 79930 169497 79933
rect 169615 79930 169681 79933
rect 169036 79928 169497 79930
rect 169036 79872 169436 79928
rect 169492 79872 169497 79928
rect 169036 79870 169497 79872
rect 169036 79868 169042 79870
rect 169431 79867 169497 79870
rect 169572 79928 169681 79930
rect 169572 79872 169620 79928
rect 169676 79872 169681 79928
rect 169572 79867 169681 79872
rect 169799 79930 169865 79933
rect 170254 79930 170260 79932
rect 169799 79928 170260 79930
rect 169799 79872 169804 79928
rect 169860 79872 170260 79928
rect 169799 79870 170260 79872
rect 169799 79867 169865 79870
rect 170254 79868 170260 79870
rect 170324 79868 170330 79932
rect 170443 79906 170448 79962
rect 170504 79906 170509 79962
rect 170627 79962 170693 79967
rect 170627 79932 170632 79962
rect 170688 79932 170693 79962
rect 170443 79901 170509 79906
rect 168557 79792 168850 79794
rect 168557 79736 168562 79792
rect 168618 79736 168850 79792
rect 168557 79734 168850 79736
rect 169017 79794 169083 79797
rect 169385 79794 169451 79797
rect 169017 79792 169451 79794
rect 169017 79736 169022 79792
rect 169078 79736 169390 79792
rect 169446 79736 169451 79792
rect 169017 79734 169451 79736
rect 169572 79794 169632 79867
rect 169753 79794 169819 79797
rect 170075 79796 170141 79797
rect 170070 79794 170076 79796
rect 169572 79792 169819 79794
rect 169572 79736 169758 79792
rect 169814 79736 169819 79792
rect 169572 79734 169819 79736
rect 169984 79734 170076 79794
rect 168557 79731 168623 79734
rect 169017 79731 169083 79734
rect 169385 79731 169451 79734
rect 169753 79731 169819 79734
rect 170070 79732 170076 79734
rect 170140 79732 170146 79796
rect 170075 79731 170141 79732
rect 170213 79658 170279 79661
rect 170446 79658 170506 79901
rect 170622 79868 170628 79932
rect 170692 79930 170698 79932
rect 170692 79870 170750 79930
rect 170995 79928 171061 79933
rect 170995 79872 171000 79928
rect 171056 79872 171061 79928
rect 170692 79868 170698 79870
rect 170995 79867 171061 79872
rect 171455 79930 171521 79933
rect 171688 79930 171748 80006
rect 172835 79930 172901 79933
rect 171455 79928 171748 79930
rect 171455 79872 171460 79928
rect 171516 79872 171748 79928
rect 171455 79870 171748 79872
rect 171455 79867 171521 79870
rect 170998 79797 171058 79867
rect 170949 79792 171058 79797
rect 170949 79736 170954 79792
rect 171010 79736 171058 79792
rect 170949 79734 171058 79736
rect 171225 79794 171291 79797
rect 171542 79794 171548 79796
rect 171225 79792 171548 79794
rect 171225 79736 171230 79792
rect 171286 79736 171548 79792
rect 171225 79734 171548 79736
rect 170949 79731 171015 79734
rect 171225 79731 171291 79734
rect 171542 79732 171548 79734
rect 171612 79732 171618 79796
rect 170213 79656 170506 79658
rect 170213 79600 170218 79656
rect 170274 79600 170506 79656
rect 170213 79598 170506 79600
rect 171317 79658 171383 79661
rect 171688 79658 171748 79870
rect 172700 79928 172901 79930
rect 172700 79872 172840 79928
rect 172896 79872 172901 79928
rect 172700 79870 172901 79872
rect 172700 79797 172760 79870
rect 172835 79867 172901 79870
rect 173382 79868 173388 79932
rect 173452 79930 173458 79932
rect 173663 79930 173729 79933
rect 173452 79928 173729 79930
rect 173452 79872 173668 79928
rect 173724 79872 173729 79928
rect 173452 79870 173729 79872
rect 173804 79930 173864 80006
rect 173942 79930 174002 80142
rect 173804 79870 174002 79930
rect 174123 79962 174189 79967
rect 174123 79906 174128 79962
rect 174184 79906 174189 79962
rect 174123 79901 174189 79906
rect 173452 79868 173458 79870
rect 173663 79867 173729 79870
rect 174126 79831 174186 79901
rect 174123 79826 174189 79831
rect 172145 79794 172211 79797
rect 172278 79794 172284 79796
rect 172145 79792 172284 79794
rect 172145 79736 172150 79792
rect 172206 79736 172284 79792
rect 172145 79734 172284 79736
rect 172145 79731 172211 79734
rect 172278 79732 172284 79734
rect 172348 79732 172354 79796
rect 172697 79792 172763 79797
rect 172697 79736 172702 79792
rect 172758 79736 172763 79792
rect 172697 79731 172763 79736
rect 172830 79732 172836 79796
rect 172900 79794 172906 79796
rect 173111 79794 173177 79797
rect 172900 79792 173177 79794
rect 172900 79736 173116 79792
rect 173172 79736 173177 79792
rect 172900 79734 173177 79736
rect 172900 79732 172906 79734
rect 173111 79731 173177 79734
rect 173387 79792 173453 79797
rect 173387 79736 173392 79792
rect 173448 79736 173453 79792
rect 173387 79731 173453 79736
rect 173566 79732 173572 79796
rect 173636 79794 173642 79796
rect 173847 79794 173913 79797
rect 173636 79792 173913 79794
rect 173636 79736 173852 79792
rect 173908 79736 173913 79792
rect 174123 79770 174128 79826
rect 174184 79770 174189 79826
rect 174123 79765 174189 79770
rect 173636 79734 173913 79736
rect 173636 79732 173642 79734
rect 173847 79731 173913 79734
rect 171317 79656 171748 79658
rect 171317 79600 171322 79656
rect 171378 79600 171748 79656
rect 171317 79598 171748 79600
rect 172789 79658 172855 79661
rect 173390 79658 173450 79731
rect 174264 79658 174324 80142
rect 181662 80140 181668 80142
rect 181732 80140 181738 80204
rect 175222 80066 175228 80068
rect 174908 80006 175228 80066
rect 174399 79930 174465 79933
rect 174767 79930 174833 79933
rect 174908 79930 174968 80006
rect 175222 80004 175228 80006
rect 175292 80004 175298 80068
rect 200798 80004 200804 80068
rect 200868 80066 200874 80068
rect 201309 80066 201375 80069
rect 200868 80064 201375 80066
rect 200868 80008 201314 80064
rect 201370 80008 201375 80064
rect 200868 80006 201375 80008
rect 200868 80004 200874 80006
rect 201309 80003 201375 80006
rect 175595 79962 175661 79967
rect 174399 79928 174508 79930
rect 174399 79872 174404 79928
rect 174460 79872 174508 79928
rect 174399 79867 174508 79872
rect 174767 79928 174968 79930
rect 174767 79872 174772 79928
rect 174828 79872 174968 79928
rect 174767 79870 174968 79872
rect 175043 79930 175109 79933
rect 175406 79930 175412 79932
rect 175043 79928 175412 79930
rect 175043 79872 175048 79928
rect 175104 79872 175412 79928
rect 175043 79870 175412 79872
rect 174767 79867 174833 79870
rect 175043 79867 175109 79870
rect 175406 79868 175412 79870
rect 175476 79868 175482 79932
rect 175595 79906 175600 79962
rect 175656 79906 175661 79962
rect 176055 79962 176121 79967
rect 176055 79930 176060 79962
rect 175595 79901 175661 79906
rect 176012 79906 176060 79930
rect 176116 79906 176121 79962
rect 176012 79901 176121 79906
rect 176239 79930 176305 79933
rect 176510 79930 176516 79932
rect 176239 79928 176516 79930
rect 172789 79656 174324 79658
rect 172789 79600 172794 79656
rect 172850 79600 174324 79656
rect 172789 79598 174324 79600
rect 174448 79658 174508 79867
rect 174670 79732 174676 79796
rect 174740 79794 174746 79796
rect 175227 79794 175293 79797
rect 174740 79792 175293 79794
rect 174740 79736 175232 79792
rect 175288 79736 175293 79792
rect 174740 79734 175293 79736
rect 174740 79732 174746 79734
rect 175227 79731 175293 79734
rect 175598 79661 175658 79901
rect 175779 79894 175845 79899
rect 175779 79838 175784 79894
rect 175840 79838 175845 79894
rect 175779 79833 175845 79838
rect 176012 79870 176118 79901
rect 176239 79872 176244 79928
rect 176300 79872 176516 79928
rect 176239 79870 176516 79872
rect 175782 79661 175842 79833
rect 176012 79796 176072 79870
rect 176239 79867 176305 79870
rect 176510 79868 176516 79870
rect 176580 79868 176586 79932
rect 177435 79930 177501 79933
rect 180517 79930 180583 79933
rect 177435 79928 180583 79930
rect 177435 79872 177440 79928
rect 177496 79872 180522 79928
rect 180578 79872 180583 79928
rect 177435 79870 180583 79872
rect 177435 79867 177501 79870
rect 180517 79867 180583 79870
rect 175958 79732 175964 79796
rect 176028 79734 176072 79796
rect 176028 79732 176034 79734
rect 174629 79658 174695 79661
rect 174448 79656 174695 79658
rect 174448 79600 174634 79656
rect 174690 79600 174695 79656
rect 174448 79598 174695 79600
rect 170213 79595 170279 79598
rect 171317 79595 171383 79598
rect 172789 79595 172855 79598
rect 174629 79595 174695 79598
rect 175549 79656 175658 79661
rect 175549 79600 175554 79656
rect 175610 79600 175658 79656
rect 175549 79598 175658 79600
rect 175733 79656 175842 79661
rect 175733 79600 175738 79656
rect 175794 79600 175842 79656
rect 175733 79598 175842 79600
rect 175549 79595 175615 79598
rect 175733 79595 175799 79598
rect 168925 79522 168991 79525
rect 190494 79522 190500 79524
rect 168925 79520 190500 79522
rect 168925 79464 168930 79520
rect 168986 79464 190500 79520
rect 168925 79462 190500 79464
rect 168925 79459 168991 79462
rect 190494 79460 190500 79462
rect 190564 79460 190570 79524
rect 192150 79386 192156 79388
rect 167269 79384 192156 79386
rect 167269 79328 167274 79384
rect 167330 79328 192156 79384
rect 167269 79326 192156 79328
rect 167269 79323 167335 79326
rect 192150 79324 192156 79326
rect 192220 79324 192226 79388
rect 108113 79250 108179 79253
rect 108665 79250 108731 79253
rect 141233 79250 141299 79253
rect 108113 79248 141299 79250
rect 108113 79192 108118 79248
rect 108174 79192 108670 79248
rect 108726 79192 141238 79248
rect 141294 79192 141299 79248
rect 108113 79190 141299 79192
rect 108113 79187 108179 79190
rect 108665 79187 108731 79190
rect 141233 79187 141299 79190
rect 141417 79250 141483 79253
rect 142245 79250 142311 79253
rect 141417 79248 142311 79250
rect 141417 79192 141422 79248
rect 141478 79192 142250 79248
rect 142306 79192 142311 79248
rect 141417 79190 142311 79192
rect 141417 79187 141483 79190
rect 142245 79187 142311 79190
rect 146753 79250 146819 79253
rect 146886 79250 146892 79252
rect 146753 79248 146892 79250
rect 146753 79192 146758 79248
rect 146814 79192 146892 79248
rect 146753 79190 146892 79192
rect 146753 79187 146819 79190
rect 146886 79188 146892 79190
rect 146956 79188 146962 79252
rect 147622 79188 147628 79252
rect 147692 79250 147698 79252
rect 147857 79250 147923 79253
rect 147692 79248 147923 79250
rect 147692 79192 147862 79248
rect 147918 79192 147923 79248
rect 147692 79190 147923 79192
rect 147692 79188 147698 79190
rect 147857 79187 147923 79190
rect 157977 79250 158043 79253
rect 162577 79250 162643 79253
rect 157977 79248 162643 79250
rect 157977 79192 157982 79248
rect 158038 79192 162582 79248
rect 162638 79192 162643 79248
rect 157977 79190 162643 79192
rect 157977 79187 158043 79190
rect 162577 79187 162643 79190
rect 162945 79250 163011 79253
rect 163998 79250 164004 79252
rect 162945 79248 164004 79250
rect 162945 79192 162950 79248
rect 163006 79192 164004 79248
rect 162945 79190 164004 79192
rect 162945 79187 163011 79190
rect 163998 79188 164004 79190
rect 164068 79188 164074 79252
rect 165521 79250 165587 79253
rect 189390 79250 189396 79252
rect 165521 79248 189396 79250
rect 165521 79192 165526 79248
rect 165582 79192 189396 79248
rect 165521 79190 189396 79192
rect 165521 79187 165587 79190
rect 189390 79188 189396 79190
rect 189460 79188 189466 79252
rect 117865 79114 117931 79117
rect 150525 79114 150591 79117
rect 151721 79114 151787 79117
rect 117865 79112 151787 79114
rect 117865 79056 117870 79112
rect 117926 79056 150530 79112
rect 150586 79056 151726 79112
rect 151782 79056 151787 79112
rect 117865 79054 151787 79056
rect 117865 79051 117931 79054
rect 150525 79051 150591 79054
rect 151721 79051 151787 79054
rect 164141 79114 164207 79117
rect 190678 79114 190684 79116
rect 164141 79112 190684 79114
rect 164141 79056 164146 79112
rect 164202 79056 190684 79112
rect 164141 79054 190684 79056
rect 164141 79051 164207 79054
rect 190678 79052 190684 79054
rect 190748 79052 190754 79116
rect 116209 78978 116275 78981
rect 155953 78978 156019 78981
rect 157006 78978 157012 78980
rect 116209 78976 149530 78978
rect 116209 78920 116214 78976
rect 116270 78920 149530 78976
rect 116209 78918 149530 78920
rect 116209 78915 116275 78918
rect 127801 78842 127867 78845
rect 128169 78842 128235 78845
rect 145189 78842 145255 78845
rect 149470 78844 149530 78918
rect 155953 78976 157012 78978
rect 155953 78920 155958 78976
rect 156014 78920 157012 78976
rect 155953 78918 157012 78920
rect 155953 78915 156019 78918
rect 157006 78916 157012 78918
rect 157076 78916 157082 78980
rect 164918 78916 164924 78980
rect 164988 78978 164994 78980
rect 165429 78978 165495 78981
rect 164988 78976 165495 78978
rect 164988 78920 165434 78976
rect 165490 78920 165495 78976
rect 164988 78918 165495 78920
rect 164988 78916 164994 78918
rect 165429 78915 165495 78918
rect 168741 78978 168807 78981
rect 169334 78978 169340 78980
rect 168741 78976 169340 78978
rect 168741 78920 168746 78976
rect 168802 78920 169340 78976
rect 168741 78918 169340 78920
rect 168741 78915 168807 78918
rect 169334 78916 169340 78918
rect 169404 78916 169410 78980
rect 172881 78978 172947 78981
rect 174261 78980 174327 78981
rect 173014 78978 173020 78980
rect 172881 78976 173020 78978
rect 172881 78920 172886 78976
rect 172942 78920 173020 78976
rect 172881 78918 173020 78920
rect 172881 78915 172947 78918
rect 173014 78916 173020 78918
rect 173084 78916 173090 78980
rect 174261 78978 174308 78980
rect 174216 78976 174308 78978
rect 174216 78920 174266 78976
rect 174216 78918 174308 78920
rect 174261 78916 174308 78918
rect 174372 78916 174378 78980
rect 178217 78978 178283 78981
rect 206134 78978 206140 78980
rect 178217 78976 206140 78978
rect 178217 78920 178222 78976
rect 178278 78920 206140 78976
rect 178217 78918 206140 78920
rect 174261 78915 174327 78916
rect 178217 78915 178283 78918
rect 206134 78916 206140 78918
rect 206204 78916 206210 78980
rect 127801 78840 145255 78842
rect 127801 78784 127806 78840
rect 127862 78784 128174 78840
rect 128230 78784 145194 78840
rect 145250 78784 145255 78840
rect 127801 78782 145255 78784
rect 127801 78779 127867 78782
rect 128169 78779 128235 78782
rect 145189 78779 145255 78782
rect 149462 78780 149468 78844
rect 149532 78842 149538 78844
rect 218697 78842 218763 78845
rect 149532 78840 218763 78842
rect 149532 78784 218702 78840
rect 218758 78784 218763 78840
rect 149532 78782 218763 78784
rect 149532 78780 149538 78782
rect 218697 78779 218763 78782
rect 137369 78706 137435 78709
rect 137870 78706 137876 78708
rect 137369 78704 137876 78706
rect 137369 78648 137374 78704
rect 137430 78648 137876 78704
rect 137369 78646 137876 78648
rect 137369 78643 137435 78646
rect 137870 78644 137876 78646
rect 137940 78644 137946 78708
rect 140630 78644 140636 78708
rect 140700 78706 140706 78708
rect 140773 78706 140839 78709
rect 140700 78704 140839 78706
rect 140700 78648 140778 78704
rect 140834 78648 140839 78704
rect 140700 78646 140839 78648
rect 140700 78644 140706 78646
rect 140773 78643 140839 78646
rect 145414 78644 145420 78708
rect 145484 78706 145490 78708
rect 145741 78706 145807 78709
rect 145484 78704 145807 78706
rect 145484 78648 145746 78704
rect 145802 78648 145807 78704
rect 145484 78646 145807 78648
rect 145484 78644 145490 78646
rect 145741 78643 145807 78646
rect 149462 78644 149468 78708
rect 149532 78706 149538 78708
rect 150433 78706 150499 78709
rect 149532 78704 150499 78706
rect 149532 78648 150438 78704
rect 150494 78648 150499 78704
rect 149532 78646 150499 78648
rect 149532 78644 149538 78646
rect 150433 78643 150499 78646
rect 151721 78706 151787 78709
rect 234613 78706 234679 78709
rect 151721 78704 234679 78706
rect 151721 78648 151726 78704
rect 151782 78648 234618 78704
rect 234674 78648 234679 78704
rect 151721 78646 234679 78648
rect 151721 78643 151787 78646
rect 234613 78643 234679 78646
rect 107510 78570 107516 78572
rect 99330 78510 107516 78570
rect 2773 77890 2839 77893
rect 99330 77890 99390 78510
rect 107510 78508 107516 78510
rect 107580 78570 107586 78572
rect 128261 78570 128327 78573
rect 107580 78568 128327 78570
rect 107580 78512 128266 78568
rect 128322 78512 128327 78568
rect 107580 78510 128327 78512
rect 107580 78508 107586 78510
rect 128261 78507 128327 78510
rect 149094 78508 149100 78572
rect 149164 78570 149170 78572
rect 150249 78570 150315 78573
rect 149164 78568 150315 78570
rect 149164 78512 150254 78568
rect 150310 78512 150315 78568
rect 149164 78510 150315 78512
rect 149164 78508 149170 78510
rect 150249 78507 150315 78510
rect 156638 78508 156644 78572
rect 156708 78570 156714 78572
rect 156965 78570 157031 78573
rect 156708 78568 157031 78570
rect 156708 78512 156970 78568
rect 157026 78512 157031 78568
rect 156708 78510 157031 78512
rect 156708 78508 156714 78510
rect 156965 78507 157031 78510
rect 157926 78508 157932 78572
rect 157996 78570 158002 78572
rect 158529 78570 158595 78573
rect 157996 78568 158595 78570
rect 157996 78512 158534 78568
rect 158590 78512 158595 78568
rect 157996 78510 158595 78512
rect 157996 78508 158002 78510
rect 158529 78507 158595 78510
rect 158805 78570 158871 78573
rect 159030 78570 159036 78572
rect 158805 78568 159036 78570
rect 158805 78512 158810 78568
rect 158866 78512 159036 78568
rect 158805 78510 159036 78512
rect 158805 78507 158871 78510
rect 159030 78508 159036 78510
rect 159100 78508 159106 78572
rect 160686 78508 160692 78572
rect 160756 78570 160762 78572
rect 161381 78570 161447 78573
rect 166625 78572 166691 78573
rect 166574 78570 166580 78572
rect 160756 78568 161447 78570
rect 160756 78512 161386 78568
rect 161442 78512 161447 78568
rect 160756 78510 161447 78512
rect 166534 78510 166580 78570
rect 166644 78568 166691 78572
rect 166686 78512 166691 78568
rect 160756 78508 160762 78510
rect 161381 78507 161447 78510
rect 166574 78508 166580 78510
rect 166644 78508 166691 78512
rect 166625 78507 166691 78508
rect 166993 78570 167059 78573
rect 167494 78570 167500 78572
rect 166993 78568 167500 78570
rect 166993 78512 166998 78568
rect 167054 78512 167500 78568
rect 166993 78510 167500 78512
rect 166993 78507 167059 78510
rect 167494 78508 167500 78510
rect 167564 78508 167570 78572
rect 168833 78568 168899 78573
rect 170581 78572 170647 78573
rect 170581 78570 170628 78572
rect 168833 78512 168838 78568
rect 168894 78512 168899 78568
rect 168833 78507 168899 78512
rect 170536 78568 170628 78570
rect 170536 78512 170586 78568
rect 170536 78510 170628 78512
rect 170581 78508 170628 78510
rect 170692 78508 170698 78572
rect 171409 78570 171475 78573
rect 181437 78570 181503 78573
rect 171409 78568 181503 78570
rect 171409 78512 171414 78568
rect 171470 78512 181442 78568
rect 181498 78512 181503 78568
rect 171409 78510 181503 78512
rect 170581 78507 170647 78508
rect 171409 78507 171475 78510
rect 181437 78507 181503 78510
rect 181621 78570 181687 78573
rect 188981 78570 189047 78573
rect 181621 78568 189047 78570
rect 181621 78512 181626 78568
rect 181682 78512 188986 78568
rect 189042 78512 189047 78568
rect 181621 78510 189047 78512
rect 181621 78507 181687 78510
rect 188981 78507 189047 78510
rect 197302 78508 197308 78572
rect 197372 78570 197378 78572
rect 197905 78570 197971 78573
rect 199009 78572 199075 78573
rect 198958 78570 198964 78572
rect 197372 78568 197971 78570
rect 197372 78512 197910 78568
rect 197966 78512 197971 78568
rect 197372 78510 197971 78512
rect 198918 78510 198964 78570
rect 199028 78568 199075 78572
rect 199070 78512 199075 78568
rect 197372 78508 197378 78510
rect 197905 78507 197971 78510
rect 198958 78508 198964 78510
rect 199028 78508 199075 78512
rect 199009 78507 199075 78508
rect 119797 78434 119863 78437
rect 120022 78434 120028 78436
rect 119797 78432 120028 78434
rect 119797 78376 119802 78432
rect 119858 78376 120028 78432
rect 119797 78374 120028 78376
rect 119797 78371 119863 78374
rect 120022 78372 120028 78374
rect 120092 78372 120098 78436
rect 122966 78372 122972 78436
rect 123036 78434 123042 78436
rect 144269 78434 144335 78437
rect 123036 78432 144335 78434
rect 123036 78376 144274 78432
rect 144330 78376 144335 78432
rect 123036 78374 144335 78376
rect 123036 78372 123042 78374
rect 144269 78371 144335 78374
rect 149278 78372 149284 78436
rect 149348 78434 149354 78436
rect 149421 78434 149487 78437
rect 167361 78436 167427 78437
rect 167310 78434 167316 78436
rect 149348 78432 149487 78434
rect 149348 78376 149426 78432
rect 149482 78376 149487 78432
rect 149348 78374 149487 78376
rect 167270 78374 167316 78434
rect 167380 78432 167427 78436
rect 167422 78376 167427 78432
rect 149348 78372 149354 78374
rect 149421 78371 149487 78374
rect 167310 78372 167316 78374
rect 167380 78372 167427 78376
rect 168836 78434 168896 78507
rect 169518 78434 169524 78436
rect 168836 78374 169524 78434
rect 169518 78372 169524 78374
rect 169588 78372 169594 78436
rect 170121 78434 170187 78437
rect 170806 78434 170812 78436
rect 170121 78432 170812 78434
rect 170121 78376 170126 78432
rect 170182 78376 170812 78432
rect 170121 78374 170812 78376
rect 167361 78371 167427 78372
rect 170121 78371 170187 78374
rect 170806 78372 170812 78374
rect 170876 78372 170882 78436
rect 172697 78434 172763 78437
rect 172830 78434 172836 78436
rect 172697 78432 172836 78434
rect 172697 78376 172702 78432
rect 172758 78376 172836 78432
rect 172697 78374 172836 78376
rect 172697 78371 172763 78374
rect 172830 78372 172836 78374
rect 172900 78372 172906 78436
rect 173382 78372 173388 78436
rect 173452 78434 173458 78436
rect 173709 78434 173775 78437
rect 173452 78432 173775 78434
rect 173452 78376 173714 78432
rect 173770 78376 173775 78432
rect 173452 78374 173775 78376
rect 173452 78372 173458 78374
rect 173709 78371 173775 78374
rect 173985 78434 174051 78437
rect 175406 78434 175412 78436
rect 173985 78432 175412 78434
rect 173985 78376 173990 78432
rect 174046 78376 175412 78432
rect 173985 78374 175412 78376
rect 173985 78371 174051 78374
rect 175406 78372 175412 78374
rect 175476 78372 175482 78436
rect 180517 78434 180583 78437
rect 180517 78432 209790 78434
rect 180517 78376 180522 78432
rect 180578 78376 209790 78432
rect 180517 78374 209790 78376
rect 180517 78371 180583 78374
rect 136817 78298 136883 78301
rect 137502 78298 137508 78300
rect 136817 78296 137508 78298
rect 136817 78240 136822 78296
rect 136878 78240 137508 78296
rect 136817 78238 137508 78240
rect 136817 78235 136883 78238
rect 137502 78236 137508 78238
rect 137572 78236 137578 78300
rect 139526 78236 139532 78300
rect 139596 78298 139602 78300
rect 139761 78298 139827 78301
rect 142245 78300 142311 78301
rect 142245 78298 142292 78300
rect 139596 78296 139827 78298
rect 139596 78240 139766 78296
rect 139822 78240 139827 78296
rect 139596 78238 139827 78240
rect 142200 78296 142292 78298
rect 142200 78240 142250 78296
rect 142200 78238 142292 78240
rect 139596 78236 139602 78238
rect 139761 78235 139827 78238
rect 142245 78236 142292 78238
rect 142356 78236 142362 78300
rect 165470 78236 165476 78300
rect 165540 78298 165546 78300
rect 165613 78298 165679 78301
rect 168925 78300 168991 78301
rect 168925 78298 168972 78300
rect 165540 78296 165679 78298
rect 165540 78240 165618 78296
rect 165674 78240 165679 78296
rect 165540 78238 165679 78240
rect 168880 78296 168972 78298
rect 168880 78240 168930 78296
rect 168880 78238 168972 78240
rect 165540 78236 165546 78238
rect 142245 78235 142311 78236
rect 165613 78235 165679 78238
rect 168925 78236 168972 78238
rect 169036 78236 169042 78300
rect 177573 78298 177639 78301
rect 177573 78296 204914 78298
rect 177573 78240 177578 78296
rect 177634 78240 204914 78296
rect 177573 78238 204914 78240
rect 168925 78235 168991 78236
rect 177573 78235 177639 78238
rect 136817 78162 136883 78165
rect 136950 78162 136956 78164
rect 136817 78160 136956 78162
rect 136817 78104 136822 78160
rect 136878 78104 136956 78160
rect 136817 78102 136956 78104
rect 136817 78099 136883 78102
rect 136950 78100 136956 78102
rect 137020 78100 137026 78164
rect 139301 78162 139367 78165
rect 139301 78160 139594 78162
rect 139301 78104 139306 78160
rect 139362 78104 139594 78160
rect 139301 78102 139594 78104
rect 139301 78099 139367 78102
rect 107326 77964 107332 78028
rect 107396 78026 107402 78028
rect 127065 78026 127131 78029
rect 107396 78024 127131 78026
rect 107396 77968 127070 78024
rect 127126 77968 127131 78024
rect 107396 77966 127131 77968
rect 107396 77964 107402 77966
rect 127065 77963 127131 77966
rect 133965 78028 134031 78029
rect 133965 78024 134012 78028
rect 134076 78026 134082 78028
rect 139534 78026 139594 78102
rect 164182 78100 164188 78164
rect 164252 78162 164258 78164
rect 164693 78162 164759 78165
rect 164252 78160 164759 78162
rect 164252 78104 164698 78160
rect 164754 78104 164759 78160
rect 164252 78102 164759 78104
rect 164252 78100 164258 78102
rect 164693 78099 164759 78102
rect 171869 78162 171935 78165
rect 178309 78162 178375 78165
rect 171869 78160 178375 78162
rect 171869 78104 171874 78160
rect 171930 78104 178314 78160
rect 178370 78104 178375 78160
rect 171869 78102 178375 78104
rect 171869 78099 171935 78102
rect 178309 78099 178375 78102
rect 181437 78162 181503 78165
rect 201401 78162 201467 78165
rect 181437 78160 201467 78162
rect 181437 78104 181442 78160
rect 181498 78104 201406 78160
rect 201462 78104 201467 78160
rect 181437 78102 201467 78104
rect 181437 78099 181503 78102
rect 201401 78099 201467 78102
rect 139894 78026 139900 78028
rect 133965 77968 133970 78024
rect 133965 77964 134012 77968
rect 134076 77966 134122 78026
rect 139534 77966 139900 78026
rect 134076 77964 134082 77966
rect 139894 77964 139900 77966
rect 139964 77964 139970 78028
rect 169569 78026 169635 78029
rect 197353 78026 197419 78029
rect 169569 78024 197419 78026
rect 169569 77968 169574 78024
rect 169630 77968 197358 78024
rect 197414 77968 197419 78024
rect 169569 77966 197419 77968
rect 204854 78026 204914 78238
rect 209730 78162 209790 78374
rect 211286 78162 211292 78164
rect 209730 78102 211292 78162
rect 211286 78100 211292 78102
rect 211356 78162 211362 78164
rect 268377 78162 268443 78165
rect 211356 78160 268443 78162
rect 211356 78104 268382 78160
rect 268438 78104 268443 78160
rect 211356 78102 268443 78104
rect 211356 78100 211362 78102
rect 268377 78099 268443 78102
rect 221457 78026 221523 78029
rect 222101 78026 222167 78029
rect 342897 78026 342963 78029
rect 204854 77966 209790 78026
rect 133965 77963 134031 77964
rect 169569 77963 169635 77966
rect 197353 77963 197419 77966
rect 2773 77888 99390 77890
rect 2773 77832 2778 77888
rect 2834 77832 99390 77888
rect 2773 77830 99390 77832
rect 127157 77890 127223 77893
rect 138933 77890 138999 77893
rect 127157 77888 138999 77890
rect 127157 77832 127162 77888
rect 127218 77832 138938 77888
rect 138994 77832 138999 77888
rect 127157 77830 138999 77832
rect 2773 77827 2839 77830
rect 127157 77827 127223 77830
rect 138933 77827 138999 77830
rect 169109 77890 169175 77893
rect 209730 77890 209790 77966
rect 221457 78024 342963 78026
rect 221457 77968 221462 78024
rect 221518 77968 222106 78024
rect 222162 77968 342902 78024
rect 342958 77968 342963 78024
rect 221457 77966 342963 77968
rect 221457 77963 221523 77966
rect 222101 77963 222167 77966
rect 342897 77963 342963 77966
rect 211102 77890 211108 77892
rect 169109 77888 175290 77890
rect 169109 77832 169114 77888
rect 169170 77832 175290 77888
rect 169109 77830 175290 77832
rect 209730 77830 211108 77890
rect 169109 77827 169175 77830
rect 130745 77754 130811 77757
rect 140865 77754 140931 77757
rect 130745 77752 140931 77754
rect 130745 77696 130750 77752
rect 130806 77696 140870 77752
rect 140926 77696 140931 77752
rect 130745 77694 140931 77696
rect 130745 77691 130811 77694
rect 140865 77691 140931 77694
rect 152457 77754 152523 77757
rect 171961 77756 172027 77757
rect 152590 77754 152596 77756
rect 152457 77752 152596 77754
rect 152457 77696 152462 77752
rect 152518 77696 152596 77752
rect 152457 77694 152596 77696
rect 152457 77691 152523 77694
rect 152590 77692 152596 77694
rect 152660 77692 152666 77756
rect 171910 77754 171916 77756
rect 171870 77694 171916 77754
rect 171980 77752 172027 77756
rect 172022 77696 172027 77752
rect 171910 77692 171916 77694
rect 171980 77692 172027 77696
rect 171961 77691 172027 77692
rect 173433 77754 173499 77757
rect 173750 77754 173756 77756
rect 173433 77752 173756 77754
rect 173433 77696 173438 77752
rect 173494 77696 173756 77752
rect 173433 77694 173756 77696
rect 173433 77691 173499 77694
rect 173750 77692 173756 77694
rect 173820 77692 173826 77756
rect 132861 77618 132927 77621
rect 133454 77618 133460 77620
rect 132861 77616 133460 77618
rect 132861 77560 132866 77616
rect 132922 77560 133460 77616
rect 132861 77558 133460 77560
rect 132861 77555 132927 77558
rect 133454 77556 133460 77558
rect 133524 77556 133530 77620
rect 144126 77556 144132 77620
rect 144196 77618 144202 77620
rect 144453 77618 144519 77621
rect 144196 77616 144519 77618
rect 144196 77560 144458 77616
rect 144514 77560 144519 77616
rect 144196 77558 144519 77560
rect 144196 77556 144202 77558
rect 144453 77555 144519 77558
rect 133270 77420 133276 77484
rect 133340 77482 133346 77484
rect 133413 77482 133479 77485
rect 133340 77480 133479 77482
rect 133340 77424 133418 77480
rect 133474 77424 133479 77480
rect 133340 77422 133479 77424
rect 133340 77420 133346 77422
rect 133413 77419 133479 77422
rect 135478 77420 135484 77484
rect 135548 77482 135554 77484
rect 135805 77482 135871 77485
rect 135548 77480 135871 77482
rect 135548 77424 135810 77480
rect 135866 77424 135871 77480
rect 135548 77422 135871 77424
rect 135548 77420 135554 77422
rect 135805 77419 135871 77422
rect 143574 77420 143580 77484
rect 143644 77482 143650 77484
rect 144085 77482 144151 77485
rect 147949 77484 148015 77485
rect 147949 77482 147996 77484
rect 143644 77480 144151 77482
rect 143644 77424 144090 77480
rect 144146 77424 144151 77480
rect 143644 77422 144151 77424
rect 147904 77480 147996 77482
rect 147904 77424 147954 77480
rect 147904 77422 147996 77424
rect 143644 77420 143650 77422
rect 144085 77419 144151 77422
rect 147949 77420 147996 77422
rect 148060 77420 148066 77484
rect 148174 77420 148180 77484
rect 148244 77482 148250 77484
rect 148409 77482 148475 77485
rect 161105 77484 161171 77485
rect 148244 77480 148475 77482
rect 148244 77424 148414 77480
rect 148470 77424 148475 77480
rect 148244 77422 148475 77424
rect 148244 77420 148250 77422
rect 147949 77419 148015 77420
rect 148409 77419 148475 77422
rect 161054 77420 161060 77484
rect 161124 77482 161171 77484
rect 175230 77482 175290 77830
rect 211102 77828 211108 77830
rect 211172 77890 211178 77892
rect 486417 77890 486483 77893
rect 211172 77888 486483 77890
rect 211172 77832 486422 77888
rect 486478 77832 486483 77888
rect 211172 77830 486483 77832
rect 211172 77828 211178 77830
rect 486417 77827 486483 77830
rect 177941 77482 178007 77485
rect 183553 77482 183619 77485
rect 161124 77480 161216 77482
rect 161166 77424 161216 77480
rect 161124 77422 161216 77424
rect 175230 77422 176670 77482
rect 161124 77420 161171 77422
rect 161105 77419 161171 77420
rect 133086 77284 133092 77348
rect 133156 77346 133162 77348
rect 133597 77346 133663 77349
rect 134609 77348 134675 77349
rect 133156 77344 133663 77346
rect 133156 77288 133602 77344
rect 133658 77288 133663 77344
rect 133156 77286 133663 77288
rect 133156 77284 133162 77286
rect 133597 77283 133663 77286
rect 134558 77284 134564 77348
rect 134628 77346 134675 77348
rect 142429 77346 142495 77349
rect 142838 77346 142844 77348
rect 134628 77344 134720 77346
rect 134670 77288 134720 77344
rect 134628 77286 134720 77288
rect 142429 77344 142844 77346
rect 142429 77288 142434 77344
rect 142490 77288 142844 77344
rect 142429 77286 142844 77288
rect 134628 77284 134675 77286
rect 134609 77283 134675 77284
rect 142429 77283 142495 77286
rect 142838 77284 142844 77286
rect 142908 77284 142914 77348
rect 142981 77346 143047 77349
rect 143206 77346 143212 77348
rect 142981 77344 143212 77346
rect 142981 77288 142986 77344
rect 143042 77288 143212 77344
rect 142981 77286 143212 77288
rect 142981 77283 143047 77286
rect 143206 77284 143212 77286
rect 143276 77284 143282 77348
rect 143993 77346 144059 77349
rect 144310 77346 144316 77348
rect 143993 77344 144316 77346
rect 143993 77288 143998 77344
rect 144054 77288 144316 77344
rect 143993 77286 144316 77288
rect 143993 77283 144059 77286
rect 144310 77284 144316 77286
rect 144380 77284 144386 77348
rect 147990 77284 147996 77348
rect 148060 77346 148066 77348
rect 148685 77346 148751 77349
rect 152549 77346 152615 77349
rect 153101 77346 153167 77349
rect 148060 77344 148751 77346
rect 148060 77288 148690 77344
rect 148746 77288 148751 77344
rect 148060 77286 148751 77288
rect 148060 77284 148066 77286
rect 148685 77283 148751 77286
rect 151770 77344 153167 77346
rect 151770 77288 152554 77344
rect 152610 77288 153106 77344
rect 153162 77288 153167 77344
rect 151770 77286 153167 77288
rect 176610 77346 176670 77422
rect 177941 77480 183619 77482
rect 177941 77424 177946 77480
rect 178002 77424 183558 77480
rect 183614 77424 183619 77480
rect 177941 77422 183619 77424
rect 177941 77419 178007 77422
rect 183553 77419 183619 77422
rect 222101 77346 222167 77349
rect 176610 77344 222167 77346
rect 176610 77288 222106 77344
rect 222162 77288 222167 77344
rect 176610 77286 222167 77288
rect 110822 77148 110828 77212
rect 110892 77210 110898 77212
rect 111241 77210 111307 77213
rect 110892 77208 111307 77210
rect 110892 77152 111246 77208
rect 111302 77152 111307 77208
rect 110892 77150 111307 77152
rect 110892 77148 110898 77150
rect 111241 77147 111307 77150
rect 117998 77148 118004 77212
rect 118068 77210 118074 77212
rect 151770 77210 151830 77286
rect 152549 77283 152615 77286
rect 153101 77283 153167 77286
rect 222101 77283 222167 77286
rect 118068 77150 151830 77210
rect 152181 77210 152247 77213
rect 152774 77210 152780 77212
rect 152181 77208 152780 77210
rect 152181 77152 152186 77208
rect 152242 77152 152780 77208
rect 152181 77150 152780 77152
rect 118068 77148 118074 77150
rect 152181 77147 152247 77150
rect 152774 77148 152780 77150
rect 152844 77148 152850 77212
rect 154246 77148 154252 77212
rect 154316 77210 154322 77212
rect 154665 77210 154731 77213
rect 154316 77208 154731 77210
rect 154316 77152 154670 77208
rect 154726 77152 154731 77208
rect 154316 77150 154731 77152
rect 154316 77148 154322 77150
rect 154665 77147 154731 77150
rect 162526 77148 162532 77212
rect 162596 77210 162602 77212
rect 162761 77210 162827 77213
rect 162596 77208 162827 77210
rect 162596 77152 162766 77208
rect 162822 77152 162827 77208
rect 162596 77150 162827 77152
rect 162596 77148 162602 77150
rect 162761 77147 162827 77150
rect 118182 77012 118188 77076
rect 118252 77074 118258 77076
rect 143349 77074 143415 77077
rect 143758 77074 143764 77076
rect 118252 77014 138030 77074
rect 118252 77012 118258 77014
rect 98729 76938 98795 76941
rect 128629 76938 128695 76941
rect 98729 76936 128695 76938
rect 98729 76880 98734 76936
rect 98790 76880 128634 76936
rect 128690 76880 128695 76936
rect 98729 76878 128695 76880
rect 98729 76875 98795 76878
rect 128629 76875 128695 76878
rect 103053 76802 103119 76805
rect 137461 76802 137527 76805
rect 99330 76800 137527 76802
rect 99330 76744 103058 76800
rect 103114 76744 137466 76800
rect 137522 76744 137527 76800
rect 99330 76742 137527 76744
rect 137970 76802 138030 77014
rect 143349 77072 143764 77074
rect 143349 77016 143354 77072
rect 143410 77016 143764 77072
rect 143349 77014 143764 77016
rect 143349 77011 143415 77014
rect 143758 77012 143764 77014
rect 143828 77012 143834 77076
rect 160829 77074 160895 77077
rect 218329 77074 218395 77077
rect 218513 77074 218579 77077
rect 160829 77072 218579 77074
rect 160829 77016 160834 77072
rect 160890 77016 218334 77072
rect 218390 77016 218518 77072
rect 218574 77016 218579 77072
rect 160829 77014 218579 77016
rect 160829 77011 160895 77014
rect 218329 77011 218395 77014
rect 218513 77011 218579 77014
rect 143758 76876 143764 76940
rect 143828 76938 143834 76940
rect 144729 76938 144795 76941
rect 143828 76936 144795 76938
rect 143828 76880 144734 76936
rect 144790 76880 144795 76936
rect 143828 76878 144795 76880
rect 143828 76876 143834 76878
rect 144729 76875 144795 76878
rect 164785 76938 164851 76941
rect 165286 76938 165292 76940
rect 164785 76936 165292 76938
rect 164785 76880 164790 76936
rect 164846 76880 165292 76936
rect 164785 76878 165292 76880
rect 164785 76875 164851 76878
rect 165286 76876 165292 76878
rect 165356 76876 165362 76940
rect 170070 76876 170076 76940
rect 170140 76938 170146 76940
rect 170990 76938 170996 76940
rect 170140 76878 170996 76938
rect 170140 76876 170146 76878
rect 170990 76876 170996 76878
rect 171060 76876 171066 76940
rect 174486 76876 174492 76940
rect 174556 76938 174562 76940
rect 174813 76938 174879 76941
rect 174556 76936 174879 76938
rect 174556 76880 174818 76936
rect 174874 76880 174879 76936
rect 174556 76878 174879 76880
rect 174556 76876 174562 76878
rect 174813 76875 174879 76878
rect 176101 76940 176167 76941
rect 176101 76936 176148 76940
rect 176212 76938 176218 76940
rect 178217 76938 178283 76941
rect 210509 76938 210575 76941
rect 211061 76938 211127 76941
rect 176101 76880 176106 76936
rect 176101 76876 176148 76880
rect 176212 76878 176258 76938
rect 178217 76936 211127 76938
rect 178217 76880 178222 76936
rect 178278 76880 210514 76936
rect 210570 76880 211066 76936
rect 211122 76880 211127 76936
rect 178217 76878 211127 76880
rect 176212 76876 176218 76878
rect 176101 76875 176167 76876
rect 178217 76875 178283 76878
rect 210509 76875 210575 76878
rect 211061 76875 211127 76878
rect 217961 76938 218027 76941
rect 218513 76938 218579 76941
rect 247677 76938 247743 76941
rect 217961 76936 247743 76938
rect 217961 76880 217966 76936
rect 218022 76880 218518 76936
rect 218574 76880 247682 76936
rect 247738 76880 247743 76936
rect 217961 76878 247743 76880
rect 217961 76875 218027 76878
rect 218513 76875 218579 76878
rect 247677 76875 247743 76878
rect 152641 76802 152707 76805
rect 260833 76802 260899 76805
rect 137970 76800 260899 76802
rect 137970 76744 152646 76800
rect 152702 76744 260838 76800
rect 260894 76744 260899 76800
rect 137970 76742 260899 76744
rect 66253 76666 66319 76669
rect 99330 76666 99390 76742
rect 103053 76739 103119 76742
rect 137461 76739 137527 76742
rect 152641 76739 152707 76742
rect 260833 76739 260899 76742
rect 66253 76664 99390 76666
rect 66253 76608 66258 76664
rect 66314 76608 99390 76664
rect 66253 76606 99390 76608
rect 66253 76603 66319 76606
rect 133822 76604 133828 76668
rect 133892 76666 133898 76668
rect 134701 76666 134767 76669
rect 133892 76664 134767 76666
rect 133892 76608 134706 76664
rect 134762 76608 134767 76664
rect 133892 76606 134767 76608
rect 133892 76604 133898 76606
rect 134701 76603 134767 76606
rect 170397 76666 170463 76669
rect 197486 76666 197492 76668
rect 170397 76664 197492 76666
rect 170397 76608 170402 76664
rect 170458 76608 197492 76664
rect 170397 76606 197492 76608
rect 170397 76603 170463 76606
rect 197486 76604 197492 76606
rect 197556 76604 197562 76668
rect 218329 76666 218395 76669
rect 367093 76666 367159 76669
rect 218329 76664 367159 76666
rect 218329 76608 218334 76664
rect 218390 76608 367098 76664
rect 367154 76608 367159 76664
rect 218329 76606 367159 76608
rect 218329 76603 218395 76606
rect 367093 76603 367159 76606
rect 13077 76530 13143 76533
rect 98729 76530 98795 76533
rect 13077 76528 98795 76530
rect 13077 76472 13082 76528
rect 13138 76472 98734 76528
rect 98790 76472 98795 76528
rect 13077 76470 98795 76472
rect 13077 76467 13143 76470
rect 98729 76467 98795 76470
rect 162669 76532 162735 76533
rect 162669 76528 162716 76532
rect 162780 76530 162786 76532
rect 170121 76530 170187 76533
rect 170254 76530 170260 76532
rect 162669 76472 162674 76528
rect 162669 76468 162716 76472
rect 162780 76470 162826 76530
rect 170121 76528 170260 76530
rect 170121 76472 170126 76528
rect 170182 76472 170260 76528
rect 170121 76470 170260 76472
rect 162780 76468 162786 76470
rect 162669 76467 162735 76468
rect 170121 76467 170187 76470
rect 170254 76468 170260 76470
rect 170324 76468 170330 76532
rect 170489 76530 170555 76533
rect 170622 76530 170628 76532
rect 170489 76528 170628 76530
rect 170489 76472 170494 76528
rect 170550 76472 170628 76528
rect 170489 76470 170628 76472
rect 170489 76467 170555 76470
rect 170622 76468 170628 76470
rect 170692 76468 170698 76532
rect 171593 76530 171659 76533
rect 172145 76532 172211 76533
rect 172329 76532 172395 76533
rect 171726 76530 171732 76532
rect 171593 76528 171732 76530
rect 171593 76472 171598 76528
rect 171654 76472 171732 76528
rect 171593 76470 171732 76472
rect 171593 76467 171659 76470
rect 171726 76468 171732 76470
rect 171796 76468 171802 76532
rect 172094 76530 172100 76532
rect 172054 76470 172100 76530
rect 172164 76528 172211 76532
rect 172206 76472 172211 76528
rect 172094 76468 172100 76470
rect 172164 76468 172211 76472
rect 172278 76468 172284 76532
rect 172348 76530 172395 76532
rect 174721 76530 174787 76533
rect 175089 76532 175155 76533
rect 174854 76530 174860 76532
rect 172348 76528 172440 76530
rect 172390 76472 172440 76528
rect 172348 76470 172440 76472
rect 174721 76528 174860 76530
rect 174721 76472 174726 76528
rect 174782 76472 174860 76528
rect 174721 76470 174860 76472
rect 172348 76468 172395 76470
rect 172145 76467 172211 76468
rect 172329 76467 172395 76468
rect 174721 76467 174787 76470
rect 174854 76468 174860 76470
rect 174924 76468 174930 76532
rect 175038 76530 175044 76532
rect 174998 76470 175044 76530
rect 175108 76528 175155 76532
rect 175150 76472 175155 76528
rect 175038 76468 175044 76470
rect 175108 76468 175155 76472
rect 175089 76467 175155 76468
rect 176193 76530 176259 76533
rect 176561 76530 176627 76533
rect 200982 76530 200988 76532
rect 176193 76528 200988 76530
rect 176193 76472 176198 76528
rect 176254 76472 176566 76528
rect 176622 76472 200988 76528
rect 176193 76470 200988 76472
rect 176193 76467 176259 76470
rect 176561 76467 176627 76470
rect 200982 76468 200988 76470
rect 201052 76468 201058 76532
rect 211061 76530 211127 76533
rect 552657 76530 552723 76533
rect 211061 76528 552723 76530
rect 211061 76472 211066 76528
rect 211122 76472 552662 76528
rect 552718 76472 552723 76528
rect 211061 76470 552723 76472
rect 211061 76467 211127 76470
rect 552657 76467 552723 76470
rect 154481 76394 154547 76397
rect 218513 76394 218579 76397
rect 154481 76392 218579 76394
rect 154481 76336 154486 76392
rect 154542 76336 218518 76392
rect 218574 76336 218579 76392
rect 154481 76334 218579 76336
rect 154481 76331 154547 76334
rect 218513 76331 218579 76334
rect 139669 76258 139735 76261
rect 140630 76258 140636 76260
rect 139669 76256 140636 76258
rect 139669 76200 139674 76256
rect 139730 76200 140636 76256
rect 139669 76198 140636 76200
rect 139669 76195 139735 76198
rect 140630 76196 140636 76198
rect 140700 76196 140706 76260
rect 145373 76258 145439 76261
rect 145598 76258 145604 76260
rect 145373 76256 145604 76258
rect 145373 76200 145378 76256
rect 145434 76200 145604 76256
rect 145373 76198 145604 76200
rect 145373 76195 145439 76198
rect 145598 76196 145604 76198
rect 145668 76196 145674 76260
rect 146886 76196 146892 76260
rect 146956 76258 146962 76260
rect 147489 76258 147555 76261
rect 146956 76256 147555 76258
rect 146956 76200 147494 76256
rect 147550 76200 147555 76256
rect 146956 76198 147555 76200
rect 146956 76196 146962 76198
rect 147489 76195 147555 76198
rect 176285 76258 176351 76261
rect 176510 76258 176516 76260
rect 176285 76256 176516 76258
rect 176285 76200 176290 76256
rect 176346 76200 176516 76256
rect 176285 76198 176516 76200
rect 176285 76195 176351 76198
rect 176510 76196 176516 76198
rect 176580 76196 176586 76260
rect 138013 76124 138079 76125
rect 138013 76120 138060 76124
rect 138124 76122 138130 76124
rect 138013 76064 138018 76120
rect 138013 76060 138060 76064
rect 138124 76062 138170 76122
rect 138124 76060 138130 76062
rect 138238 76060 138244 76124
rect 138308 76122 138314 76124
rect 138657 76122 138723 76125
rect 138308 76120 138723 76122
rect 138308 76064 138662 76120
rect 138718 76064 138723 76120
rect 138308 76062 138723 76064
rect 138308 76060 138314 76062
rect 138013 76059 138079 76060
rect 138657 76059 138723 76062
rect 170438 76060 170444 76124
rect 170508 76122 170514 76124
rect 171041 76122 171107 76125
rect 170508 76120 171107 76122
rect 170508 76064 171046 76120
rect 171102 76064 171107 76120
rect 170508 76062 171107 76064
rect 170508 76060 170514 76062
rect 171041 76059 171107 76062
rect 163630 75924 163636 75988
rect 163700 75986 163706 75988
rect 163865 75986 163931 75989
rect 165337 75988 165403 75989
rect 165286 75986 165292 75988
rect 163700 75984 163931 75986
rect 163700 75928 163870 75984
rect 163926 75928 163931 75984
rect 163700 75926 163931 75928
rect 165246 75926 165292 75986
rect 165356 75984 165403 75988
rect 165398 75928 165403 75984
rect 163700 75924 163706 75926
rect 163865 75923 163931 75926
rect 165286 75924 165292 75926
rect 165356 75924 165403 75928
rect 165654 75924 165660 75988
rect 165724 75986 165730 75988
rect 165797 75986 165863 75989
rect 165724 75984 165863 75986
rect 165724 75928 165802 75984
rect 165858 75928 165863 75984
rect 165724 75926 165863 75928
rect 165724 75924 165730 75926
rect 165337 75923 165403 75924
rect 165797 75923 165863 75926
rect 166993 75986 167059 75989
rect 167729 75988 167795 75989
rect 167310 75986 167316 75988
rect 166993 75984 167316 75986
rect 166993 75928 166998 75984
rect 167054 75928 167316 75984
rect 166993 75926 167316 75928
rect 166993 75923 167059 75926
rect 167310 75924 167316 75926
rect 167380 75924 167386 75988
rect 167678 75986 167684 75988
rect 167638 75926 167684 75986
rect 167748 75984 167795 75988
rect 167790 75928 167795 75984
rect 167678 75924 167684 75926
rect 167748 75924 167795 75928
rect 167729 75923 167795 75924
rect 122741 75850 122807 75853
rect 123109 75850 123175 75853
rect 122741 75848 123175 75850
rect 122741 75792 122746 75848
rect 122802 75792 123114 75848
rect 123170 75792 123175 75848
rect 122741 75790 123175 75792
rect 122741 75787 122807 75790
rect 123109 75787 123175 75790
rect 138749 75850 138815 75853
rect 138974 75850 138980 75852
rect 138749 75848 138980 75850
rect 138749 75792 138754 75848
rect 138810 75792 138980 75848
rect 138749 75790 138980 75792
rect 138749 75787 138815 75790
rect 138974 75788 138980 75790
rect 139044 75788 139050 75852
rect 171542 75788 171548 75852
rect 171612 75850 171618 75852
rect 172237 75850 172303 75853
rect 171612 75848 172303 75850
rect 171612 75792 172242 75848
rect 172298 75792 172303 75848
rect 171612 75790 172303 75792
rect 171612 75788 171618 75790
rect 172237 75787 172303 75790
rect 205541 75852 205607 75853
rect 205541 75848 205588 75852
rect 205652 75850 205658 75852
rect 205541 75792 205546 75848
rect 205541 75788 205588 75792
rect 205652 75790 205698 75850
rect 205652 75788 205658 75790
rect 205766 75788 205772 75852
rect 205836 75850 205842 75852
rect 206277 75850 206343 75853
rect 205836 75848 206343 75850
rect 205836 75792 206282 75848
rect 206338 75792 206343 75848
rect 205836 75790 206343 75792
rect 205836 75788 205842 75790
rect 205541 75787 205607 75788
rect 206277 75787 206343 75790
rect 114461 75714 114527 75717
rect 147254 75714 147260 75716
rect 114461 75712 147260 75714
rect 114461 75656 114466 75712
rect 114522 75656 147260 75712
rect 114461 75654 147260 75656
rect 114461 75651 114527 75654
rect 147254 75652 147260 75654
rect 147324 75652 147330 75716
rect 173249 75714 173315 75717
rect 173249 75712 205834 75714
rect 173249 75656 173254 75712
rect 173310 75656 205834 75712
rect 173249 75654 205834 75656
rect 173249 75651 173315 75654
rect 112713 75578 112779 75581
rect 175181 75580 175247 75581
rect 145414 75578 145420 75580
rect 112713 75576 145420 75578
rect 112713 75520 112718 75576
rect 112774 75520 145420 75576
rect 112713 75518 145420 75520
rect 112713 75515 112779 75518
rect 145414 75516 145420 75518
rect 145484 75516 145490 75580
rect 175181 75578 175228 75580
rect 175136 75576 175228 75578
rect 175136 75520 175186 75576
rect 175136 75518 175228 75520
rect 175181 75516 175228 75518
rect 175292 75516 175298 75580
rect 176101 75578 176167 75581
rect 203374 75578 203380 75580
rect 176101 75576 203380 75578
rect 176101 75520 176106 75576
rect 176162 75520 203380 75576
rect 176101 75518 203380 75520
rect 175181 75515 175247 75516
rect 176101 75515 176167 75518
rect 203374 75516 203380 75518
rect 203444 75516 203450 75580
rect 115197 75442 115263 75445
rect 147581 75442 147647 75445
rect 196198 75442 196204 75444
rect 115197 75440 151830 75442
rect 115197 75384 115202 75440
rect 115258 75384 147586 75440
rect 147642 75384 151830 75440
rect 115197 75382 151830 75384
rect 115197 75379 115263 75382
rect 147581 75379 147647 75382
rect 118417 75306 118483 75309
rect 146477 75306 146543 75309
rect 118417 75304 146543 75306
rect 118417 75248 118422 75304
rect 118478 75248 146482 75304
rect 146538 75248 146543 75304
rect 118417 75246 146543 75248
rect 118417 75243 118483 75246
rect 146477 75243 146543 75246
rect 7557 75170 7623 75173
rect 97206 75170 97212 75172
rect 7557 75168 97212 75170
rect 7557 75112 7562 75168
rect 7618 75112 97212 75168
rect 7557 75110 97212 75112
rect 7557 75107 7623 75110
rect 97206 75108 97212 75110
rect 97276 75170 97282 75172
rect 97349 75170 97415 75173
rect 97276 75168 97415 75170
rect 97276 75112 97354 75168
rect 97410 75112 97415 75168
rect 97276 75110 97415 75112
rect 97276 75108 97282 75110
rect 97349 75107 97415 75110
rect 111149 75170 111215 75173
rect 129733 75170 129799 75173
rect 130929 75170 130995 75173
rect 111149 75168 130995 75170
rect 111149 75112 111154 75168
rect 111210 75112 129738 75168
rect 129794 75112 130934 75168
rect 130990 75112 130995 75168
rect 111149 75110 130995 75112
rect 111149 75107 111215 75110
rect 129733 75107 129799 75110
rect 130929 75107 130995 75110
rect 138105 75170 138171 75173
rect 138606 75170 138612 75172
rect 138105 75168 138612 75170
rect 138105 75112 138110 75168
rect 138166 75112 138612 75168
rect 138105 75110 138612 75112
rect 138105 75107 138171 75110
rect 138606 75108 138612 75110
rect 138676 75108 138682 75172
rect 140814 75108 140820 75172
rect 140884 75170 140890 75172
rect 141325 75170 141391 75173
rect 140884 75168 141391 75170
rect 140884 75112 141330 75168
rect 141386 75112 141391 75168
rect 140884 75110 141391 75112
rect 140884 75108 140890 75110
rect 141325 75107 141391 75110
rect 145414 75108 145420 75172
rect 145484 75170 145490 75172
rect 146201 75170 146267 75173
rect 145484 75168 146267 75170
rect 145484 75112 146206 75168
rect 146262 75112 146267 75168
rect 145484 75110 146267 75112
rect 151770 75170 151830 75382
rect 171918 75382 196204 75442
rect 168925 75306 168991 75309
rect 169477 75306 169543 75309
rect 171918 75306 171978 75382
rect 196198 75380 196204 75382
rect 196268 75380 196274 75444
rect 168925 75304 171978 75306
rect 168925 75248 168930 75304
rect 168986 75248 169482 75304
rect 169538 75248 171978 75304
rect 168925 75246 171978 75248
rect 172237 75306 172303 75309
rect 199142 75306 199148 75308
rect 172237 75304 199148 75306
rect 172237 75248 172242 75304
rect 172298 75248 199148 75304
rect 172237 75246 199148 75248
rect 168925 75243 168991 75246
rect 169477 75243 169543 75246
rect 172237 75243 172303 75246
rect 199142 75244 199148 75246
rect 199212 75244 199218 75308
rect 194041 75170 194107 75173
rect 151770 75168 194107 75170
rect 151770 75112 194046 75168
rect 194102 75112 194107 75168
rect 151770 75110 194107 75112
rect 205774 75170 205834 75654
rect 207105 75306 207171 75309
rect 207473 75306 207539 75309
rect 493317 75306 493383 75309
rect 207105 75304 493383 75306
rect 207105 75248 207110 75304
rect 207166 75248 207478 75304
rect 207534 75248 493322 75304
rect 493378 75248 493383 75304
rect 207105 75246 493383 75248
rect 207105 75243 207171 75246
rect 207473 75243 207539 75246
rect 493317 75243 493383 75246
rect 207381 75170 207447 75173
rect 521653 75170 521719 75173
rect 205774 75168 521719 75170
rect 205774 75112 207386 75168
rect 207442 75112 521658 75168
rect 521714 75112 521719 75168
rect 205774 75110 521719 75112
rect 145484 75108 145490 75110
rect 146201 75107 146267 75110
rect 194041 75107 194107 75110
rect 207381 75107 207447 75110
rect 521653 75107 521719 75110
rect 144310 74972 144316 75036
rect 144380 75034 144386 75036
rect 144545 75034 144611 75037
rect 144380 75032 144611 75034
rect 144380 74976 144550 75032
rect 144606 74976 144611 75032
rect 144380 74974 144611 74976
rect 144380 74972 144386 74974
rect 144545 74971 144611 74974
rect 178033 75034 178099 75037
rect 207105 75034 207171 75037
rect 178033 75032 207171 75034
rect 178033 74976 178038 75032
rect 178094 74976 207110 75032
rect 207166 74976 207171 75032
rect 178033 74974 207171 74976
rect 178033 74971 178099 74974
rect 207105 74971 207171 74974
rect 115606 74836 115612 74900
rect 115676 74898 115682 74900
rect 176193 74898 176259 74901
rect 177297 74898 177363 74901
rect 115676 74838 138030 74898
rect 115676 74836 115682 74838
rect 137970 74762 138030 74838
rect 176193 74896 177363 74898
rect 176193 74840 176198 74896
rect 176254 74840 177302 74896
rect 177358 74840 177363 74896
rect 176193 74838 177363 74840
rect 176193 74835 176259 74838
rect 177297 74835 177363 74838
rect 152917 74762 152983 74765
rect 137970 74760 152983 74762
rect 137970 74704 152922 74760
rect 152978 74704 152983 74760
rect 137970 74702 152983 74704
rect 152917 74699 152983 74702
rect 112662 74564 112668 74628
rect 112732 74626 112738 74628
rect 113265 74626 113331 74629
rect 112732 74624 113331 74626
rect 112732 74568 113270 74624
rect 113326 74568 113331 74624
rect 112732 74566 113331 74568
rect 112732 74564 112738 74566
rect 113265 74563 113331 74566
rect 119838 74428 119844 74492
rect 119908 74490 119914 74492
rect 154021 74490 154087 74493
rect 154481 74490 154547 74493
rect 119908 74488 154547 74490
rect 119908 74432 154026 74488
rect 154082 74432 154486 74488
rect 154542 74432 154547 74488
rect 119908 74430 154547 74432
rect 119908 74428 119914 74430
rect 154021 74427 154087 74430
rect 154481 74427 154547 74430
rect 118366 74292 118372 74356
rect 118436 74354 118442 74356
rect 118436 74294 151002 74354
rect 118436 74292 118442 74294
rect 116669 74218 116735 74221
rect 149462 74218 149468 74220
rect 116669 74216 149468 74218
rect 116669 74160 116674 74216
rect 116730 74160 149468 74216
rect 116669 74158 149468 74160
rect 116669 74155 116735 74158
rect 149462 74156 149468 74158
rect 149532 74218 149538 74220
rect 149830 74218 149836 74220
rect 149532 74158 149836 74218
rect 149532 74156 149538 74158
rect 149830 74156 149836 74158
rect 149900 74156 149906 74220
rect 117681 74082 117747 74085
rect 150942 74082 151002 74294
rect 152774 74292 152780 74356
rect 152844 74354 152850 74356
rect 218145 74354 218211 74357
rect 152844 74352 218211 74354
rect 152844 74296 218150 74352
rect 218206 74296 218211 74352
rect 152844 74294 218211 74296
rect 152844 74292 152850 74294
rect 218145 74291 218211 74294
rect 151118 74156 151124 74220
rect 151188 74218 151194 74220
rect 215753 74218 215819 74221
rect 151188 74216 219450 74218
rect 151188 74160 215758 74216
rect 215814 74160 219450 74216
rect 151188 74158 219450 74160
rect 151188 74156 151194 74158
rect 215753 74155 215819 74158
rect 152549 74082 152615 74085
rect 176285 74082 176351 74085
rect 204897 74082 204963 74085
rect 117681 74080 138030 74082
rect 117681 74024 117686 74080
rect 117742 74024 138030 74080
rect 117681 74022 138030 74024
rect 150942 74080 157350 74082
rect 150942 74024 152554 74080
rect 152610 74024 157350 74080
rect 150942 74022 157350 74024
rect 117681 74019 117747 74022
rect 54477 73946 54543 73949
rect 106273 73946 106339 73949
rect 106774 73946 106780 73948
rect 54477 73944 106780 73946
rect 54477 73888 54482 73944
rect 54538 73888 106278 73944
rect 106334 73888 106780 73944
rect 54477 73886 106780 73888
rect 54477 73883 54543 73886
rect 106273 73883 106339 73886
rect 106774 73884 106780 73886
rect 106844 73884 106850 73948
rect 137970 73946 138030 74022
rect 152549 74019 152615 74022
rect 149278 73946 149284 73948
rect 137970 73886 149284 73946
rect 149278 73884 149284 73886
rect 149348 73884 149354 73948
rect 14457 73810 14523 73813
rect 103094 73810 103100 73812
rect 14457 73808 103100 73810
rect 14457 73752 14462 73808
rect 14518 73752 103100 73808
rect 14457 73750 103100 73752
rect 14457 73747 14523 73750
rect 103094 73748 103100 73750
rect 103164 73810 103170 73812
rect 130377 73810 130443 73813
rect 103164 73808 130443 73810
rect 103164 73752 130382 73808
rect 130438 73752 130443 73808
rect 103164 73750 130443 73752
rect 103164 73748 103170 73750
rect 130377 73747 130443 73750
rect 142337 73810 142403 73813
rect 143022 73810 143028 73812
rect 142337 73808 143028 73810
rect 142337 73752 142342 73808
rect 142398 73752 143028 73808
rect 142337 73750 143028 73752
rect 142337 73747 142403 73750
rect 143022 73748 143028 73750
rect 143092 73748 143098 73812
rect 157290 73810 157350 74022
rect 176285 74080 204963 74082
rect 176285 74024 176290 74080
rect 176346 74024 204902 74080
rect 204958 74024 204963 74080
rect 176285 74022 204963 74024
rect 219390 74082 219450 74158
rect 237373 74082 237439 74085
rect 219390 74080 237439 74082
rect 219390 74024 237378 74080
rect 237434 74024 237439 74080
rect 219390 74022 237439 74024
rect 176285 74019 176351 74022
rect 204897 74019 204963 74022
rect 237373 74019 237439 74022
rect 218145 73946 218211 73949
rect 255313 73946 255379 73949
rect 218145 73944 255379 73946
rect 218145 73888 218150 73944
rect 218206 73888 255318 73944
rect 255374 73888 255379 73944
rect 218145 73886 255379 73888
rect 218145 73883 218211 73886
rect 255313 73883 255379 73886
rect 261477 73810 261543 73813
rect 157290 73808 261543 73810
rect 157290 73752 261482 73808
rect 261538 73752 261543 73808
rect 157290 73750 261543 73752
rect 261477 73747 261543 73750
rect 154430 73612 154436 73676
rect 154500 73674 154506 73676
rect 221273 73674 221339 73677
rect 154500 73672 221339 73674
rect 154500 73616 221278 73672
rect 221334 73616 221339 73672
rect 154500 73614 221339 73616
rect 154500 73612 154506 73614
rect 221273 73611 221339 73614
rect 221273 73266 221339 73269
rect 224217 73266 224283 73269
rect 221273 73264 224283 73266
rect 221273 73208 221278 73264
rect 221334 73208 224222 73264
rect 224278 73208 224283 73264
rect 221273 73206 224283 73208
rect 221273 73203 221339 73206
rect 224217 73203 224283 73206
rect 104709 73130 104775 73133
rect 131757 73130 131823 73133
rect 151997 73130 152063 73133
rect 152549 73130 152615 73133
rect 104709 73128 131823 73130
rect 104709 73072 104714 73128
rect 104770 73072 131762 73128
rect 131818 73072 131823 73128
rect 104709 73070 131823 73072
rect 104709 73067 104775 73070
rect 131757 73067 131823 73070
rect 147630 73128 152615 73130
rect 147630 73072 152002 73128
rect 152058 73072 152554 73128
rect 152610 73072 152615 73128
rect 147630 73070 152615 73072
rect 99925 72994 99991 72997
rect 130469 72994 130535 72997
rect 99330 72992 130535 72994
rect 99330 72936 99930 72992
rect 99986 72936 130474 72992
rect 130530 72936 130535 72992
rect 99330 72934 130535 72936
rect 8293 72450 8359 72453
rect 99330 72450 99390 72934
rect 99925 72931 99991 72934
rect 130469 72931 130535 72934
rect 120625 72858 120691 72861
rect 147630 72858 147690 73070
rect 151997 73067 152063 73070
rect 152549 73067 152615 73070
rect 157190 73068 157196 73132
rect 157260 73130 157266 73132
rect 220997 73130 221063 73133
rect 157260 73128 229110 73130
rect 157260 73072 221002 73128
rect 221058 73072 229110 73128
rect 157260 73070 229110 73072
rect 157260 73068 157266 73070
rect 220997 73067 221063 73070
rect 158478 72932 158484 72996
rect 158548 72994 158554 72996
rect 219617 72994 219683 72997
rect 158548 72992 219683 72994
rect 158548 72936 219622 72992
rect 219678 72936 219683 72992
rect 158548 72934 219683 72936
rect 158548 72932 158554 72934
rect 120625 72856 147690 72858
rect 120625 72800 120630 72856
rect 120686 72800 147690 72856
rect 120625 72798 147690 72800
rect 174261 72858 174327 72861
rect 174445 72858 174511 72861
rect 175917 72858 175983 72861
rect 176377 72858 176443 72861
rect 210325 72858 210391 72861
rect 174261 72856 175106 72858
rect 174261 72800 174266 72856
rect 174322 72800 174450 72856
rect 174506 72800 175106 72856
rect 174261 72798 175106 72800
rect 120625 72795 120691 72798
rect 174261 72795 174327 72798
rect 174445 72795 174511 72798
rect 112437 72724 112503 72725
rect 112437 72720 112484 72724
rect 112548 72722 112554 72724
rect 118233 72722 118299 72725
rect 148358 72722 148364 72724
rect 112437 72664 112442 72720
rect 112437 72660 112484 72664
rect 112548 72662 112594 72722
rect 118233 72720 148364 72722
rect 118233 72664 118238 72720
rect 118294 72664 148364 72720
rect 118233 72662 148364 72664
rect 112548 72660 112554 72662
rect 112437 72659 112503 72660
rect 118233 72659 118299 72662
rect 148358 72660 148364 72662
rect 148428 72722 148434 72724
rect 148726 72722 148732 72724
rect 148428 72662 148732 72722
rect 148428 72660 148434 72662
rect 148726 72660 148732 72662
rect 148796 72660 148802 72724
rect 175046 72722 175106 72798
rect 175917 72856 210391 72858
rect 175917 72800 175922 72856
rect 175978 72800 176382 72856
rect 176438 72800 210330 72856
rect 210386 72800 210391 72856
rect 175917 72798 210391 72800
rect 175917 72795 175983 72798
rect 176377 72795 176443 72798
rect 210325 72795 210391 72798
rect 208761 72722 208827 72725
rect 175046 72720 208827 72722
rect 175046 72664 208766 72720
rect 208822 72664 208827 72720
rect 175046 72662 208827 72664
rect 208761 72659 208827 72662
rect 104617 72586 104683 72589
rect 176193 72586 176259 72589
rect 176469 72586 176535 72589
rect 207933 72586 207999 72589
rect 104617 72584 122850 72586
rect 104617 72528 104622 72584
rect 104678 72528 122850 72584
rect 104617 72526 122850 72528
rect 104617 72523 104683 72526
rect 8293 72448 99390 72450
rect 8293 72392 8298 72448
rect 8354 72392 99390 72448
rect 8293 72390 99390 72392
rect 122790 72450 122850 72526
rect 176193 72584 207999 72586
rect 176193 72528 176198 72584
rect 176254 72528 176474 72584
rect 176530 72528 207938 72584
rect 207994 72528 207999 72584
rect 176193 72526 207999 72528
rect 176193 72523 176259 72526
rect 176469 72523 176535 72526
rect 207933 72523 207999 72526
rect 133965 72450 134031 72453
rect 122790 72448 134031 72450
rect 122790 72392 133970 72448
rect 134026 72392 134031 72448
rect 122790 72390 134031 72392
rect 8293 72387 8359 72390
rect 133965 72387 134031 72390
rect 169109 72450 169175 72453
rect 192477 72450 192543 72453
rect 169109 72448 192543 72450
rect 169109 72392 169114 72448
rect 169170 72392 192482 72448
rect 192538 72392 192543 72448
rect 169109 72390 192543 72392
rect 219390 72450 219450 72934
rect 219617 72931 219683 72934
rect 229050 72586 229110 73070
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect 318793 72586 318859 72589
rect 229050 72584 318859 72586
rect 229050 72528 318798 72584
rect 318854 72528 318859 72584
rect 229050 72526 318859 72528
rect 318793 72523 318859 72526
rect 332593 72450 332659 72453
rect 219390 72448 332659 72450
rect 219390 72392 332598 72448
rect 332654 72392 332659 72448
rect 219390 72390 332659 72392
rect 169109 72387 169175 72390
rect 192477 72387 192543 72390
rect 332593 72387 332659 72390
rect 112805 71770 112871 71773
rect 147070 71770 147076 71772
rect 112805 71768 147076 71770
rect -960 71634 480 71724
rect 112805 71712 112810 71768
rect 112866 71712 147076 71768
rect 112805 71710 147076 71712
rect 112805 71707 112871 71710
rect 147070 71708 147076 71710
rect 147140 71708 147146 71772
rect 170673 71770 170739 71773
rect 214741 71770 214807 71773
rect 170673 71768 214807 71770
rect 170673 71712 170678 71768
rect 170734 71712 214746 71768
rect 214802 71712 214807 71768
rect 170673 71710 214807 71712
rect 170673 71707 170739 71710
rect 214741 71707 214807 71710
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 98453 71634 98519 71637
rect 132861 71634 132927 71637
rect 98453 71632 132927 71634
rect 98453 71576 98458 71632
rect 98514 71576 132866 71632
rect 132922 71576 132927 71632
rect 98453 71574 132927 71576
rect 98453 71571 98519 71574
rect 132861 71571 132927 71574
rect 173433 71634 173499 71637
rect 207238 71634 207244 71636
rect 173433 71632 207244 71634
rect 173433 71576 173438 71632
rect 173494 71576 207244 71632
rect 173433 71574 207244 71576
rect 173433 71571 173499 71574
rect 207238 71572 207244 71574
rect 207308 71634 207314 71636
rect 207308 71574 214666 71634
rect 207308 71572 207314 71574
rect 116853 71498 116919 71501
rect 149278 71498 149284 71500
rect 116853 71496 149284 71498
rect 116853 71440 116858 71496
rect 116914 71440 149284 71496
rect 116853 71438 149284 71440
rect 116853 71435 116919 71438
rect 149278 71436 149284 71438
rect 149348 71498 149354 71500
rect 149646 71498 149652 71500
rect 149348 71438 149652 71498
rect 149348 71436 149354 71438
rect 149646 71436 149652 71438
rect 149716 71436 149722 71500
rect 177757 71498 177823 71501
rect 211429 71498 211495 71501
rect 177757 71496 211495 71498
rect 177757 71440 177762 71496
rect 177818 71440 211434 71496
rect 211490 71440 211495 71496
rect 177757 71438 211495 71440
rect 177757 71435 177823 71438
rect 211429 71435 211495 71438
rect 122414 71300 122420 71364
rect 122484 71362 122490 71364
rect 152406 71362 152412 71364
rect 122484 71302 152412 71362
rect 122484 71300 122490 71302
rect 152406 71300 152412 71302
rect 152476 71300 152482 71364
rect 174997 71362 175063 71365
rect 174997 71360 200130 71362
rect 174997 71304 175002 71360
rect 175058 71304 200130 71360
rect 174997 71302 200130 71304
rect 174997 71299 175063 71302
rect 9673 71226 9739 71229
rect 98453 71226 98519 71229
rect 9673 71224 98519 71226
rect 9673 71168 9678 71224
rect 9734 71168 98458 71224
rect 98514 71168 98519 71224
rect 9673 71166 98519 71168
rect 9673 71163 9739 71166
rect 98453 71163 98519 71166
rect 120901 71226 120967 71229
rect 148174 71226 148180 71228
rect 120901 71224 148180 71226
rect 120901 71168 120906 71224
rect 120962 71168 148180 71224
rect 120901 71166 148180 71168
rect 120901 71163 120967 71166
rect 148174 71164 148180 71166
rect 148244 71164 148250 71228
rect 9029 71090 9095 71093
rect 104893 71090 104959 71093
rect 106038 71090 106044 71092
rect 9029 71088 106044 71090
rect 9029 71032 9034 71088
rect 9090 71032 104898 71088
rect 104954 71032 106044 71088
rect 9029 71030 106044 71032
rect 9029 71027 9095 71030
rect 104893 71027 104959 71030
rect 106038 71028 106044 71030
rect 106108 71028 106114 71092
rect 146477 71090 146543 71093
rect 178033 71090 178099 71093
rect 146477 71088 178099 71090
rect 146477 71032 146482 71088
rect 146538 71032 178038 71088
rect 178094 71032 178099 71088
rect 146477 71030 178099 71032
rect 200070 71090 200130 71302
rect 214606 71226 214666 71574
rect 214741 71362 214807 71365
rect 494053 71362 494119 71365
rect 214741 71360 494119 71362
rect 214741 71304 214746 71360
rect 214802 71304 494058 71360
rect 494114 71304 494119 71360
rect 214741 71302 494119 71304
rect 214741 71299 214807 71302
rect 494053 71299 494119 71302
rect 531313 71226 531379 71229
rect 214606 71224 531379 71226
rect 214606 71168 531318 71224
rect 531374 71168 531379 71224
rect 214606 71166 531379 71168
rect 531313 71163 531379 71166
rect 201718 71090 201724 71092
rect 200070 71030 201724 71090
rect 146477 71027 146543 71030
rect 178033 71027 178099 71030
rect 201718 71028 201724 71030
rect 201788 71090 201794 71092
rect 547873 71090 547939 71093
rect 201788 71088 547939 71090
rect 201788 71032 547878 71088
rect 547934 71032 547939 71088
rect 201788 71030 547939 71032
rect 201788 71028 201794 71030
rect 547873 71027 547939 71030
rect 97257 70274 97323 70277
rect 144310 70274 144316 70276
rect 97257 70272 144316 70274
rect 97257 70216 97262 70272
rect 97318 70216 144316 70272
rect 97257 70214 144316 70216
rect 97257 70211 97323 70214
rect 144310 70212 144316 70214
rect 144380 70212 144386 70276
rect 171726 70212 171732 70276
rect 171796 70274 171802 70276
rect 171796 70214 209790 70274
rect 171796 70212 171802 70214
rect 113582 70076 113588 70140
rect 113652 70138 113658 70140
rect 154113 70138 154179 70141
rect 113652 70136 154179 70138
rect 113652 70080 154118 70136
rect 154174 70080 154179 70136
rect 113652 70078 154179 70080
rect 113652 70076 113658 70078
rect 154113 70075 154179 70078
rect 175549 70138 175615 70141
rect 205214 70138 205220 70140
rect 175549 70136 205220 70138
rect 175549 70080 175554 70136
rect 175610 70080 205220 70136
rect 175549 70078 205220 70080
rect 175549 70075 175615 70078
rect 205214 70076 205220 70078
rect 205284 70076 205290 70140
rect 118550 69940 118556 70004
rect 118620 70002 118626 70004
rect 154205 70002 154271 70005
rect 118620 70000 154271 70002
rect 118620 69944 154210 70000
rect 154266 69944 154271 70000
rect 118620 69942 154271 69944
rect 118620 69940 118626 69942
rect 154205 69939 154271 69942
rect 164693 70002 164759 70005
rect 191598 70002 191604 70004
rect 164693 70000 191604 70002
rect 164693 69944 164698 70000
rect 164754 69944 191604 70000
rect 164693 69942 191604 69944
rect 164693 69939 164759 69942
rect 191598 69940 191604 69942
rect 191668 69940 191674 70004
rect 102777 69868 102843 69869
rect 102726 69866 102732 69868
rect 102686 69806 102732 69866
rect 102796 69864 102843 69868
rect 102838 69808 102843 69864
rect 102726 69804 102732 69806
rect 102796 69804 102843 69808
rect 121310 69804 121316 69868
rect 121380 69866 121386 69868
rect 121380 69806 142170 69866
rect 121380 69804 121386 69806
rect 102777 69803 102843 69804
rect 142110 69730 142170 69806
rect 150617 69730 150683 69733
rect 142110 69728 150683 69730
rect 142110 69672 150622 69728
rect 150678 69672 150683 69728
rect 142110 69670 150683 69672
rect 209730 69730 209790 70214
rect 214465 69730 214531 69733
rect 502977 69730 503043 69733
rect 209730 69728 503043 69730
rect 209730 69672 214470 69728
rect 214526 69672 502982 69728
rect 503038 69672 503043 69728
rect 209730 69670 503043 69672
rect 150617 69667 150683 69670
rect 214465 69667 214531 69670
rect 502977 69667 503043 69670
rect 18597 69594 18663 69597
rect 102777 69594 102843 69597
rect 18597 69592 102843 69594
rect 18597 69536 18602 69592
rect 18658 69536 102782 69592
rect 102838 69536 102843 69592
rect 18597 69534 102843 69536
rect 18597 69531 18663 69534
rect 102777 69531 102843 69534
rect 205214 69532 205220 69596
rect 205284 69594 205290 69596
rect 557533 69594 557599 69597
rect 205284 69592 557599 69594
rect 205284 69536 557538 69592
rect 557594 69536 557599 69592
rect 205284 69534 557599 69536
rect 205284 69532 205290 69534
rect 557533 69531 557599 69534
rect 150617 69050 150683 69053
rect 151445 69050 151511 69053
rect 150617 69048 151511 69050
rect 150617 68992 150622 69048
rect 150678 68992 151450 69048
rect 151506 68992 151511 69048
rect 150617 68990 151511 68992
rect 150617 68987 150683 68990
rect 151445 68987 151511 68990
rect 154205 69050 154271 69053
rect 154389 69050 154455 69053
rect 154205 69048 154455 69050
rect 154205 68992 154210 69048
rect 154266 68992 154394 69048
rect 154450 68992 154455 69048
rect 154205 68990 154455 68992
rect 154205 68987 154271 68990
rect 154389 68987 154455 68990
rect 102910 68852 102916 68916
rect 102980 68914 102986 68916
rect 103145 68914 103211 68917
rect 102980 68912 103211 68914
rect 102980 68856 103150 68912
rect 103206 68856 103211 68912
rect 102980 68854 103211 68856
rect 102980 68852 102986 68854
rect 103145 68851 103211 68854
rect 114134 68852 114140 68916
rect 114204 68914 114210 68916
rect 147990 68914 147996 68916
rect 114204 68854 147996 68914
rect 114204 68852 114210 68854
rect 147990 68852 147996 68854
rect 148060 68914 148066 68916
rect 148542 68914 148548 68916
rect 148060 68854 148548 68914
rect 148060 68852 148066 68854
rect 148542 68852 148548 68854
rect 148612 68852 148618 68916
rect 177113 68914 177179 68917
rect 177113 68912 200130 68914
rect 177113 68856 177118 68912
rect 177174 68856 200130 68912
rect 177113 68854 200130 68856
rect 177113 68851 177179 68854
rect 112846 68716 112852 68780
rect 112916 68778 112922 68780
rect 146518 68778 146524 68780
rect 112916 68718 146524 68778
rect 112916 68716 112922 68718
rect 146518 68716 146524 68718
rect 146588 68716 146594 68780
rect 118325 68642 118391 68645
rect 149094 68642 149100 68644
rect 118325 68640 149100 68642
rect 118325 68584 118330 68640
rect 118386 68584 149100 68640
rect 118325 68582 149100 68584
rect 118325 68579 118391 68582
rect 149094 68580 149100 68582
rect 149164 68642 149170 68644
rect 150014 68642 150020 68644
rect 149164 68582 150020 68642
rect 149164 68580 149170 68582
rect 150014 68580 150020 68582
rect 150084 68580 150090 68644
rect 122046 68444 122052 68508
rect 122116 68506 122122 68508
rect 147806 68506 147812 68508
rect 122116 68446 147812 68506
rect 122116 68444 122122 68446
rect 147806 68444 147812 68446
rect 147876 68506 147882 68508
rect 148174 68506 148180 68508
rect 147876 68446 148180 68506
rect 147876 68444 147882 68446
rect 148174 68444 148180 68446
rect 148244 68444 148250 68508
rect 26233 68234 26299 68237
rect 103145 68234 103211 68237
rect 26233 68232 103211 68234
rect 26233 68176 26238 68232
rect 26294 68176 103150 68232
rect 103206 68176 103211 68232
rect 26233 68174 103211 68176
rect 200070 68234 200130 68854
rect 203190 68234 203196 68236
rect 200070 68174 203196 68234
rect 26233 68171 26299 68174
rect 103145 68171 103211 68174
rect 203190 68172 203196 68174
rect 203260 68234 203266 68236
rect 574737 68234 574803 68237
rect 203260 68232 574803 68234
rect 203260 68176 574742 68232
rect 574798 68176 574803 68232
rect 203260 68174 574803 68176
rect 203260 68172 203266 68174
rect 574737 68171 574803 68174
rect 119654 67492 119660 67556
rect 119724 67554 119730 67556
rect 153561 67554 153627 67557
rect 119724 67552 153627 67554
rect 119724 67496 153566 67552
rect 153622 67496 153627 67552
rect 119724 67494 153627 67496
rect 119724 67492 119730 67494
rect 153561 67491 153627 67494
rect 161473 67554 161539 67557
rect 162485 67554 162551 67557
rect 189206 67554 189212 67556
rect 161473 67552 189212 67554
rect 161473 67496 161478 67552
rect 161534 67496 162490 67552
rect 162546 67496 189212 67552
rect 161473 67494 189212 67496
rect 161473 67491 161539 67494
rect 162485 67491 162551 67494
rect 189206 67492 189212 67494
rect 189276 67492 189282 67556
rect 204897 67554 204963 67557
rect 205030 67554 205036 67556
rect 204897 67552 205036 67554
rect 204897 67496 204902 67552
rect 204958 67496 205036 67552
rect 204897 67494 205036 67496
rect 204897 67491 204963 67494
rect 205030 67492 205036 67494
rect 205100 67492 205106 67556
rect 133454 67418 133460 67420
rect 108990 67358 133460 67418
rect 7649 66874 7715 66877
rect 99230 66874 99236 66876
rect 7649 66872 99236 66874
rect 7649 66816 7654 66872
rect 7710 66816 99236 66872
rect 7649 66814 99236 66816
rect 7649 66811 7715 66814
rect 99230 66812 99236 66814
rect 99300 66874 99306 66876
rect 108990 66874 109050 67358
rect 133454 67356 133460 67358
rect 133524 67356 133530 67420
rect 168741 67418 168807 67421
rect 169661 67418 169727 67421
rect 187734 67418 187740 67420
rect 168741 67416 187740 67418
rect 168741 67360 168746 67416
rect 168802 67360 169666 67416
rect 169722 67360 187740 67416
rect 168741 67358 187740 67360
rect 168741 67355 168807 67358
rect 169661 67355 169727 67358
rect 187734 67356 187740 67358
rect 187804 67356 187810 67420
rect 99300 66814 109050 66874
rect 99300 66812 99306 66814
rect 149462 66812 149468 66876
rect 149532 66874 149538 66876
rect 227713 66874 227779 66877
rect 149532 66872 227779 66874
rect 149532 66816 227718 66872
rect 227774 66816 227779 66872
rect 149532 66814 227779 66816
rect 149532 66812 149538 66814
rect 227713 66811 227779 66814
rect 153561 66330 153627 66333
rect 153929 66330 153995 66333
rect 153561 66328 153995 66330
rect 153561 66272 153566 66328
rect 153622 66272 153934 66328
rect 153990 66272 153995 66328
rect 153561 66270 153995 66272
rect 153561 66267 153627 66270
rect 153929 66267 153995 66270
rect 104433 66196 104499 66197
rect 104382 66194 104388 66196
rect 104342 66134 104388 66194
rect 104452 66192 104499 66196
rect 104494 66136 104499 66192
rect 104382 66132 104388 66134
rect 104452 66132 104499 66136
rect 104433 66131 104499 66132
rect 110137 66194 110203 66197
rect 143942 66194 143948 66196
rect 110137 66192 143948 66194
rect 110137 66136 110142 66192
rect 110198 66136 143948 66192
rect 110137 66134 143948 66136
rect 110137 66131 110203 66134
rect 143942 66132 143948 66134
rect 144012 66194 144018 66196
rect 144678 66194 144684 66196
rect 144012 66134 144684 66194
rect 144012 66132 144018 66134
rect 144678 66132 144684 66134
rect 144748 66132 144754 66196
rect 155534 66132 155540 66196
rect 155604 66194 155610 66196
rect 215661 66194 215727 66197
rect 155604 66192 219450 66194
rect 155604 66136 215666 66192
rect 215722 66136 219450 66192
rect 155604 66134 219450 66136
rect 155604 66132 155610 66134
rect 215661 66131 215727 66134
rect 122598 65996 122604 66060
rect 122668 66058 122674 66060
rect 156597 66058 156663 66061
rect 122668 66056 156663 66058
rect 122668 66000 156602 66056
rect 156658 66000 156663 66056
rect 122668 65998 156663 66000
rect 122668 65996 122674 65998
rect 156597 65995 156663 65998
rect 170438 65996 170444 66060
rect 170508 66058 170514 66060
rect 214005 66058 214071 66061
rect 170508 66056 214482 66058
rect 170508 66000 214010 66056
rect 214066 66000 214482 66056
rect 170508 65998 214482 66000
rect 170508 65996 170514 65998
rect 214005 65995 214071 65998
rect 110689 65922 110755 65925
rect 143758 65922 143764 65924
rect 110689 65920 143764 65922
rect 110689 65864 110694 65920
rect 110750 65864 143764 65920
rect 110689 65862 143764 65864
rect 110689 65859 110755 65862
rect 143758 65860 143764 65862
rect 143828 65860 143834 65924
rect 171910 65860 171916 65924
rect 171980 65922 171986 65924
rect 171980 65862 200130 65922
rect 171980 65860 171986 65862
rect 59353 65650 59419 65653
rect 104433 65650 104499 65653
rect 59353 65648 104499 65650
rect 59353 65592 59358 65648
rect 59414 65592 104438 65648
rect 104494 65592 104499 65648
rect 59353 65590 104499 65592
rect 59353 65587 59419 65590
rect 104433 65587 104499 65590
rect 57973 65514 58039 65517
rect 108246 65514 108252 65516
rect 57973 65512 108252 65514
rect 57973 65456 57978 65512
rect 58034 65456 108252 65512
rect 57973 65454 108252 65456
rect 57973 65451 58039 65454
rect 108246 65452 108252 65454
rect 108316 65452 108322 65516
rect 117221 65514 117287 65517
rect 140998 65514 141004 65516
rect 117221 65512 141004 65514
rect 117221 65456 117226 65512
rect 117282 65456 141004 65512
rect 117221 65454 141004 65456
rect 117221 65451 117287 65454
rect 140998 65452 141004 65454
rect 141068 65452 141074 65516
rect 147254 65452 147260 65516
rect 147324 65514 147330 65516
rect 188337 65514 188403 65517
rect 147324 65512 188403 65514
rect 147324 65456 188342 65512
rect 188398 65456 188403 65512
rect 147324 65454 188403 65456
rect 200070 65514 200130 65862
rect 214422 65650 214482 65998
rect 219390 65786 219450 66134
rect 295333 65786 295399 65789
rect 219390 65784 295399 65786
rect 219390 65728 295338 65784
rect 295394 65728 295399 65784
rect 219390 65726 295399 65728
rect 295333 65723 295399 65726
rect 498193 65650 498259 65653
rect 214422 65648 498259 65650
rect 214422 65592 498198 65648
rect 498254 65592 498259 65648
rect 214422 65590 498259 65592
rect 498193 65587 498259 65590
rect 214281 65514 214347 65517
rect 507853 65514 507919 65517
rect 200070 65512 507919 65514
rect 200070 65456 214286 65512
rect 214342 65456 507858 65512
rect 507914 65456 507919 65512
rect 200070 65454 507919 65456
rect 147324 65452 147330 65454
rect 188337 65451 188403 65454
rect 214281 65451 214347 65454
rect 507853 65451 507919 65454
rect 97901 64834 97967 64837
rect 143574 64834 143580 64836
rect 97901 64832 143580 64834
rect 97901 64776 97906 64832
rect 97962 64776 143580 64832
rect 97901 64774 143580 64776
rect 97901 64771 97967 64774
rect 143574 64772 143580 64774
rect 143644 64772 143650 64836
rect 153193 64834 153259 64837
rect 154297 64834 154363 64837
rect 147630 64832 154363 64834
rect 147630 64776 153198 64832
rect 153254 64776 154302 64832
rect 154358 64776 154363 64832
rect 147630 64774 154363 64776
rect 116342 64636 116348 64700
rect 116412 64698 116418 64700
rect 147630 64698 147690 64774
rect 153193 64771 153259 64774
rect 154297 64771 154363 64774
rect 172094 64772 172100 64836
rect 172164 64834 172170 64836
rect 200614 64834 200620 64836
rect 172164 64774 200620 64834
rect 172164 64772 172170 64774
rect 116412 64638 147690 64698
rect 116412 64636 116418 64638
rect 121126 64500 121132 64564
rect 121196 64562 121202 64564
rect 154849 64562 154915 64565
rect 121196 64560 154915 64562
rect 121196 64504 154854 64560
rect 154910 64504 154915 64560
rect 121196 64502 154915 64504
rect 121196 64500 121202 64502
rect 154849 64499 154915 64502
rect 57237 64290 57303 64293
rect 103789 64290 103855 64293
rect 104198 64290 104204 64292
rect 57237 64288 104204 64290
rect 57237 64232 57242 64288
rect 57298 64232 103794 64288
rect 103850 64232 104204 64288
rect 57237 64230 104204 64232
rect 57237 64227 57303 64230
rect 103789 64227 103855 64230
rect 104198 64228 104204 64230
rect 104268 64228 104274 64292
rect 4797 64154 4863 64157
rect 103973 64156 104039 64157
rect 103973 64154 104020 64156
rect 4797 64152 104020 64154
rect 104084 64154 104090 64156
rect 200070 64154 200130 64774
rect 200614 64772 200620 64774
rect 200684 64772 200690 64836
rect 511993 64154 512059 64157
rect 4797 64096 4802 64152
rect 4858 64096 103978 64152
rect 4797 64094 104020 64096
rect 4797 64091 4863 64094
rect 103973 64092 104020 64094
rect 104084 64094 104166 64154
rect 200070 64152 512059 64154
rect 200070 64096 511998 64152
rect 512054 64096 512059 64152
rect 200070 64094 512059 64096
rect 104084 64092 104090 64094
rect 103973 64091 104039 64092
rect 511993 64091 512059 64094
rect 143574 63548 143580 63612
rect 143644 63610 143650 63612
rect 144494 63610 144500 63612
rect 143644 63550 144500 63610
rect 143644 63548 143650 63550
rect 144494 63548 144500 63550
rect 144564 63548 144570 63612
rect 151486 63412 151492 63476
rect 151556 63474 151562 63476
rect 217593 63474 217659 63477
rect 151556 63472 219450 63474
rect 151556 63416 217598 63472
rect 217654 63416 219450 63472
rect 151556 63414 219450 63416
rect 151556 63412 151562 63414
rect 217593 63411 217659 63414
rect 175958 63276 175964 63340
rect 176028 63338 176034 63340
rect 217317 63338 217383 63341
rect 176028 63336 217383 63338
rect 176028 63280 217322 63336
rect 217378 63280 217383 63336
rect 176028 63278 217383 63280
rect 176028 63276 176034 63278
rect 217317 63275 217383 63278
rect 166206 63140 166212 63204
rect 166276 63202 166282 63204
rect 219390 63202 219450 63414
rect 245653 63202 245719 63205
rect 166276 63142 200130 63202
rect 219390 63200 245719 63202
rect 219390 63144 245658 63200
rect 245714 63144 245719 63200
rect 219390 63142 245719 63144
rect 166276 63140 166282 63142
rect 200070 63066 200130 63142
rect 245653 63139 245719 63142
rect 200389 63066 200455 63069
rect 430573 63066 430639 63069
rect 200070 63064 430639 63066
rect 200070 63008 200394 63064
rect 200450 63008 430578 63064
rect 430634 63008 430639 63064
rect 200070 63006 430639 63008
rect 200389 63003 200455 63006
rect 430573 63003 430639 63006
rect 172278 62868 172284 62932
rect 172348 62930 172354 62932
rect 201534 62930 201540 62932
rect 172348 62870 201540 62930
rect 172348 62868 172354 62870
rect 201534 62868 201540 62870
rect 201604 62930 201610 62932
rect 514017 62930 514083 62933
rect 201604 62928 514083 62930
rect 201604 62872 514022 62928
rect 514078 62872 514083 62928
rect 201604 62870 514083 62872
rect 201604 62868 201610 62870
rect 514017 62867 514083 62870
rect 148726 62732 148732 62796
rect 148796 62794 148802 62796
rect 214005 62794 214071 62797
rect 148796 62792 214071 62794
rect 148796 62736 214010 62792
rect 214066 62736 214071 62792
rect 148796 62734 214071 62736
rect 148796 62732 148802 62734
rect 214005 62731 214071 62734
rect 217317 62794 217383 62797
rect 561673 62794 561739 62797
rect 217317 62792 561739 62794
rect 217317 62736 217322 62792
rect 217378 62736 561678 62792
rect 561734 62736 561739 62792
rect 217317 62734 561739 62736
rect 217317 62731 217383 62734
rect 561673 62731 561739 62734
rect 100293 62114 100359 62117
rect 134190 62114 134196 62116
rect 100293 62112 134196 62114
rect 100293 62056 100298 62112
rect 100354 62056 134196 62112
rect 100293 62054 134196 62056
rect 100293 62051 100359 62054
rect 134190 62052 134196 62054
rect 134260 62052 134266 62116
rect 164918 62052 164924 62116
rect 164988 62114 164994 62116
rect 199101 62114 199167 62117
rect 199837 62114 199903 62117
rect 164988 62112 199903 62114
rect 164988 62056 199106 62112
rect 199162 62056 199842 62112
rect 199898 62056 199903 62112
rect 164988 62054 199903 62056
rect 164988 62052 164994 62054
rect 199101 62051 199167 62054
rect 199837 62051 199903 62054
rect 138606 61978 138612 61980
rect 108990 61918 138612 61978
rect 75177 61570 75243 61573
rect 105997 61570 106063 61573
rect 108990 61570 109050 61918
rect 138606 61916 138612 61918
rect 138676 61916 138682 61980
rect 176142 61916 176148 61980
rect 176212 61978 176218 61980
rect 203006 61978 203012 61980
rect 176212 61918 203012 61978
rect 176212 61916 176218 61918
rect 203006 61916 203012 61918
rect 203076 61978 203082 61980
rect 204110 61978 204116 61980
rect 203076 61918 204116 61978
rect 203076 61916 203082 61918
rect 204110 61916 204116 61918
rect 204180 61916 204186 61980
rect 116945 61842 117011 61845
rect 140814 61842 140820 61844
rect 116945 61840 140820 61842
rect 116945 61784 116950 61840
rect 117006 61784 140820 61840
rect 116945 61782 140820 61784
rect 116945 61779 117011 61782
rect 140814 61780 140820 61782
rect 140884 61780 140890 61844
rect 150014 61644 150020 61708
rect 150084 61706 150090 61708
rect 230473 61706 230539 61709
rect 150084 61704 230539 61706
rect 150084 61648 230478 61704
rect 230534 61648 230539 61704
rect 150084 61646 230539 61648
rect 150084 61644 150090 61646
rect 230473 61643 230539 61646
rect 75177 61568 109050 61570
rect 75177 61512 75182 61568
rect 75238 61512 106002 61568
rect 106058 61512 109050 61568
rect 75177 61510 109050 61512
rect 199837 61570 199903 61573
rect 422937 61570 423003 61573
rect 199837 61568 423003 61570
rect 199837 61512 199842 61568
rect 199898 61512 422942 61568
rect 422998 61512 423003 61568
rect 199837 61510 423003 61512
rect 75177 61507 75243 61510
rect 105997 61507 106063 61510
rect 199837 61507 199903 61510
rect 422937 61507 423003 61510
rect 23473 61434 23539 61437
rect 100293 61434 100359 61437
rect 23473 61432 100359 61434
rect 23473 61376 23478 61432
rect 23534 61376 100298 61432
rect 100354 61376 100359 61432
rect 23473 61374 100359 61376
rect 23473 61371 23539 61374
rect 100293 61371 100359 61374
rect 204110 61372 204116 61436
rect 204180 61434 204186 61436
rect 563697 61434 563763 61437
rect 204180 61432 563763 61434
rect 204180 61376 563702 61432
rect 563758 61376 563763 61432
rect 204180 61374 563763 61376
rect 204180 61372 204186 61374
rect 563697 61371 563763 61374
rect 193673 60620 193739 60621
rect 193622 60618 193628 60620
rect 193582 60558 193628 60618
rect 193692 60616 193739 60620
rect 193734 60560 193739 60616
rect 193622 60556 193628 60558
rect 193692 60556 193739 60560
rect 193673 60555 193739 60556
rect 173566 60420 173572 60484
rect 173636 60482 173642 60484
rect 212625 60482 212691 60485
rect 213821 60482 213887 60485
rect 173636 60480 213887 60482
rect 173636 60424 212630 60480
rect 212686 60424 213826 60480
rect 213882 60424 213887 60480
rect 173636 60422 213887 60424
rect 173636 60420 173642 60422
rect 212625 60419 212691 60422
rect 213821 60419 213887 60422
rect 165102 60284 165108 60348
rect 165172 60346 165178 60348
rect 219525 60346 219591 60349
rect 165172 60344 219591 60346
rect 165172 60288 219530 60344
rect 219586 60288 219591 60344
rect 165172 60286 219591 60288
rect 165172 60284 165178 60286
rect 219390 60074 219450 60286
rect 219525 60283 219591 60286
rect 412633 60074 412699 60077
rect 219390 60072 412699 60074
rect 219390 60016 412638 60072
rect 412694 60016 412699 60072
rect 219390 60014 412699 60016
rect 412633 60011 412699 60014
rect 213821 59938 213887 59941
rect 527817 59938 527883 59941
rect 213821 59936 527883 59938
rect 213821 59880 213826 59936
rect 213882 59880 527822 59936
rect 527878 59880 527883 59936
rect 213821 59878 527883 59880
rect 213821 59875 213887 59878
rect 527817 59875 527883 59878
rect 580625 59666 580691 59669
rect 583520 59666 584960 59756
rect 580625 59664 584960 59666
rect 580625 59608 580630 59664
rect 580686 59608 584960 59664
rect 580625 59606 584960 59608
rect 580625 59603 580691 59606
rect 583520 59516 584960 59606
rect 139894 59258 139900 59260
rect 113130 59198 139900 59258
rect -960 58578 480 58668
rect 93853 58578 93919 58581
rect 108798 58578 108804 58580
rect -960 58518 674 58578
rect -960 58442 480 58518
rect 614 58442 674 58518
rect 93853 58576 108804 58578
rect 93853 58520 93858 58576
rect 93914 58520 108804 58576
rect 93853 58518 108804 58520
rect 93853 58515 93919 58518
rect 108798 58516 108804 58518
rect 108868 58578 108874 58580
rect 113130 58578 113190 59198
rect 139894 59196 139900 59198
rect 139964 59196 139970 59260
rect 151670 59196 151676 59260
rect 151740 59258 151746 59260
rect 217041 59258 217107 59261
rect 151740 59256 229110 59258
rect 151740 59200 217046 59256
rect 217102 59200 229110 59256
rect 151740 59198 229110 59200
rect 151740 59196 151746 59198
rect 217041 59195 217107 59198
rect 154062 59060 154068 59124
rect 154132 59122 154138 59124
rect 215385 59122 215451 59125
rect 154132 59120 219450 59122
rect 154132 59064 215390 59120
rect 215446 59064 219450 59120
rect 154132 59062 219450 59064
rect 154132 59060 154138 59062
rect 215385 59059 215451 59062
rect 170622 58924 170628 58988
rect 170692 58986 170698 58988
rect 170692 58926 209790 58986
rect 170692 58924 170698 58926
rect 174486 58788 174492 58852
rect 174556 58850 174562 58852
rect 174556 58790 200130 58850
rect 174556 58788 174562 58790
rect 108868 58518 113190 58578
rect 200070 58578 200130 58790
rect 209730 58714 209790 58926
rect 219390 58850 219450 59062
rect 229050 58986 229110 59198
rect 249793 58986 249859 58989
rect 229050 58984 249859 58986
rect 229050 58928 249798 58984
rect 249854 58928 249859 58984
rect 229050 58926 249859 58928
rect 249793 58923 249859 58926
rect 281533 58850 281599 58853
rect 219390 58848 281599 58850
rect 219390 58792 281538 58848
rect 281594 58792 281599 58848
rect 219390 58790 281599 58792
rect 281533 58787 281599 58790
rect 214189 58714 214255 58717
rect 489177 58714 489243 58717
rect 209730 58712 489243 58714
rect 209730 58656 214194 58712
rect 214250 58656 489182 58712
rect 489238 58656 489243 58712
rect 209730 58654 489243 58656
rect 214189 58651 214255 58654
rect 489177 58651 489243 58654
rect 208577 58578 208643 58581
rect 538857 58578 538923 58581
rect 200070 58576 538923 58578
rect 200070 58520 208582 58576
rect 208638 58520 538862 58576
rect 538918 58520 538923 58576
rect 200070 58518 538923 58520
rect 108868 58516 108874 58518
rect 208577 58515 208643 58518
rect 538857 58515 538923 58518
rect -960 58428 674 58442
rect 246 58382 674 58428
rect 246 58034 306 58382
rect 111006 58034 111012 58036
rect 246 57974 111012 58034
rect 111006 57972 111012 57974
rect 111076 57972 111082 58036
rect 106181 57898 106247 57901
rect 138422 57898 138428 57900
rect 84150 57896 138428 57898
rect 84150 57840 106186 57896
rect 106242 57840 138428 57896
rect 84150 57838 138428 57840
rect 80053 57354 80119 57357
rect 84150 57354 84210 57838
rect 106181 57835 106247 57838
rect 138422 57836 138428 57838
rect 138492 57836 138498 57900
rect 174670 57836 174676 57900
rect 174740 57898 174746 57900
rect 217225 57898 217291 57901
rect 174740 57896 217291 57898
rect 174740 57840 217230 57896
rect 217286 57840 217291 57896
rect 174740 57838 217291 57840
rect 174740 57836 174746 57838
rect 217225 57835 217291 57838
rect 134006 57762 134012 57764
rect 80053 57352 84210 57354
rect 80053 57296 80058 57352
rect 80114 57296 84210 57352
rect 80053 57294 84210 57296
rect 103470 57702 134012 57762
rect 80053 57291 80119 57294
rect 25497 57218 25563 57221
rect 101990 57218 101996 57220
rect 25497 57216 101996 57218
rect 25497 57160 25502 57216
rect 25558 57160 101996 57216
rect 25497 57158 101996 57160
rect 25497 57155 25563 57158
rect 101990 57156 101996 57158
rect 102060 57218 102066 57220
rect 103470 57218 103530 57702
rect 134006 57700 134012 57702
rect 134076 57700 134082 57764
rect 166390 57700 166396 57764
rect 166460 57762 166466 57764
rect 200297 57762 200363 57765
rect 166460 57760 200363 57762
rect 166460 57704 200302 57760
rect 200358 57704 200363 57760
rect 166460 57702 200363 57704
rect 166460 57700 166466 57702
rect 200070 57354 200130 57702
rect 200297 57699 200363 57702
rect 432597 57354 432663 57357
rect 200070 57352 432663 57354
rect 200070 57296 432602 57352
rect 432658 57296 432663 57352
rect 200070 57294 432663 57296
rect 432597 57291 432663 57294
rect 102060 57158 103530 57218
rect 217225 57218 217291 57221
rect 545757 57218 545823 57221
rect 217225 57216 545823 57218
rect 217225 57160 217230 57216
rect 217286 57160 545762 57216
rect 545818 57160 545823 57216
rect 217225 57158 545823 57160
rect 102060 57156 102066 57158
rect 217225 57155 217291 57158
rect 545757 57155 545823 57158
rect 99414 56476 99420 56540
rect 99484 56538 99490 56540
rect 100334 56538 100340 56540
rect 99484 56478 100340 56538
rect 99484 56476 99490 56478
rect 100334 56476 100340 56478
rect 100404 56538 100410 56540
rect 133270 56538 133276 56540
rect 100404 56478 133276 56538
rect 100404 56476 100410 56478
rect 133270 56476 133276 56478
rect 133340 56476 133346 56540
rect 144678 56476 144684 56540
rect 144748 56538 144754 56540
rect 149789 56538 149855 56541
rect 144748 56536 149855 56538
rect 144748 56480 149794 56536
rect 149850 56480 149855 56536
rect 144748 56478 149855 56480
rect 144748 56476 144754 56478
rect 149789 56475 149855 56478
rect 104750 56402 104756 56404
rect 103470 56342 104756 56402
rect 56593 55994 56659 55997
rect 103470 55994 103530 56342
rect 104750 56340 104756 56342
rect 104820 56402 104826 56404
rect 137502 56402 137508 56404
rect 104820 56342 137508 56402
rect 104820 56340 104826 56342
rect 137502 56340 137508 56342
rect 137572 56340 137578 56404
rect 56593 55992 103530 55994
rect 56593 55936 56598 55992
rect 56654 55936 103530 55992
rect 56593 55934 103530 55936
rect 56593 55931 56659 55934
rect 12433 55858 12499 55861
rect 99414 55858 99420 55860
rect 12433 55856 99420 55858
rect 12433 55800 12438 55856
rect 12494 55800 99420 55856
rect 12433 55798 99420 55800
rect 12433 55795 12499 55798
rect 99414 55796 99420 55798
rect 99484 55796 99490 55860
rect 101949 55178 102015 55181
rect 135846 55178 135852 55180
rect 101949 55176 135852 55178
rect 101949 55120 101954 55176
rect 102010 55120 135852 55176
rect 101949 55118 135852 55120
rect 101949 55115 102015 55118
rect 135846 55116 135852 55118
rect 135916 55116 135922 55180
rect 156822 55116 156828 55180
rect 156892 55178 156898 55180
rect 210049 55178 210115 55181
rect 156892 55176 219450 55178
rect 156892 55120 210054 55176
rect 210110 55120 219450 55176
rect 156892 55118 219450 55120
rect 156892 55116 156898 55118
rect 210049 55115 210115 55118
rect 170806 54980 170812 55044
rect 170876 55042 170882 55044
rect 211245 55042 211311 55045
rect 170876 55040 211311 55042
rect 170876 54984 211250 55040
rect 211306 54984 211311 55040
rect 170876 54982 211311 54984
rect 170876 54980 170882 54982
rect 211245 54979 211311 54982
rect 160870 54844 160876 54908
rect 160940 54906 160946 54908
rect 194593 54906 194659 54909
rect 160940 54904 194659 54906
rect 160940 54848 194598 54904
rect 194654 54848 194659 54904
rect 160940 54846 194659 54848
rect 160940 54844 160946 54846
rect 194593 54843 194659 54846
rect 219390 54770 219450 55118
rect 315297 54770 315363 54773
rect 219390 54768 315363 54770
rect 219390 54712 315302 54768
rect 315358 54712 315363 54768
rect 219390 54710 315363 54712
rect 315297 54707 315363 54710
rect 84193 54634 84259 54637
rect 109585 54636 109651 54637
rect 109534 54634 109540 54636
rect 84193 54632 109540 54634
rect 109604 54634 109651 54636
rect 194593 54634 194659 54637
rect 364977 54634 365043 54637
rect 109604 54632 109732 54634
rect 84193 54576 84198 54632
rect 84254 54576 109540 54632
rect 109646 54576 109732 54632
rect 84193 54574 109540 54576
rect 84193 54571 84259 54574
rect 109534 54572 109540 54574
rect 109604 54574 109732 54576
rect 194593 54632 365043 54634
rect 194593 54576 194598 54632
rect 194654 54576 364982 54632
rect 365038 54576 365043 54632
rect 194593 54574 365043 54576
rect 109604 54572 109651 54574
rect 109585 54571 109651 54572
rect 194593 54571 194659 54574
rect 364977 54571 365043 54574
rect 41413 54498 41479 54501
rect 101949 54498 102015 54501
rect 41413 54496 102015 54498
rect 41413 54440 41418 54496
rect 41474 54440 101954 54496
rect 102010 54440 102015 54496
rect 41413 54438 102015 54440
rect 41413 54435 41479 54438
rect 101949 54435 102015 54438
rect 148542 54436 148548 54500
rect 148612 54498 148618 54500
rect 210049 54498 210115 54501
rect 148612 54496 210115 54498
rect 148612 54440 210054 54496
rect 210110 54440 210115 54496
rect 148612 54438 210115 54440
rect 148612 54436 148618 54438
rect 210049 54435 210115 54438
rect 211245 54498 211311 54501
rect 486509 54498 486575 54501
rect 211245 54496 486575 54498
rect 211245 54440 211250 54496
rect 211306 54440 486514 54496
rect 486570 54440 486575 54496
rect 211245 54438 486575 54440
rect 211245 54435 211311 54438
rect 486509 54435 486575 54438
rect 92473 53818 92539 53821
rect 105445 53818 105511 53821
rect 139710 53818 139716 53820
rect 92473 53816 139716 53818
rect 92473 53760 92478 53816
rect 92534 53760 105450 53816
rect 105506 53760 139716 53816
rect 92473 53758 139716 53760
rect 92473 53755 92539 53758
rect 105445 53755 105511 53758
rect 139710 53756 139716 53758
rect 139780 53756 139786 53820
rect 154246 53756 154252 53820
rect 154316 53818 154322 53820
rect 215293 53818 215359 53821
rect 154316 53816 215359 53818
rect 154316 53760 215298 53816
rect 215354 53760 215359 53816
rect 154316 53758 215359 53760
rect 154316 53756 154322 53758
rect 215293 53755 215359 53758
rect 100518 53620 100524 53684
rect 100588 53682 100594 53684
rect 133086 53682 133092 53684
rect 100588 53622 133092 53682
rect 100588 53620 100594 53622
rect 133086 53620 133092 53622
rect 133156 53620 133162 53684
rect 162158 53620 162164 53684
rect 162228 53682 162234 53684
rect 196065 53682 196131 53685
rect 162228 53680 200130 53682
rect 162228 53624 196070 53680
rect 196126 53624 200130 53680
rect 162228 53622 200130 53624
rect 162228 53620 162234 53622
rect 196065 53619 196131 53622
rect 166574 53484 166580 53548
rect 166644 53546 166650 53548
rect 194542 53546 194548 53548
rect 166644 53486 194548 53546
rect 166644 53484 166650 53486
rect 194542 53484 194548 53486
rect 194612 53484 194618 53548
rect 200070 53274 200130 53622
rect 215293 53410 215359 53413
rect 284385 53410 284451 53413
rect 215293 53408 284451 53410
rect 215293 53352 215298 53408
rect 215354 53352 284390 53408
rect 284446 53352 284451 53408
rect 215293 53350 284451 53352
rect 215293 53347 215359 53350
rect 284385 53347 284451 53350
rect 382917 53274 382983 53277
rect 200070 53272 382983 53274
rect 200070 53216 382922 53272
rect 382978 53216 382983 53272
rect 200070 53214 382983 53216
rect 382917 53211 382983 53214
rect 17953 53138 18019 53141
rect 100518 53138 100524 53140
rect 17953 53136 100524 53138
rect 17953 53080 17958 53136
rect 18014 53080 100524 53136
rect 17953 53078 100524 53080
rect 17953 53075 18019 53078
rect 100518 53076 100524 53078
rect 100588 53076 100594 53140
rect 194542 53076 194548 53140
rect 194612 53138 194618 53140
rect 437473 53138 437539 53141
rect 194612 53136 437539 53138
rect 194612 53080 437478 53136
rect 437534 53080 437539 53136
rect 194612 53078 437539 53080
rect 194612 53076 194618 53078
rect 437473 53075 437539 53078
rect 107142 52396 107148 52460
rect 107212 52458 107218 52460
rect 138238 52458 138244 52460
rect 107212 52398 138244 52458
rect 107212 52396 107218 52398
rect 138238 52396 138244 52398
rect 138308 52396 138314 52460
rect 163262 52396 163268 52460
rect 163332 52458 163338 52460
rect 197445 52458 197511 52461
rect 163332 52456 197511 52458
rect 163332 52400 197450 52456
rect 197506 52400 197511 52456
rect 163332 52398 197511 52400
rect 163332 52396 163338 52398
rect 197445 52395 197511 52398
rect 167494 52260 167500 52324
rect 167564 52322 167570 52324
rect 201677 52322 201743 52325
rect 202781 52322 202847 52325
rect 167564 52320 202847 52322
rect 167564 52264 201682 52320
rect 201738 52264 202786 52320
rect 202842 52264 202847 52320
rect 167564 52262 202847 52264
rect 167564 52260 167570 52262
rect 201677 52259 201743 52262
rect 202781 52259 202847 52262
rect 161054 52124 161060 52188
rect 161124 52186 161130 52188
rect 193581 52186 193647 52189
rect 369853 52186 369919 52189
rect 161124 52184 369919 52186
rect 161124 52128 193586 52184
rect 193642 52128 369858 52184
rect 369914 52128 369919 52184
rect 161124 52126 369919 52128
rect 161124 52124 161130 52126
rect 193581 52123 193647 52126
rect 369853 52123 369919 52126
rect 189625 52050 189691 52053
rect 189758 52050 189764 52052
rect 189625 52048 189764 52050
rect 189625 51992 189630 52048
rect 189686 51992 189764 52048
rect 189625 51990 189764 51992
rect 189625 51987 189691 51990
rect 189758 51988 189764 51990
rect 189828 51988 189834 52052
rect 197445 52050 197511 52053
rect 400857 52050 400923 52053
rect 197445 52048 400923 52050
rect 197445 51992 197450 52048
rect 197506 51992 400862 52048
rect 400918 51992 400923 52048
rect 197445 51990 400923 51992
rect 197445 51987 197511 51990
rect 400857 51987 400923 51990
rect 202781 51914 202847 51917
rect 450537 51914 450603 51917
rect 202781 51912 450603 51914
rect 202781 51856 202786 51912
rect 202842 51856 450542 51912
rect 450598 51856 450603 51912
rect 202781 51854 450603 51856
rect 202781 51851 202847 51854
rect 450537 51851 450603 51854
rect 81433 51778 81499 51781
rect 107142 51778 107148 51780
rect 81433 51776 107148 51778
rect 81433 51720 81438 51776
rect 81494 51720 107148 51776
rect 81433 51718 107148 51720
rect 81433 51715 81499 51718
rect 107142 51716 107148 51718
rect 107212 51716 107218 51780
rect 174854 51716 174860 51780
rect 174924 51778 174930 51780
rect 208485 51778 208551 51781
rect 542353 51778 542419 51781
rect 174924 51776 542419 51778
rect 174924 51720 208490 51776
rect 208546 51720 542358 51776
rect 542414 51720 542419 51776
rect 174924 51718 542419 51720
rect 174924 51716 174930 51718
rect 208485 51715 208551 51718
rect 542353 51715 542419 51718
rect 99465 50962 99531 50965
rect 100661 50962 100727 50965
rect 133822 50962 133828 50964
rect 99465 50960 133828 50962
rect 99465 50904 99470 50960
rect 99526 50904 100666 50960
rect 100722 50904 133828 50960
rect 99465 50902 133828 50904
rect 99465 50899 99531 50902
rect 100661 50899 100727 50902
rect 133822 50900 133828 50902
rect 133892 50900 133898 50964
rect 160686 50900 160692 50964
rect 160756 50962 160762 50964
rect 216949 50962 217015 50965
rect 160756 50960 219450 50962
rect 160756 50904 216954 50960
rect 217010 50904 219450 50960
rect 160756 50902 219450 50904
rect 160756 50900 160762 50902
rect 216949 50899 217015 50902
rect 176326 50764 176332 50828
rect 176396 50826 176402 50828
rect 209814 50826 209820 50828
rect 176396 50766 209820 50826
rect 176396 50764 176402 50766
rect 209814 50764 209820 50766
rect 209884 50826 209890 50828
rect 211102 50826 211108 50828
rect 209884 50766 211108 50826
rect 209884 50764 209890 50766
rect 211102 50764 211108 50766
rect 211172 50764 211178 50828
rect 165286 50628 165292 50692
rect 165356 50690 165362 50692
rect 198733 50690 198799 50693
rect 165356 50688 200130 50690
rect 165356 50632 198738 50688
rect 198794 50632 200130 50688
rect 165356 50630 200130 50632
rect 165356 50628 165362 50630
rect 198733 50627 198799 50630
rect 200070 50418 200130 50630
rect 219390 50554 219450 50902
rect 373993 50554 374059 50557
rect 219390 50552 374059 50554
rect 219390 50496 373998 50552
rect 374054 50496 374059 50552
rect 219390 50494 374059 50496
rect 373993 50491 374059 50494
rect 423765 50418 423831 50421
rect 200070 50416 423831 50418
rect 200070 50360 423770 50416
rect 423826 50360 423831 50416
rect 200070 50358 423831 50360
rect 423765 50355 423831 50358
rect 30373 50282 30439 50285
rect 99465 50282 99531 50285
rect 30373 50280 99531 50282
rect 30373 50224 30378 50280
rect 30434 50224 99470 50280
rect 99526 50224 99531 50280
rect 30373 50222 99531 50224
rect 30373 50219 30439 50222
rect 99465 50219 99531 50222
rect 147070 50220 147076 50284
rect 147140 50282 147146 50284
rect 193305 50282 193371 50285
rect 147140 50280 193371 50282
rect 147140 50224 193310 50280
rect 193366 50224 193371 50280
rect 147140 50222 193371 50224
rect 147140 50220 147146 50222
rect 193305 50219 193371 50222
rect 211102 50220 211108 50284
rect 211172 50282 211178 50284
rect 560937 50282 561003 50285
rect 211172 50280 561003 50282
rect 211172 50224 560942 50280
rect 560998 50224 561003 50280
rect 211172 50222 561003 50224
rect 211172 50220 211178 50222
rect 560937 50219 561003 50222
rect 100753 49602 100819 49605
rect 102041 49602 102107 49605
rect 135662 49602 135668 49604
rect 100753 49600 135668 49602
rect 100753 49544 100758 49600
rect 100814 49544 102046 49600
rect 102102 49544 135668 49600
rect 100753 49542 135668 49544
rect 100753 49539 100819 49542
rect 102041 49539 102107 49542
rect 135662 49540 135668 49542
rect 135732 49540 135738 49604
rect 167678 49540 167684 49604
rect 167748 49602 167754 49604
rect 202413 49602 202479 49605
rect 202781 49602 202847 49605
rect 167748 49600 202847 49602
rect 167748 49544 202418 49600
rect 202474 49544 202786 49600
rect 202842 49544 202847 49600
rect 167748 49542 202847 49544
rect 167748 49540 167754 49542
rect 202413 49539 202479 49542
rect 202781 49539 202847 49542
rect 162342 49404 162348 49468
rect 162412 49466 162418 49468
rect 195973 49466 196039 49469
rect 162412 49464 196039 49466
rect 162412 49408 195978 49464
rect 196034 49408 196039 49464
rect 162412 49406 196039 49408
rect 162412 49404 162418 49406
rect 195973 49403 196039 49406
rect 158846 49268 158852 49332
rect 158916 49330 158922 49332
rect 191782 49330 191788 49332
rect 158916 49270 191788 49330
rect 158916 49268 158922 49270
rect 191782 49268 191788 49270
rect 191852 49330 191858 49332
rect 356053 49330 356119 49333
rect 191852 49328 356119 49330
rect 191852 49272 356058 49328
rect 356114 49272 356119 49328
rect 191852 49270 356119 49272
rect 191852 49268 191858 49270
rect 356053 49267 356119 49270
rect 195973 49194 196039 49197
rect 387793 49194 387859 49197
rect 195973 49192 387859 49194
rect 195973 49136 195978 49192
rect 196034 49136 387798 49192
rect 387854 49136 387859 49192
rect 195973 49134 387859 49136
rect 195973 49131 196039 49134
rect 387793 49131 387859 49134
rect 202781 49058 202847 49061
rect 455413 49058 455479 49061
rect 202781 49056 455479 49058
rect 202781 49000 202786 49056
rect 202842 49000 455418 49056
rect 455474 49000 455479 49056
rect 202781 48998 455479 49000
rect 202781 48995 202847 48998
rect 455413 48995 455479 48998
rect 39297 48922 39363 48925
rect 100753 48922 100819 48925
rect 39297 48920 100819 48922
rect 39297 48864 39302 48920
rect 39358 48864 100758 48920
rect 100814 48864 100819 48920
rect 39297 48862 100819 48864
rect 39297 48859 39363 48862
rect 100753 48859 100819 48862
rect 176510 48860 176516 48924
rect 176580 48922 176586 48924
rect 210141 48922 210207 48925
rect 556153 48922 556219 48925
rect 176580 48920 556219 48922
rect 176580 48864 210146 48920
rect 210202 48864 556158 48920
rect 556214 48864 556219 48920
rect 176580 48862 556219 48864
rect 176580 48860 176586 48862
rect 210141 48859 210207 48862
rect 556153 48859 556219 48862
rect 103278 48180 103284 48244
rect 103348 48242 103354 48244
rect 135478 48242 135484 48244
rect 103348 48182 135484 48242
rect 103348 48180 103354 48182
rect 44265 47562 44331 47565
rect 103470 47562 103530 48182
rect 135478 48180 135484 48182
rect 135548 48180 135554 48244
rect 169334 48180 169340 48244
rect 169404 48242 169410 48244
rect 203333 48242 203399 48245
rect 204161 48242 204227 48245
rect 169404 48240 204227 48242
rect 169404 48184 203338 48240
rect 203394 48184 204166 48240
rect 204222 48184 204227 48240
rect 169404 48182 204227 48184
rect 169404 48180 169410 48182
rect 203333 48179 203399 48182
rect 204161 48179 204227 48182
rect 163630 48044 163636 48108
rect 163700 48106 163706 48108
rect 197445 48106 197511 48109
rect 163700 48104 197511 48106
rect 163700 48048 197450 48104
rect 197506 48048 197511 48104
rect 163700 48046 197511 48048
rect 163700 48044 163706 48046
rect 197445 48043 197511 48046
rect 169518 47908 169524 47972
rect 169588 47970 169594 47972
rect 202965 47970 203031 47973
rect 204069 47970 204135 47973
rect 169588 47968 204135 47970
rect 169588 47912 202970 47968
rect 203026 47912 204074 47968
rect 204130 47912 204135 47968
rect 169588 47910 204135 47912
rect 169588 47908 169594 47910
rect 202965 47907 203031 47910
rect 204069 47907 204135 47910
rect 197445 47834 197511 47837
rect 405733 47834 405799 47837
rect 197445 47832 405799 47834
rect 197445 47776 197450 47832
rect 197506 47776 405738 47832
rect 405794 47776 405799 47832
rect 197445 47774 405799 47776
rect 197445 47771 197511 47774
rect 405733 47771 405799 47774
rect 204161 47698 204227 47701
rect 466453 47698 466519 47701
rect 204161 47696 466519 47698
rect 204161 47640 204166 47696
rect 204222 47640 466458 47696
rect 466514 47640 466519 47696
rect 204161 47638 466519 47640
rect 204161 47635 204227 47638
rect 466453 47635 466519 47638
rect 44265 47560 103530 47562
rect 44265 47504 44270 47560
rect 44326 47504 103530 47560
rect 44265 47502 103530 47504
rect 204069 47562 204135 47565
rect 468477 47562 468543 47565
rect 204069 47560 468543 47562
rect 204069 47504 204074 47560
rect 204130 47504 468482 47560
rect 468538 47504 468543 47560
rect 204069 47502 468543 47504
rect 44265 47499 44331 47502
rect 204069 47499 204135 47502
rect 468477 47499 468543 47502
rect 100753 46882 100819 46885
rect 101581 46882 101647 46885
rect 135294 46882 135300 46884
rect 100753 46880 135300 46882
rect 100753 46824 100758 46880
rect 100814 46824 101586 46880
rect 101642 46824 135300 46880
rect 100753 46822 135300 46824
rect 100753 46819 100819 46822
rect 101581 46819 101647 46822
rect 135294 46820 135300 46822
rect 135364 46820 135370 46884
rect 152590 46820 152596 46884
rect 152660 46882 152666 46884
rect 220905 46882 220971 46885
rect 152660 46880 229110 46882
rect 152660 46824 220910 46880
rect 220966 46824 229110 46880
rect 152660 46822 229110 46824
rect 152660 46820 152666 46822
rect 220905 46819 220971 46822
rect 165470 46684 165476 46748
rect 165540 46746 165546 46748
rect 219433 46746 219499 46749
rect 165540 46744 219499 46746
rect 165540 46688 219438 46744
rect 219494 46688 219499 46744
rect 165540 46686 219499 46688
rect 165540 46684 165546 46686
rect 219390 46683 219499 46686
rect 170990 46548 170996 46612
rect 171060 46610 171066 46612
rect 171060 46550 200130 46610
rect 171060 46548 171066 46550
rect 49693 46202 49759 46205
rect 100753 46202 100819 46205
rect 49693 46200 100819 46202
rect 49693 46144 49698 46200
rect 49754 46144 100758 46200
rect 100814 46144 100819 46200
rect 49693 46142 100819 46144
rect 49693 46139 49759 46142
rect 100753 46139 100819 46142
rect 144494 46140 144500 46204
rect 144564 46202 144570 46204
rect 151905 46202 151971 46205
rect 144564 46200 151971 46202
rect 144564 46144 151910 46200
rect 151966 46144 151971 46200
rect 144564 46142 151971 46144
rect 200070 46202 200130 46550
rect 219390 46338 219450 46683
rect 229050 46474 229110 46822
rect 259545 46474 259611 46477
rect 229050 46472 259611 46474
rect 229050 46416 259550 46472
rect 259606 46416 259611 46472
rect 229050 46414 259611 46416
rect 259545 46411 259611 46414
rect 425053 46338 425119 46341
rect 219390 46336 425119 46338
rect 219390 46280 425058 46336
rect 425114 46280 425119 46336
rect 219390 46278 425119 46280
rect 425053 46275 425119 46278
rect 580533 46338 580599 46341
rect 583520 46338 584960 46428
rect 580533 46336 584960 46338
rect 580533 46280 580538 46336
rect 580594 46280 584960 46336
rect 580533 46278 584960 46280
rect 580533 46275 580599 46278
rect 204713 46202 204779 46205
rect 484393 46202 484459 46205
rect 200070 46200 484459 46202
rect 200070 46144 204718 46200
rect 204774 46144 484398 46200
rect 484454 46144 484459 46200
rect 583520 46188 584960 46278
rect 200070 46142 484459 46144
rect 144564 46140 144570 46142
rect 151905 46139 151971 46142
rect 204713 46139 204779 46142
rect 484393 46139 484459 46142
rect -960 45522 480 45612
rect 205909 45524 205975 45525
rect -960 45462 674 45522
rect -960 45386 480 45462
rect 614 45386 674 45462
rect 108614 45460 108620 45524
rect 108684 45522 108690 45524
rect 139526 45522 139532 45524
rect 108684 45462 139532 45522
rect 108684 45460 108690 45462
rect 139526 45460 139532 45462
rect 139596 45460 139602 45524
rect 162526 45460 162532 45524
rect 162596 45522 162602 45524
rect 196014 45522 196020 45524
rect 162596 45462 196020 45522
rect 162596 45460 162602 45462
rect 196014 45460 196020 45462
rect 196084 45460 196090 45524
rect 205909 45520 205956 45524
rect 206020 45522 206026 45524
rect 205909 45464 205914 45520
rect 205909 45460 205956 45464
rect 206020 45462 206066 45522
rect 206020 45460 206026 45462
rect 205909 45459 205975 45460
rect -960 45372 674 45386
rect 246 45326 674 45372
rect 246 44842 306 45326
rect 166758 45324 166764 45388
rect 166828 45386 166834 45388
rect 200205 45386 200271 45389
rect 201401 45386 201467 45389
rect 166828 45384 201467 45386
rect 166828 45328 200210 45384
rect 200266 45328 201406 45384
rect 201462 45328 201467 45384
rect 166828 45326 201467 45328
rect 166828 45324 166834 45326
rect 200205 45323 200271 45326
rect 201401 45323 201467 45326
rect 149830 45188 149836 45252
rect 149900 45250 149906 45252
rect 231853 45250 231919 45253
rect 149900 45248 231919 45250
rect 149900 45192 231858 45248
rect 231914 45192 231919 45248
rect 149900 45190 231919 45192
rect 149900 45188 149906 45190
rect 231853 45187 231919 45190
rect 196014 45052 196020 45116
rect 196084 45114 196090 45116
rect 390553 45114 390619 45117
rect 196084 45112 390619 45114
rect 196084 45056 390558 45112
rect 390614 45056 390619 45112
rect 196084 45054 390619 45056
rect 196084 45052 196090 45054
rect 390553 45051 390619 45054
rect 201401 44978 201467 44981
rect 444373 44978 444439 44981
rect 201401 44976 444439 44978
rect 201401 44920 201406 44976
rect 201462 44920 444378 44976
rect 444434 44920 444439 44976
rect 201401 44918 444439 44920
rect 201401 44915 201467 44918
rect 444373 44915 444439 44918
rect 95233 44842 95299 44845
rect 108614 44842 108620 44844
rect 246 44782 6930 44842
rect 6870 44298 6930 44782
rect 95233 44840 108620 44842
rect 95233 44784 95238 44840
rect 95294 44784 108620 44840
rect 95233 44782 108620 44784
rect 95233 44779 95299 44782
rect 108614 44780 108620 44782
rect 108684 44780 108690 44844
rect 173750 44780 173756 44844
rect 173820 44842 173826 44844
rect 207054 44842 207060 44844
rect 173820 44782 207060 44842
rect 173820 44780 173826 44782
rect 207054 44780 207060 44782
rect 207124 44842 207130 44844
rect 528553 44842 528619 44845
rect 207124 44840 528619 44842
rect 207124 44784 528558 44840
rect 528614 44784 528619 44840
rect 207124 44782 528619 44784
rect 207124 44780 207130 44782
rect 528553 44779 528619 44782
rect 116526 44298 116532 44300
rect 6870 44238 116532 44298
rect 116526 44236 116532 44238
rect 116596 44236 116602 44300
rect 102133 44162 102199 44165
rect 102685 44162 102751 44165
rect 136582 44162 136588 44164
rect 102133 44160 136588 44162
rect 102133 44104 102138 44160
rect 102194 44104 102690 44160
rect 102746 44104 136588 44160
rect 102133 44102 136588 44104
rect 102133 44099 102199 44102
rect 102685 44099 102751 44102
rect 136582 44100 136588 44102
rect 136652 44100 136658 44164
rect 175038 44100 175044 44164
rect 175108 44162 175114 44164
rect 208393 44162 208459 44165
rect 175108 44160 208459 44162
rect 175108 44104 208398 44160
rect 208454 44104 208459 44160
rect 175108 44102 208459 44104
rect 175108 44100 175114 44102
rect 208393 44099 208459 44102
rect 209998 44100 210004 44164
rect 210068 44162 210074 44164
rect 210141 44162 210207 44165
rect 210068 44160 210207 44162
rect 210068 44104 210146 44160
rect 210202 44104 210207 44160
rect 210068 44102 210207 44104
rect 210068 44100 210074 44102
rect 210141 44099 210207 44102
rect 63493 43482 63559 43485
rect 102133 43482 102199 43485
rect 63493 43480 102199 43482
rect 63493 43424 63498 43480
rect 63554 43424 102138 43480
rect 102194 43424 102199 43480
rect 63493 43422 102199 43424
rect 63493 43419 63559 43422
rect 102133 43419 102199 43422
rect 146886 43420 146892 43484
rect 146956 43482 146962 43484
rect 191833 43482 191899 43485
rect 146956 43480 191899 43482
rect 146956 43424 191838 43480
rect 191894 43424 191899 43480
rect 146956 43422 191899 43424
rect 146956 43420 146962 43422
rect 191833 43419 191899 43422
rect 208393 43482 208459 43485
rect 549253 43482 549319 43485
rect 208393 43480 549319 43482
rect 208393 43424 208398 43480
rect 208454 43424 549258 43480
rect 549314 43424 549319 43480
rect 208393 43422 549319 43424
rect 208393 43419 208459 43422
rect 549253 43419 549319 43422
rect 96245 41306 96311 41309
rect 96521 41306 96587 41309
rect 138054 41306 138060 41308
rect 96245 41304 138060 41306
rect 96245 41248 96250 41304
rect 96306 41248 96526 41304
rect 96582 41248 138060 41304
rect 96245 41246 138060 41248
rect 96245 41243 96311 41246
rect 96521 41243 96587 41246
rect 138054 41244 138060 41246
rect 138124 41244 138130 41308
rect 158110 41244 158116 41308
rect 158180 41306 158186 41308
rect 204713 41306 204779 41309
rect 158180 41304 204779 41306
rect 158180 41248 204718 41304
rect 204774 41248 204779 41304
rect 158180 41246 204779 41248
rect 158180 41244 158186 41246
rect 204713 41243 204779 41246
rect 149646 40700 149652 40764
rect 149716 40762 149722 40764
rect 229093 40762 229159 40765
rect 149716 40760 229159 40762
rect 149716 40704 229098 40760
rect 229154 40704 229159 40760
rect 149716 40702 229159 40704
rect 149716 40700 149722 40702
rect 229093 40699 229159 40702
rect 74533 40626 74599 40629
rect 96521 40626 96587 40629
rect 74533 40624 96587 40626
rect 74533 40568 74538 40624
rect 74594 40568 96526 40624
rect 96582 40568 96587 40624
rect 74533 40566 96587 40568
rect 74533 40563 74599 40566
rect 96521 40563 96587 40566
rect 204713 40626 204779 40629
rect 324313 40626 324379 40629
rect 204713 40624 324379 40626
rect 204713 40568 204718 40624
rect 204774 40568 324318 40624
rect 324374 40568 324379 40624
rect 204713 40566 324379 40568
rect 204713 40563 204779 40566
rect 324313 40563 324379 40566
rect 153878 39884 153884 39948
rect 153948 39946 153954 39948
rect 191925 39946 191991 39949
rect 193029 39946 193095 39949
rect 153948 39944 193095 39946
rect 153948 39888 191930 39944
rect 191986 39888 193034 39944
rect 193090 39888 193095 39944
rect 153948 39886 193095 39888
rect 153948 39884 153954 39886
rect 191925 39883 191991 39886
rect 193029 39883 193095 39886
rect 193029 39266 193095 39269
rect 276105 39266 276171 39269
rect 193029 39264 276171 39266
rect 193029 39208 193034 39264
rect 193090 39208 276110 39264
rect 276166 39208 276171 39264
rect 193029 39206 276171 39208
rect 193029 39203 193095 39206
rect 276105 39203 276171 39206
rect 155718 38524 155724 38588
rect 155788 38586 155794 38588
rect 216857 38586 216923 38589
rect 217041 38586 217107 38589
rect 155788 38584 217107 38586
rect 155788 38528 216862 38584
rect 216918 38528 217046 38584
rect 217102 38528 217107 38584
rect 155788 38526 217107 38528
rect 155788 38524 155794 38526
rect 216857 38523 216923 38526
rect 217041 38523 217107 38526
rect 217041 37906 217107 37909
rect 293953 37906 294019 37909
rect 217041 37904 294019 37906
rect 217041 37848 217046 37904
rect 217102 37848 293958 37904
rect 294014 37848 294019 37904
rect 217041 37846 294019 37848
rect 217041 37843 217107 37846
rect 293953 37843 294019 37846
rect 96429 37226 96495 37229
rect 102133 37226 102199 37229
rect 96429 37224 102199 37226
rect 96429 37168 96434 37224
rect 96490 37168 102138 37224
rect 102194 37168 102199 37224
rect 96429 37166 102199 37168
rect 96429 37163 96495 37166
rect 102133 37163 102199 37166
rect 102133 36546 102199 36549
rect 139342 36546 139348 36548
rect 102133 36544 139348 36546
rect 102133 36488 102138 36544
rect 102194 36488 139348 36544
rect 102133 36486 139348 36488
rect 102133 36483 102199 36486
rect 139342 36484 139348 36486
rect 139412 36484 139418 36548
rect 157006 35804 157012 35868
rect 157076 35866 157082 35868
rect 204805 35866 204871 35869
rect 157076 35864 204871 35866
rect 157076 35808 204810 35864
rect 204866 35808 204871 35864
rect 157076 35806 204871 35808
rect 157076 35804 157082 35806
rect 204805 35803 204871 35806
rect 167862 35668 167868 35732
rect 167932 35730 167938 35732
rect 214097 35730 214163 35733
rect 167932 35728 214163 35730
rect 167932 35672 214102 35728
rect 214158 35672 214163 35728
rect 167932 35670 214163 35672
rect 167932 35668 167938 35670
rect 214097 35667 214163 35670
rect 204805 35322 204871 35325
rect 303613 35322 303679 35325
rect 204805 35320 303679 35322
rect 204805 35264 204810 35320
rect 204866 35264 303618 35320
rect 303674 35264 303679 35320
rect 204805 35262 303679 35264
rect 204805 35259 204871 35262
rect 303613 35259 303679 35262
rect 214097 35186 214163 35189
rect 454033 35186 454099 35189
rect 214097 35184 454099 35186
rect 214097 35128 214102 35184
rect 214158 35128 454038 35184
rect 454094 35128 454099 35184
rect 214097 35126 454099 35128
rect 214097 35123 214163 35126
rect 454033 35123 454099 35126
rect 168046 33084 168052 33148
rect 168116 33146 168122 33148
rect 215569 33146 215635 33149
rect 168116 33144 215635 33146
rect 168116 33088 215574 33144
rect 215630 33088 215635 33144
rect 168116 33086 215635 33088
rect 168116 33084 168122 33086
rect 215569 33083 215635 33086
rect 580441 33146 580507 33149
rect 583520 33146 584960 33236
rect 580441 33144 584960 33146
rect 580441 33088 580446 33144
rect 580502 33088 584960 33144
rect 580441 33086 584960 33088
rect 580441 33083 580507 33086
rect 162710 32948 162716 33012
rect 162780 33010 162786 33012
rect 209865 33010 209931 33013
rect 162780 33008 209931 33010
rect 162780 32952 209870 33008
rect 209926 32952 209931 33008
rect 583520 32996 584960 33086
rect 162780 32950 209931 32952
rect 162780 32948 162786 32950
rect 209730 32602 209790 32950
rect 209865 32947 209931 32950
rect 390645 32602 390711 32605
rect 209730 32600 390711 32602
rect -960 32466 480 32556
rect 209730 32544 390650 32600
rect 390706 32544 390711 32600
rect 209730 32542 390711 32544
rect 390645 32539 390711 32542
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 215569 32466 215635 32469
rect 456793 32466 456859 32469
rect 215569 32464 456859 32466
rect 215569 32408 215574 32464
rect 215630 32408 456798 32464
rect 456854 32408 456859 32464
rect 215569 32406 456859 32408
rect 215569 32403 215635 32406
rect 456793 32403 456859 32406
rect 148358 30908 148364 30972
rect 148428 30970 148434 30972
rect 208393 30970 208459 30973
rect 148428 30968 208459 30970
rect 148428 30912 208398 30968
rect 208454 30912 208459 30968
rect 148428 30910 208459 30912
rect 148428 30908 148434 30910
rect 208393 30907 208459 30910
rect 158294 30228 158300 30292
rect 158364 30290 158370 30292
rect 205725 30290 205791 30293
rect 206001 30290 206067 30293
rect 158364 30288 206067 30290
rect 158364 30232 205730 30288
rect 205786 30232 206006 30288
rect 206062 30232 206067 30288
rect 158364 30230 206067 30232
rect 158364 30228 158370 30230
rect 205725 30227 205791 30230
rect 206001 30227 206067 30230
rect 205725 29610 205791 29613
rect 333973 29610 334039 29613
rect 205725 29608 334039 29610
rect 205725 29552 205730 29608
rect 205786 29552 333978 29608
rect 334034 29552 334039 29608
rect 205725 29550 334039 29552
rect 205725 29547 205791 29550
rect 333973 29547 334039 29550
rect 148174 28188 148180 28252
rect 148244 28250 148250 28252
rect 212533 28250 212599 28253
rect 148244 28248 212599 28250
rect 148244 28192 212538 28248
rect 212594 28192 212599 28248
rect 148244 28190 212599 28192
rect 148244 28188 148250 28190
rect 212533 28187 212599 28190
rect 145414 22612 145420 22676
rect 145484 22674 145490 22676
rect 173157 22674 173223 22677
rect 145484 22672 173223 22674
rect 145484 22616 173162 22672
rect 173218 22616 173223 22672
rect 145484 22614 173223 22616
rect 145484 22612 145490 22614
rect 173157 22611 173223 22614
rect 157926 21932 157932 21996
rect 157996 21994 158002 21996
rect 216673 21994 216739 21997
rect 157996 21992 219450 21994
rect 157996 21936 216678 21992
rect 216734 21936 219450 21992
rect 157996 21934 219450 21936
rect 157996 21932 158002 21934
rect 216673 21931 216739 21934
rect 159030 21796 159036 21860
rect 159100 21858 159106 21860
rect 207013 21858 207079 21861
rect 159100 21856 209790 21858
rect 159100 21800 207018 21856
rect 207074 21800 209790 21856
rect 159100 21798 209790 21800
rect 159100 21796 159106 21798
rect 207013 21795 207079 21798
rect 163446 21660 163452 21724
rect 163516 21722 163522 21724
rect 163516 21662 200130 21722
rect 163516 21660 163522 21662
rect 200070 21314 200130 21662
rect 209730 21450 209790 21798
rect 219390 21586 219450 21934
rect 336733 21586 336799 21589
rect 219390 21584 336799 21586
rect 219390 21528 336738 21584
rect 336794 21528 336799 21584
rect 219390 21526 336799 21528
rect 336733 21523 336799 21526
rect 342989 21450 343055 21453
rect 209730 21448 343055 21450
rect 209730 21392 342994 21448
rect 343050 21392 343055 21448
rect 209730 21390 343055 21392
rect 342989 21387 343055 21390
rect 209773 21314 209839 21317
rect 347773 21314 347839 21317
rect 200070 21312 347839 21314
rect 200070 21256 209778 21312
rect 209834 21256 347778 21312
rect 347834 21256 347839 21312
rect 200070 21254 347839 21256
rect 209773 21251 209839 21254
rect 347773 21251 347839 21254
rect 580349 19818 580415 19821
rect 583520 19818 584960 19908
rect 580349 19816 584960 19818
rect 580349 19760 580354 19816
rect 580410 19760 584960 19816
rect 580349 19758 584960 19760
rect 580349 19755 580415 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 152406 18532 152412 18596
rect 152476 18594 152482 18596
rect 266353 18594 266419 18597
rect 152476 18592 266419 18594
rect 152476 18536 266358 18592
rect 266414 18536 266419 18592
rect 152476 18534 266419 18536
rect 152476 18532 152482 18534
rect 266353 18531 266419 18534
rect 156638 17852 156644 17916
rect 156708 17914 156714 17916
rect 211153 17914 211219 17917
rect 212441 17914 212507 17917
rect 156708 17912 212507 17914
rect 156708 17856 211158 17912
rect 211214 17856 212446 17912
rect 212502 17856 212507 17912
rect 156708 17854 212507 17856
rect 156708 17852 156714 17854
rect 211153 17851 211219 17854
rect 212441 17851 212507 17854
rect 212441 17234 212507 17237
rect 316125 17234 316191 17237
rect 212441 17232 316191 17234
rect 212441 17176 212446 17232
rect 212502 17176 316130 17232
rect 316186 17176 316191 17232
rect 212441 17174 316191 17176
rect 212441 17171 212507 17174
rect 316125 17171 316191 17174
rect 144310 15812 144316 15876
rect 144380 15874 144386 15876
rect 161105 15874 161171 15877
rect 144380 15872 161171 15874
rect 144380 15816 161110 15872
rect 161166 15816 161171 15872
rect 144380 15814 161171 15816
rect 144380 15812 144386 15814
rect 161105 15811 161171 15814
rect 144126 7516 144132 7580
rect 144196 7578 144202 7580
rect 160093 7578 160159 7581
rect 144196 7576 160159 7578
rect 144196 7520 160098 7576
rect 160154 7520 160159 7576
rect 144196 7518 160159 7520
rect 144196 7516 144202 7518
rect 160093 7515 160159 7518
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 189028 289852 189092 289916
rect 187004 281556 187068 281620
rect 111564 265100 111628 265164
rect 111380 264964 111444 265028
rect 198780 264964 198844 265028
rect 115796 263740 115860 263804
rect 117084 263604 117148 263668
rect 109540 262516 109604 262580
rect 193444 262516 193508 262580
rect 193260 262380 193324 262444
rect 118372 260340 118436 260404
rect 114140 260204 114204 260268
rect 118556 260068 118620 260132
rect 113036 259932 113100 259996
rect 116900 259796 116964 259860
rect 113956 259660 114020 259724
rect 111196 259524 111260 259588
rect 186084 259388 186148 259452
rect 186084 212468 186148 212532
rect 137876 200636 137940 200700
rect 103100 200500 103164 200564
rect 136036 200500 136100 200564
rect 102732 200364 102796 200428
rect 171364 200364 171428 200428
rect 139348 199956 139412 200020
rect 134748 199880 134812 199884
rect 134748 199824 134752 199880
rect 134752 199824 134808 199880
rect 134808 199824 134812 199880
rect 134748 199820 134812 199824
rect 134196 199684 134260 199748
rect 135484 199858 135488 199884
rect 135488 199858 135544 199884
rect 135544 199858 135548 199884
rect 135484 199820 135548 199858
rect 136404 199858 136408 199884
rect 136408 199858 136464 199884
rect 136464 199858 136468 199884
rect 136404 199820 136468 199858
rect 136772 199858 136776 199884
rect 136776 199858 136832 199884
rect 136832 199858 136836 199884
rect 136772 199820 136836 199858
rect 136036 199684 136100 199748
rect 138244 199820 138308 199884
rect 138060 199684 138124 199748
rect 139164 199858 139168 199884
rect 139168 199858 139224 199884
rect 139224 199858 139228 199884
rect 166212 200092 166276 200156
rect 139164 199820 139228 199858
rect 140636 199858 140640 199884
rect 140640 199858 140696 199884
rect 140696 199858 140700 199884
rect 140636 199820 140700 199858
rect 141464 199914 141528 199918
rect 141464 199858 141468 199914
rect 141468 199858 141524 199914
rect 141524 199858 141528 199914
rect 137876 199548 137940 199612
rect 141464 199854 141528 199858
rect 141924 199820 141988 199884
rect 142108 199820 142172 199884
rect 142844 199858 142848 199884
rect 142848 199858 142904 199884
rect 142904 199858 142908 199884
rect 142844 199820 142908 199858
rect 143212 199820 143276 199884
rect 142660 199684 142724 199748
rect 144132 199820 144196 199884
rect 145420 199858 145424 199884
rect 145424 199858 145480 199884
rect 145480 199858 145484 199884
rect 145420 199820 145484 199858
rect 145052 199744 145116 199748
rect 145052 199688 145066 199744
rect 145066 199688 145116 199744
rect 145052 199684 145116 199688
rect 146524 199858 146528 199884
rect 146528 199858 146584 199884
rect 146584 199858 146588 199884
rect 146524 199820 146588 199858
rect 146524 199744 146588 199748
rect 146524 199688 146574 199744
rect 146574 199688 146588 199744
rect 146524 199684 146588 199688
rect 147260 199858 147264 199884
rect 147264 199858 147320 199884
rect 147320 199858 147324 199884
rect 147260 199820 147324 199858
rect 148180 199820 148244 199884
rect 152780 199820 152844 199884
rect 147628 199744 147692 199748
rect 147628 199688 147642 199744
rect 147642 199688 147692 199744
rect 147628 199684 147692 199688
rect 147812 199684 147876 199748
rect 148916 199744 148980 199748
rect 148916 199688 148930 199744
rect 148930 199688 148980 199744
rect 148916 199684 148980 199688
rect 157012 199744 157076 199748
rect 157012 199688 157016 199744
rect 157016 199688 157072 199744
rect 157072 199688 157076 199744
rect 157012 199684 157076 199688
rect 158300 199858 158304 199884
rect 158304 199858 158360 199884
rect 158360 199858 158364 199884
rect 158300 199820 158364 199858
rect 158668 199858 158672 199884
rect 158672 199858 158728 199884
rect 158728 199858 158732 199884
rect 158668 199820 158732 199858
rect 160876 199820 160940 199884
rect 161244 199880 161308 199884
rect 161244 199824 161248 199880
rect 161248 199824 161304 199880
rect 161304 199824 161308 199880
rect 161244 199820 161308 199824
rect 161244 199684 161308 199748
rect 162532 199820 162596 199884
rect 164740 199858 164744 199884
rect 164744 199858 164800 199884
rect 164800 199858 164804 199884
rect 164740 199820 164804 199858
rect 165108 199820 165172 199884
rect 165476 199858 165480 199884
rect 165480 199858 165536 199884
rect 165536 199858 165540 199884
rect 165476 199820 165540 199858
rect 165844 199880 165908 199884
rect 165844 199824 165848 199880
rect 165848 199824 165904 199880
rect 165904 199824 165908 199880
rect 165844 199820 165908 199824
rect 166580 199820 166644 199884
rect 165476 199684 165540 199748
rect 168604 199858 168608 199884
rect 168608 199858 168664 199884
rect 168664 199858 168668 199884
rect 168604 199820 168668 199858
rect 169156 199858 169160 199884
rect 169160 199858 169216 199884
rect 169216 199858 169220 199884
rect 169156 199820 169220 199858
rect 169892 199820 169956 199884
rect 163820 199608 163884 199612
rect 163820 199552 163834 199608
rect 163834 199552 163884 199608
rect 163820 199548 163884 199552
rect 166028 199548 166092 199612
rect 168052 199548 168116 199612
rect 169340 199548 169404 199612
rect 170996 199858 171000 199884
rect 171000 199858 171056 199884
rect 171056 199858 171060 199884
rect 170996 199820 171060 199858
rect 171916 199820 171980 199884
rect 172652 199820 172716 199884
rect 171548 199548 171612 199612
rect 173572 199858 173576 199884
rect 173576 199858 173632 199884
rect 173632 199858 173636 199884
rect 173572 199820 173636 199858
rect 173756 199684 173820 199748
rect 174860 199820 174924 199884
rect 176332 199820 176396 199884
rect 171364 199412 171428 199476
rect 203012 199276 203076 199340
rect 138428 198868 138492 198932
rect 145052 199140 145116 199204
rect 145420 199200 145484 199204
rect 145420 199144 145434 199200
rect 145434 199144 145484 199200
rect 145420 199140 145484 199144
rect 146340 199140 146404 199204
rect 168604 199140 168668 199204
rect 173756 199200 173820 199204
rect 173756 199144 173770 199200
rect 173770 199144 173820 199200
rect 173756 199140 173820 199144
rect 200804 199140 200868 199204
rect 205036 199004 205100 199068
rect 144316 198868 144380 198932
rect 205220 198868 205284 198932
rect 139164 198596 139228 198660
rect 146524 198596 146588 198660
rect 160692 198596 160756 198660
rect 167868 198596 167932 198660
rect 169156 198656 169220 198660
rect 169156 198600 169206 198656
rect 169206 198600 169220 198656
rect 169156 198596 169220 198600
rect 169524 198596 169588 198660
rect 124076 198460 124140 198524
rect 150020 198460 150084 198524
rect 171916 198460 171980 198524
rect 201540 198460 201604 198524
rect 106044 198324 106108 198388
rect 136404 198384 136468 198388
rect 136404 198328 136454 198384
rect 136454 198328 136468 198384
rect 136404 198324 136468 198328
rect 151492 198324 151556 198388
rect 173572 198324 173636 198388
rect 107516 198188 107580 198252
rect 141924 198188 141988 198252
rect 107332 198052 107396 198116
rect 148180 198052 148244 198116
rect 157196 198052 157260 198116
rect 102916 197916 102980 197980
rect 147444 197916 147508 197980
rect 171548 197916 171612 197980
rect 134196 197780 134260 197844
rect 202828 197780 202892 197844
rect 164740 197644 164804 197708
rect 142844 197432 142908 197436
rect 142844 197376 142858 197432
rect 142858 197376 142908 197432
rect 142844 197372 142908 197376
rect 143212 197372 143276 197436
rect 200620 197372 200684 197436
rect 165108 197236 165172 197300
rect 135484 197024 135548 197028
rect 135484 196968 135534 197024
rect 135534 196968 135548 197024
rect 135484 196964 135548 196968
rect 142108 196964 142172 197028
rect 147260 196964 147324 197028
rect 161060 196964 161124 197028
rect 134012 196828 134076 196892
rect 134748 196828 134812 196892
rect 135484 196888 135548 196892
rect 135484 196832 135498 196888
rect 135498 196832 135548 196888
rect 135484 196828 135548 196832
rect 139532 196828 139596 196892
rect 140636 196888 140700 196892
rect 140636 196832 140650 196888
rect 140650 196832 140700 196888
rect 140636 196828 140700 196832
rect 142292 196828 142356 196892
rect 161060 196888 161124 196892
rect 161060 196832 161110 196888
rect 161110 196832 161124 196888
rect 161060 196828 161124 196832
rect 196020 196828 196084 196892
rect 106780 196692 106844 196756
rect 136588 196692 136652 196756
rect 143764 196692 143828 196756
rect 160876 196752 160940 196756
rect 160876 196696 160926 196752
rect 160926 196696 160940 196752
rect 160876 196692 160940 196696
rect 165844 196692 165908 196756
rect 134196 196480 134260 196484
rect 134196 196424 134210 196480
rect 134210 196424 134260 196480
rect 134196 196420 134260 196424
rect 142476 196420 142540 196484
rect 147628 196420 147692 196484
rect 169892 196420 169956 196484
rect 166028 196344 166092 196348
rect 166028 196288 166042 196344
rect 166042 196288 166092 196344
rect 166028 196284 166092 196288
rect 135668 196012 135732 196076
rect 143580 196012 143644 196076
rect 144316 196072 144380 196076
rect 144316 196016 144330 196072
rect 144330 196016 144380 196072
rect 144316 196012 144380 196016
rect 158300 196012 158364 196076
rect 170996 196012 171060 196076
rect 135300 195876 135364 195940
rect 154068 195876 154132 195940
rect 161428 195876 161492 195940
rect 168052 195876 168116 195940
rect 170996 195936 171060 195940
rect 170996 195880 171010 195936
rect 171010 195880 171060 195936
rect 170996 195876 171060 195880
rect 201724 195876 201788 195940
rect 148916 195604 148980 195668
rect 158668 195604 158732 195668
rect 118188 194516 118252 194580
rect 122972 194380 123036 194444
rect 144132 194380 144196 194444
rect 207060 194380 207124 194444
rect 122420 194244 122484 194308
rect 152780 194244 152844 194308
rect 172652 194244 172716 194308
rect 205588 194244 205652 194308
rect 101996 194108 102060 194172
rect 205772 194108 205836 194172
rect 122604 193972 122668 194036
rect 97212 193836 97276 193900
rect 154252 193292 154316 193356
rect 147812 193156 147876 193220
rect 159036 193156 159100 193220
rect 104020 193020 104084 193084
rect 196204 193020 196268 193084
rect 187740 192884 187804 192948
rect 119844 192748 119908 192812
rect 147996 192612 148060 192676
rect 148180 192476 148244 192540
rect 108804 191524 108868 191588
rect 100524 191388 100588 191452
rect 138428 191252 138492 191316
rect 100340 191116 100404 191180
rect 162348 191116 162412 191180
rect 134012 190980 134076 191044
rect 165292 190980 165356 191044
rect 104388 190300 104452 190364
rect 104204 190164 104268 190228
rect 176332 190164 176396 190228
rect 209820 190164 209884 190228
rect 142292 190028 142356 190092
rect 174676 190028 174740 190092
rect 142476 189892 142540 189956
rect 159036 189892 159100 189956
rect 143764 189756 143828 189820
rect 157012 189756 157076 189820
rect 143580 189620 143644 189684
rect 154252 189620 154316 189684
rect 124812 189484 124876 189548
rect 138244 187580 138308 187644
rect 103284 187444 103348 187508
rect 135668 187444 135732 187508
rect 120580 187308 120644 187372
rect 99236 187172 99300 187236
rect 135484 187036 135548 187100
rect 187188 187036 187252 187100
rect 115612 186900 115676 186964
rect 167868 186900 167932 186964
rect 147628 186416 147692 186420
rect 147628 186360 147642 186416
rect 147642 186360 147692 186416
rect 147628 186356 147692 186360
rect 168052 158068 168116 158132
rect 211108 157932 211172 157996
rect 165476 155756 165540 155820
rect 154068 155620 154132 155684
rect 169340 155484 169404 155548
rect 211292 155348 211356 155412
rect 168236 155212 168300 155276
rect 139532 153716 139596 153780
rect 203196 152764 203260 152828
rect 157196 152628 157260 152692
rect 161060 152492 161124 152556
rect 112852 152356 112916 152420
rect 210004 152356 210068 152420
rect 166580 151268 166644 151332
rect 196388 151268 196452 151332
rect 104756 151132 104820 151196
rect 136772 151132 136836 151196
rect 197308 151132 197372 151196
rect 134196 150996 134260 151060
rect 160692 150996 160756 151060
rect 200988 150044 201052 150108
rect 206140 149908 206204 149972
rect 205956 149772 206020 149836
rect 207244 149636 207308 149700
rect 140820 148820 140884 148884
rect 108436 148684 108500 148748
rect 121316 148548 121380 148612
rect 193628 148548 193692 148612
rect 122052 148412 122116 148476
rect 163820 148412 163884 148476
rect 191604 148412 191668 148476
rect 135300 148276 135364 148340
rect 169524 148276 169588 148340
rect 112668 147596 112732 147660
rect 187924 147596 187988 147660
rect 142660 147460 142724 147524
rect 197676 147460 197740 147524
rect 112484 147324 112548 147388
rect 197492 147324 197556 147388
rect 108620 147188 108684 147252
rect 139348 147188 139412 147252
rect 166212 147188 166276 147252
rect 199148 147188 199212 147252
rect 110828 147052 110892 147116
rect 170996 147052 171060 147116
rect 107148 146916 107212 146980
rect 138060 146916 138124 146980
rect 150020 146916 150084 146980
rect 119660 146780 119724 146844
rect 136588 146780 136652 146844
rect 109540 146236 109604 146300
rect 115796 146100 115860 146164
rect 191788 146100 191852 146164
rect 111564 145964 111628 146028
rect 189212 145964 189276 146028
rect 113956 145828 114020 145892
rect 191972 145828 192036 145892
rect 116348 145692 116412 145756
rect 198780 145692 198844 145756
rect 111380 145556 111444 145620
rect 147444 145556 147508 145620
rect 113036 144740 113100 144804
rect 189764 144740 189828 144804
rect 118188 144604 118252 144668
rect 193260 144604 193324 144668
rect 147628 144468 147692 144532
rect 193444 144468 193508 144532
rect 118188 144332 118252 144396
rect 189028 144332 189092 144396
rect 115244 144196 115308 144260
rect 113956 144060 114020 144124
rect 187004 144060 187068 144124
rect 118372 143380 118436 143444
rect 118372 143244 118436 143308
rect 118556 143108 118620 143172
rect 117084 142972 117148 143036
rect 116900 142836 116964 142900
rect 111012 142700 111076 142764
rect 111196 142564 111260 142628
rect 189580 141476 189644 141540
rect 114140 141340 114204 141404
rect 116532 141204 116596 141268
rect 118556 140796 118620 140860
rect 193444 140660 193508 140724
rect 120028 140524 120092 140588
rect 188292 140388 188356 140452
rect 118004 140252 118068 140316
rect 130332 140252 130396 140316
rect 190684 140252 190748 140316
rect 120764 140116 120828 140180
rect 194548 140116 194612 140180
rect 109540 139980 109604 140044
rect 151492 139980 151556 140044
rect 190500 139844 190564 139908
rect 113772 139708 113836 139772
rect 192156 139708 192220 139772
rect 116716 139572 116780 139636
rect 189396 139436 189460 139500
rect 114140 139028 114204 139092
rect 130332 139028 130396 139092
rect 121132 138076 121196 138140
rect 123156 138076 123220 138140
rect 198964 138076 199028 138140
rect 122788 138000 122852 138004
rect 122788 137944 122802 138000
rect 122802 137944 122852 138000
rect 122788 137940 122852 137944
rect 187924 137940 187988 138004
rect 124812 137804 124876 137868
rect 187188 137804 187252 137868
rect 188292 137804 188356 137868
rect 105124 137260 105188 137324
rect 120580 137260 120644 137324
rect 119660 130324 119724 130388
rect 120028 130324 120092 130388
rect 122788 128480 122852 128484
rect 122788 128424 122802 128480
rect 122802 128424 122852 128480
rect 122788 128420 122852 128424
rect 123156 123388 123220 123452
rect 122788 122980 122852 123044
rect 122236 122164 122300 122228
rect 122604 122164 122668 122228
rect 191604 114412 191668 114476
rect 189580 113868 189644 113932
rect 115244 113732 115308 113796
rect 122236 113732 122300 113796
rect 122604 113732 122668 113796
rect 189396 113324 189460 113388
rect 189580 113324 189644 113388
rect 122236 112644 122300 112708
rect 122604 112644 122668 112708
rect 119476 112372 119540 112436
rect 119476 111828 119540 111892
rect 122052 111828 122116 111892
rect 122052 110604 122116 110668
rect 189396 110604 189460 110668
rect 113588 110468 113652 110532
rect 120764 110468 120828 110532
rect 189396 109244 189460 109308
rect 189396 107068 189460 107132
rect 122236 103532 122300 103596
rect 122604 103532 122668 103596
rect 122236 103124 122300 103188
rect 122604 103124 122668 103188
rect 116716 96596 116780 96660
rect 122236 94012 122300 94076
rect 122604 94012 122668 94076
rect 122236 93604 122300 93668
rect 122604 93604 122668 93668
rect 122236 84492 122300 84556
rect 122604 84492 122668 84556
rect 122788 83948 122852 84012
rect 196388 82180 196452 82244
rect 191604 81500 191668 81564
rect 105124 81424 105188 81428
rect 105124 81368 105174 81424
rect 105174 81368 105188 81424
rect 105124 81364 105188 81368
rect 124076 81228 124140 81292
rect 147812 81228 147876 81292
rect 164004 81228 164068 81292
rect 191972 81228 192036 81292
rect 175412 81092 175476 81156
rect 151308 80956 151372 81020
rect 174308 80956 174372 81020
rect 148916 80820 148980 80884
rect 172284 80820 172348 80884
rect 146340 80684 146404 80748
rect 181668 80684 181732 80748
rect 197676 80548 197740 80612
rect 113956 80412 114020 80476
rect 173020 80412 173084 80476
rect 193444 80412 193508 80476
rect 108252 80276 108316 80340
rect 135300 80004 135364 80068
rect 134196 79906 134200 79932
rect 134200 79906 134256 79932
rect 134256 79906 134260 79932
rect 134196 79868 134260 79906
rect 134564 79906 134568 79932
rect 134568 79906 134624 79932
rect 134624 79906 134628 79932
rect 134564 79868 134628 79906
rect 135852 79868 135916 79932
rect 135668 79732 135732 79796
rect 139348 80140 139412 80204
rect 136956 79906 136960 79932
rect 136960 79906 137016 79932
rect 137016 79906 137020 79932
rect 136956 79868 137020 79906
rect 137876 79928 137940 79932
rect 137876 79872 137880 79928
rect 137880 79872 137936 79928
rect 137936 79872 137940 79928
rect 137876 79868 137940 79872
rect 138612 79928 138676 79932
rect 138612 79872 138616 79928
rect 138616 79872 138672 79928
rect 138672 79872 138676 79928
rect 138612 79868 138676 79872
rect 138980 79868 139044 79932
rect 143396 80140 143460 80204
rect 147076 80140 147140 80204
rect 151676 80004 151740 80068
rect 139716 79868 139780 79932
rect 139900 79928 139964 79932
rect 139900 79872 139904 79928
rect 139904 79872 139960 79928
rect 139960 79872 139964 79928
rect 139900 79868 139964 79872
rect 140636 79868 140700 79932
rect 141188 79868 141252 79932
rect 142292 79906 142296 79932
rect 142296 79906 142352 79932
rect 142352 79906 142356 79932
rect 142292 79868 142356 79906
rect 142660 79906 142664 79932
rect 142664 79906 142720 79932
rect 142720 79906 142724 79932
rect 142660 79868 142724 79906
rect 143028 79868 143092 79932
rect 143212 79868 143276 79932
rect 143764 79906 143768 79932
rect 143768 79906 143824 79932
rect 143824 79906 143828 79932
rect 143764 79868 143828 79906
rect 144316 79868 144380 79932
rect 144684 79928 144748 79932
rect 144684 79872 144688 79928
rect 144688 79872 144744 79928
rect 144744 79872 144748 79928
rect 144684 79868 144748 79872
rect 145052 79906 145056 79932
rect 145056 79906 145112 79932
rect 145112 79906 145116 79932
rect 145052 79868 145116 79906
rect 145420 79928 145484 79932
rect 145420 79872 145424 79928
rect 145424 79872 145480 79928
rect 145480 79872 145484 79928
rect 145420 79868 145484 79872
rect 145604 79868 145668 79932
rect 146524 79868 146588 79932
rect 147628 79868 147692 79932
rect 147996 79868 148060 79932
rect 148364 79868 148428 79932
rect 149468 79868 149532 79932
rect 149652 79868 149716 79932
rect 151124 79868 151188 79932
rect 151308 79906 151312 79932
rect 151312 79906 151368 79932
rect 151368 79906 151372 79932
rect 151308 79868 151372 79906
rect 158116 80140 158180 80204
rect 158852 80004 158916 80068
rect 143028 79596 143092 79660
rect 146340 79596 146404 79660
rect 147260 79596 147324 79660
rect 147812 79596 147876 79660
rect 148916 79656 148980 79660
rect 148916 79600 148966 79656
rect 148966 79600 148980 79656
rect 148916 79596 148980 79600
rect 140820 79460 140884 79524
rect 142660 79460 142724 79524
rect 143396 79460 143460 79524
rect 144684 79460 144748 79524
rect 145052 79520 145116 79524
rect 145052 79464 145066 79520
rect 145066 79464 145116 79520
rect 145052 79460 145116 79464
rect 147812 79460 147876 79524
rect 151492 79792 151556 79796
rect 151492 79736 151496 79792
rect 151496 79736 151552 79792
rect 151552 79736 151556 79792
rect 151492 79732 151556 79736
rect 152412 79460 152476 79524
rect 153884 79928 153948 79932
rect 153884 79872 153888 79928
rect 153888 79872 153944 79928
rect 153944 79872 153948 79928
rect 153884 79868 153948 79872
rect 154252 79906 154256 79932
rect 154256 79906 154312 79932
rect 154312 79906 154316 79932
rect 154252 79868 154316 79906
rect 155724 79868 155788 79932
rect 156828 79868 156892 79932
rect 157196 79928 157260 79932
rect 157196 79872 157200 79928
rect 157200 79872 157256 79928
rect 157256 79872 157260 79928
rect 157196 79868 157260 79872
rect 158300 79868 158364 79932
rect 165108 80140 165172 80204
rect 187740 80276 187804 80340
rect 154436 79792 154500 79796
rect 154436 79736 154450 79792
rect 154450 79736 154500 79792
rect 154436 79732 154500 79736
rect 155540 79732 155604 79796
rect 158484 79732 158548 79796
rect 160876 79928 160940 79932
rect 160876 79872 160880 79928
rect 160880 79872 160936 79928
rect 160936 79872 160940 79928
rect 160876 79868 160940 79872
rect 113772 79324 113836 79388
rect 136588 79324 136652 79388
rect 139900 79324 139964 79388
rect 151308 79324 151372 79388
rect 162164 79596 162228 79660
rect 162348 79596 162412 79660
rect 163268 79868 163332 79932
rect 164004 79928 164068 79932
rect 164004 79872 164008 79928
rect 164008 79872 164064 79928
rect 164064 79872 164068 79928
rect 164004 79868 164068 79872
rect 164188 79868 164252 79932
rect 165292 79868 165356 79932
rect 165660 79928 165724 79932
rect 165660 79872 165664 79928
rect 165664 79872 165720 79928
rect 165720 79872 165724 79928
rect 165660 79868 165724 79872
rect 165844 79928 165908 79932
rect 165844 79872 165848 79928
rect 165848 79872 165904 79928
rect 165904 79872 165908 79928
rect 165844 79868 165908 79872
rect 166396 79868 166460 79932
rect 167868 79868 167932 79932
rect 166764 79732 166828 79796
rect 168052 79732 168116 79796
rect 163452 79324 163516 79388
rect 168972 79868 169036 79932
rect 170260 79868 170324 79932
rect 170076 79792 170140 79796
rect 170076 79736 170080 79792
rect 170080 79736 170136 79792
rect 170136 79736 170140 79792
rect 170076 79732 170140 79736
rect 170628 79906 170632 79932
rect 170632 79906 170688 79932
rect 170688 79906 170692 79932
rect 170628 79868 170692 79906
rect 171548 79732 171612 79796
rect 173388 79868 173452 79932
rect 172284 79732 172348 79796
rect 172836 79732 172900 79796
rect 173572 79732 173636 79796
rect 181668 80140 181732 80204
rect 175228 80004 175292 80068
rect 200804 80004 200868 80068
rect 175412 79868 175476 79932
rect 174676 79732 174740 79796
rect 176516 79868 176580 79932
rect 175964 79732 176028 79796
rect 190500 79460 190564 79524
rect 192156 79324 192220 79388
rect 146892 79188 146956 79252
rect 147628 79188 147692 79252
rect 164004 79188 164068 79252
rect 189396 79188 189460 79252
rect 190684 79052 190748 79116
rect 157012 78916 157076 78980
rect 164924 78916 164988 78980
rect 169340 78916 169404 78980
rect 173020 78916 173084 78980
rect 174308 78976 174372 78980
rect 174308 78920 174322 78976
rect 174322 78920 174372 78976
rect 174308 78916 174372 78920
rect 206140 78916 206204 78980
rect 149468 78780 149532 78844
rect 137876 78644 137940 78708
rect 140636 78644 140700 78708
rect 145420 78644 145484 78708
rect 149468 78644 149532 78708
rect 107516 78508 107580 78572
rect 149100 78508 149164 78572
rect 156644 78508 156708 78572
rect 157932 78508 157996 78572
rect 159036 78508 159100 78572
rect 160692 78508 160756 78572
rect 166580 78568 166644 78572
rect 166580 78512 166630 78568
rect 166630 78512 166644 78568
rect 166580 78508 166644 78512
rect 167500 78508 167564 78572
rect 170628 78568 170692 78572
rect 170628 78512 170642 78568
rect 170642 78512 170692 78568
rect 170628 78508 170692 78512
rect 197308 78508 197372 78572
rect 198964 78568 199028 78572
rect 198964 78512 199014 78568
rect 199014 78512 199028 78568
rect 198964 78508 199028 78512
rect 120028 78372 120092 78436
rect 122972 78372 123036 78436
rect 149284 78372 149348 78436
rect 167316 78432 167380 78436
rect 167316 78376 167366 78432
rect 167366 78376 167380 78432
rect 167316 78372 167380 78376
rect 169524 78372 169588 78436
rect 170812 78372 170876 78436
rect 172836 78372 172900 78436
rect 173388 78372 173452 78436
rect 175412 78372 175476 78436
rect 137508 78236 137572 78300
rect 139532 78236 139596 78300
rect 142292 78296 142356 78300
rect 142292 78240 142306 78296
rect 142306 78240 142356 78296
rect 142292 78236 142356 78240
rect 165476 78236 165540 78300
rect 168972 78296 169036 78300
rect 168972 78240 168986 78296
rect 168986 78240 169036 78296
rect 168972 78236 169036 78240
rect 136956 78100 137020 78164
rect 107332 77964 107396 78028
rect 134012 78024 134076 78028
rect 164188 78100 164252 78164
rect 134012 77968 134026 78024
rect 134026 77968 134076 78024
rect 134012 77964 134076 77968
rect 139900 77964 139964 78028
rect 211292 78100 211356 78164
rect 152596 77692 152660 77756
rect 171916 77752 171980 77756
rect 171916 77696 171966 77752
rect 171966 77696 171980 77752
rect 171916 77692 171980 77696
rect 173756 77692 173820 77756
rect 133460 77556 133524 77620
rect 144132 77556 144196 77620
rect 133276 77420 133340 77484
rect 135484 77420 135548 77484
rect 143580 77420 143644 77484
rect 147996 77480 148060 77484
rect 147996 77424 148010 77480
rect 148010 77424 148060 77480
rect 147996 77420 148060 77424
rect 148180 77420 148244 77484
rect 161060 77480 161124 77484
rect 211108 77828 211172 77892
rect 161060 77424 161110 77480
rect 161110 77424 161124 77480
rect 161060 77420 161124 77424
rect 133092 77284 133156 77348
rect 134564 77344 134628 77348
rect 134564 77288 134614 77344
rect 134614 77288 134628 77344
rect 134564 77284 134628 77288
rect 142844 77284 142908 77348
rect 143212 77284 143276 77348
rect 144316 77284 144380 77348
rect 147996 77284 148060 77348
rect 110828 77148 110892 77212
rect 118004 77148 118068 77212
rect 152780 77148 152844 77212
rect 154252 77148 154316 77212
rect 162532 77148 162596 77212
rect 118188 77012 118252 77076
rect 143764 77012 143828 77076
rect 143764 76876 143828 76940
rect 165292 76876 165356 76940
rect 170076 76876 170140 76940
rect 170996 76876 171060 76940
rect 174492 76876 174556 76940
rect 176148 76936 176212 76940
rect 176148 76880 176162 76936
rect 176162 76880 176212 76936
rect 176148 76876 176212 76880
rect 133828 76604 133892 76668
rect 197492 76604 197556 76668
rect 162716 76528 162780 76532
rect 162716 76472 162730 76528
rect 162730 76472 162780 76528
rect 162716 76468 162780 76472
rect 170260 76468 170324 76532
rect 170628 76468 170692 76532
rect 171732 76468 171796 76532
rect 172100 76528 172164 76532
rect 172100 76472 172150 76528
rect 172150 76472 172164 76528
rect 172100 76468 172164 76472
rect 172284 76528 172348 76532
rect 172284 76472 172334 76528
rect 172334 76472 172348 76528
rect 172284 76468 172348 76472
rect 174860 76468 174924 76532
rect 175044 76528 175108 76532
rect 175044 76472 175094 76528
rect 175094 76472 175108 76528
rect 175044 76468 175108 76472
rect 200988 76468 201052 76532
rect 140636 76196 140700 76260
rect 145604 76196 145668 76260
rect 146892 76196 146956 76260
rect 176516 76196 176580 76260
rect 138060 76120 138124 76124
rect 138060 76064 138074 76120
rect 138074 76064 138124 76120
rect 138060 76060 138124 76064
rect 138244 76060 138308 76124
rect 170444 76060 170508 76124
rect 163636 75924 163700 75988
rect 165292 75984 165356 75988
rect 165292 75928 165342 75984
rect 165342 75928 165356 75984
rect 165292 75924 165356 75928
rect 165660 75924 165724 75988
rect 167316 75924 167380 75988
rect 167684 75984 167748 75988
rect 167684 75928 167734 75984
rect 167734 75928 167748 75984
rect 167684 75924 167748 75928
rect 138980 75788 139044 75852
rect 171548 75788 171612 75852
rect 205588 75848 205652 75852
rect 205588 75792 205602 75848
rect 205602 75792 205652 75848
rect 205588 75788 205652 75792
rect 205772 75788 205836 75852
rect 147260 75652 147324 75716
rect 145420 75516 145484 75580
rect 175228 75576 175292 75580
rect 175228 75520 175242 75576
rect 175242 75520 175292 75576
rect 175228 75516 175292 75520
rect 203380 75516 203444 75580
rect 97212 75108 97276 75172
rect 138612 75108 138676 75172
rect 140820 75108 140884 75172
rect 145420 75108 145484 75172
rect 196204 75380 196268 75444
rect 199148 75244 199212 75308
rect 144316 74972 144380 75036
rect 115612 74836 115676 74900
rect 112668 74564 112732 74628
rect 119844 74428 119908 74492
rect 118372 74292 118436 74356
rect 149468 74156 149532 74220
rect 149836 74156 149900 74220
rect 152780 74292 152844 74356
rect 151124 74156 151188 74220
rect 106780 73884 106844 73948
rect 149284 73884 149348 73948
rect 103100 73748 103164 73812
rect 143028 73748 143092 73812
rect 154436 73612 154500 73676
rect 157196 73068 157260 73132
rect 158484 72932 158548 72996
rect 112484 72720 112548 72724
rect 112484 72664 112498 72720
rect 112498 72664 112548 72720
rect 112484 72660 112548 72664
rect 148364 72660 148428 72724
rect 148732 72660 148796 72724
rect 147076 71708 147140 71772
rect 207244 71572 207308 71636
rect 149284 71436 149348 71500
rect 149652 71436 149716 71500
rect 122420 71300 122484 71364
rect 152412 71300 152476 71364
rect 148180 71164 148244 71228
rect 106044 71028 106108 71092
rect 201724 71028 201788 71092
rect 144316 70212 144380 70276
rect 171732 70212 171796 70276
rect 113588 70076 113652 70140
rect 205220 70076 205284 70140
rect 118556 69940 118620 70004
rect 191604 69940 191668 70004
rect 102732 69864 102796 69868
rect 102732 69808 102782 69864
rect 102782 69808 102796 69864
rect 102732 69804 102796 69808
rect 121316 69804 121380 69868
rect 205220 69532 205284 69596
rect 102916 68852 102980 68916
rect 114140 68852 114204 68916
rect 147996 68852 148060 68916
rect 148548 68852 148612 68916
rect 112852 68716 112916 68780
rect 146524 68716 146588 68780
rect 149100 68580 149164 68644
rect 150020 68580 150084 68644
rect 122052 68444 122116 68508
rect 147812 68444 147876 68508
rect 148180 68444 148244 68508
rect 203196 68172 203260 68236
rect 119660 67492 119724 67556
rect 189212 67492 189276 67556
rect 205036 67492 205100 67556
rect 99236 66812 99300 66876
rect 133460 67356 133524 67420
rect 187740 67356 187804 67420
rect 149468 66812 149532 66876
rect 104388 66192 104452 66196
rect 104388 66136 104438 66192
rect 104438 66136 104452 66192
rect 104388 66132 104452 66136
rect 143948 66132 144012 66196
rect 144684 66132 144748 66196
rect 155540 66132 155604 66196
rect 122604 65996 122668 66060
rect 170444 65996 170508 66060
rect 143764 65860 143828 65924
rect 171916 65860 171980 65924
rect 108252 65452 108316 65516
rect 141004 65452 141068 65516
rect 147260 65452 147324 65516
rect 143580 64772 143644 64836
rect 116348 64636 116412 64700
rect 172100 64772 172164 64836
rect 121132 64500 121196 64564
rect 104204 64228 104268 64292
rect 104020 64152 104084 64156
rect 200620 64772 200684 64836
rect 104020 64096 104034 64152
rect 104034 64096 104084 64152
rect 104020 64092 104084 64096
rect 143580 63548 143644 63612
rect 144500 63548 144564 63612
rect 151492 63412 151556 63476
rect 175964 63276 176028 63340
rect 166212 63140 166276 63204
rect 172284 62868 172348 62932
rect 201540 62868 201604 62932
rect 148732 62732 148796 62796
rect 134196 62052 134260 62116
rect 164924 62052 164988 62116
rect 138612 61916 138676 61980
rect 176148 61916 176212 61980
rect 203012 61916 203076 61980
rect 204116 61916 204180 61980
rect 140820 61780 140884 61844
rect 150020 61644 150084 61708
rect 204116 61372 204180 61436
rect 193628 60616 193692 60620
rect 193628 60560 193678 60616
rect 193678 60560 193692 60616
rect 193628 60556 193692 60560
rect 173572 60420 173636 60484
rect 165108 60284 165172 60348
rect 108804 58516 108868 58580
rect 139900 59196 139964 59260
rect 151676 59196 151740 59260
rect 154068 59060 154132 59124
rect 170628 58924 170692 58988
rect 174492 58788 174556 58852
rect 111012 57972 111076 58036
rect 138428 57836 138492 57900
rect 174676 57836 174740 57900
rect 101996 57156 102060 57220
rect 134012 57700 134076 57764
rect 166396 57700 166460 57764
rect 99420 56476 99484 56540
rect 100340 56476 100404 56540
rect 133276 56476 133340 56540
rect 144684 56476 144748 56540
rect 104756 56340 104820 56404
rect 137508 56340 137572 56404
rect 99420 55796 99484 55860
rect 135852 55116 135916 55180
rect 156828 55116 156892 55180
rect 170812 54980 170876 55044
rect 160876 54844 160940 54908
rect 109540 54632 109604 54636
rect 109540 54576 109590 54632
rect 109590 54576 109604 54632
rect 109540 54572 109604 54576
rect 148548 54436 148612 54500
rect 139716 53756 139780 53820
rect 154252 53756 154316 53820
rect 100524 53620 100588 53684
rect 133092 53620 133156 53684
rect 162164 53620 162228 53684
rect 166580 53484 166644 53548
rect 194548 53484 194612 53548
rect 100524 53076 100588 53140
rect 194548 53076 194612 53140
rect 107148 52396 107212 52460
rect 138244 52396 138308 52460
rect 163268 52396 163332 52460
rect 167500 52260 167564 52324
rect 161060 52124 161124 52188
rect 189764 51988 189828 52052
rect 107148 51716 107212 51780
rect 174860 51716 174924 51780
rect 133828 50900 133892 50964
rect 160692 50900 160756 50964
rect 176332 50764 176396 50828
rect 209820 50764 209884 50828
rect 211108 50764 211172 50828
rect 165292 50628 165356 50692
rect 147076 50220 147140 50284
rect 211108 50220 211172 50284
rect 135668 49540 135732 49604
rect 167684 49540 167748 49604
rect 162348 49404 162412 49468
rect 158852 49268 158916 49332
rect 191788 49268 191852 49332
rect 176516 48860 176580 48924
rect 103284 48180 103348 48244
rect 135484 48180 135548 48244
rect 169340 48180 169404 48244
rect 163636 48044 163700 48108
rect 169524 47908 169588 47972
rect 135300 46820 135364 46884
rect 152596 46820 152660 46884
rect 165476 46684 165540 46748
rect 170996 46548 171060 46612
rect 144500 46140 144564 46204
rect 108620 45460 108684 45524
rect 139532 45460 139596 45524
rect 162532 45460 162596 45524
rect 196020 45460 196084 45524
rect 205956 45520 206020 45524
rect 205956 45464 205970 45520
rect 205970 45464 206020 45520
rect 205956 45460 206020 45464
rect 166764 45324 166828 45388
rect 149836 45188 149900 45252
rect 196020 45052 196084 45116
rect 108620 44780 108684 44844
rect 173756 44780 173820 44844
rect 207060 44780 207124 44844
rect 116532 44236 116596 44300
rect 136588 44100 136652 44164
rect 175044 44100 175108 44164
rect 210004 44100 210068 44164
rect 146892 43420 146956 43484
rect 138060 41244 138124 41308
rect 158116 41244 158180 41308
rect 149652 40700 149716 40764
rect 153884 39884 153948 39948
rect 155724 38524 155788 38588
rect 139348 36484 139412 36548
rect 157012 35804 157076 35868
rect 167868 35668 167932 35732
rect 168052 33084 168116 33148
rect 162716 32948 162780 33012
rect 148364 30908 148428 30972
rect 158300 30228 158364 30292
rect 148180 28188 148244 28252
rect 145420 22612 145484 22676
rect 157932 21932 157996 21996
rect 159036 21796 159100 21860
rect 163452 21660 163516 21724
rect 152412 18532 152476 18596
rect 156644 17852 156708 17916
rect 144316 15812 144380 15876
rect 144132 7516 144196 7580
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 97211 193900 97277 193901
rect 97211 193836 97212 193900
rect 97276 193836 97277 193900
rect 97211 193835 97277 193836
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 97214 75173 97274 193835
rect 100523 191452 100589 191453
rect 100523 191388 100524 191452
rect 100588 191388 100589 191452
rect 100523 191387 100589 191388
rect 100339 191180 100405 191181
rect 100339 191116 100340 191180
rect 100404 191116 100405 191180
rect 100339 191115 100405 191116
rect 99235 187236 99301 187237
rect 99235 187172 99236 187236
rect 99300 187172 99301 187236
rect 99235 187171 99301 187172
rect 97211 75172 97277 75173
rect 97211 75108 97212 75172
rect 97276 75108 97277 75172
rect 97211 75107 97277 75108
rect 99238 66877 99298 187171
rect 99235 66876 99301 66877
rect 99235 66812 99236 66876
rect 99300 66812 99301 66876
rect 99235 66811 99301 66812
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 100342 56541 100402 191115
rect 99419 56540 99485 56541
rect 99419 56476 99420 56540
rect 99484 56476 99485 56540
rect 99419 56475 99485 56476
rect 100339 56540 100405 56541
rect 100339 56476 100340 56540
rect 100404 56476 100405 56540
rect 100339 56475 100405 56476
rect 99422 55861 99482 56475
rect 99419 55860 99485 55861
rect 99419 55796 99420 55860
rect 99484 55796 99485 55860
rect 99419 55795 99485 55796
rect 100526 53685 100586 191387
rect 100794 174454 101414 209898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109539 262580 109605 262581
rect 109539 262516 109540 262580
rect 109604 262516 109605 262580
rect 109539 262515 109605 262516
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 103099 200564 103165 200565
rect 103099 200500 103100 200564
rect 103164 200500 103165 200564
rect 103099 200499 103165 200500
rect 102731 200428 102797 200429
rect 102731 200364 102732 200428
rect 102796 200364 102797 200428
rect 102731 200363 102797 200364
rect 101995 194172 102061 194173
rect 101995 194108 101996 194172
rect 102060 194108 102061 194172
rect 101995 194107 102061 194108
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100523 53684 100589 53685
rect 100523 53620 100524 53684
rect 100588 53620 100589 53684
rect 100523 53619 100589 53620
rect 100526 53141 100586 53619
rect 100523 53140 100589 53141
rect 100523 53076 100524 53140
rect 100588 53076 100589 53140
rect 100523 53075 100589 53076
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 30454 101414 65898
rect 101998 57221 102058 194107
rect 102734 69869 102794 200363
rect 102915 197980 102981 197981
rect 102915 197916 102916 197980
rect 102980 197916 102981 197980
rect 102915 197915 102981 197916
rect 102731 69868 102797 69869
rect 102731 69804 102732 69868
rect 102796 69804 102797 69868
rect 102731 69803 102797 69804
rect 102918 68917 102978 197915
rect 103102 73813 103162 200499
rect 104019 193084 104085 193085
rect 104019 193020 104020 193084
rect 104084 193020 104085 193084
rect 104019 193019 104085 193020
rect 103283 187508 103349 187509
rect 103283 187444 103284 187508
rect 103348 187444 103349 187508
rect 103283 187443 103349 187444
rect 103099 73812 103165 73813
rect 103099 73748 103100 73812
rect 103164 73748 103165 73812
rect 103099 73747 103165 73748
rect 102915 68916 102981 68917
rect 102915 68852 102916 68916
rect 102980 68852 102981 68916
rect 102915 68851 102981 68852
rect 101995 57220 102061 57221
rect 101995 57156 101996 57220
rect 102060 57156 102061 57220
rect 101995 57155 102061 57156
rect 103286 48245 103346 187443
rect 104022 64157 104082 193019
rect 104387 190364 104453 190365
rect 104387 190300 104388 190364
rect 104452 190300 104453 190364
rect 104387 190299 104453 190300
rect 104203 190228 104269 190229
rect 104203 190164 104204 190228
rect 104268 190164 104269 190228
rect 104203 190163 104269 190164
rect 104206 64293 104266 190163
rect 104390 66197 104450 190299
rect 105294 178954 105914 214398
rect 106043 198388 106109 198389
rect 106043 198324 106044 198388
rect 106108 198324 106109 198388
rect 106043 198323 106109 198324
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 104755 151196 104821 151197
rect 104755 151132 104756 151196
rect 104820 151132 104821 151196
rect 104755 151131 104821 151132
rect 104387 66196 104453 66197
rect 104387 66132 104388 66196
rect 104452 66132 104453 66196
rect 104387 66131 104453 66132
rect 104203 64292 104269 64293
rect 104203 64228 104204 64292
rect 104268 64228 104269 64292
rect 104203 64227 104269 64228
rect 104019 64156 104085 64157
rect 104019 64092 104020 64156
rect 104084 64092 104085 64156
rect 104019 64091 104085 64092
rect 104758 56405 104818 151131
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105123 137324 105189 137325
rect 105123 137260 105124 137324
rect 105188 137260 105189 137324
rect 105123 137259 105189 137260
rect 105126 81429 105186 137259
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105123 81428 105189 81429
rect 105123 81364 105124 81428
rect 105188 81364 105189 81428
rect 105123 81363 105189 81364
rect 105294 70954 105914 106398
rect 106046 71093 106106 198323
rect 107515 198252 107581 198253
rect 107515 198188 107516 198252
rect 107580 198188 107581 198252
rect 107515 198187 107581 198188
rect 107331 198116 107397 198117
rect 107331 198052 107332 198116
rect 107396 198052 107397 198116
rect 107331 198051 107397 198052
rect 106779 196756 106845 196757
rect 106779 196692 106780 196756
rect 106844 196692 106845 196756
rect 106779 196691 106845 196692
rect 106782 73949 106842 196691
rect 107147 146980 107213 146981
rect 107147 146916 107148 146980
rect 107212 146916 107213 146980
rect 107147 146915 107213 146916
rect 106779 73948 106845 73949
rect 106779 73884 106780 73948
rect 106844 73884 106845 73948
rect 106779 73883 106845 73884
rect 106043 71092 106109 71093
rect 106043 71028 106044 71092
rect 106108 71028 106109 71092
rect 106043 71027 106109 71028
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 104755 56404 104821 56405
rect 104755 56340 104756 56404
rect 104820 56340 104821 56404
rect 104755 56339 104821 56340
rect 103283 48244 103349 48245
rect 103283 48180 103284 48244
rect 103348 48180 103349 48244
rect 103283 48179 103349 48180
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 34954 105914 70398
rect 107150 52461 107210 146915
rect 107334 78029 107394 198051
rect 107518 78573 107578 198187
rect 108803 191588 108869 191589
rect 108803 191524 108804 191588
rect 108868 191524 108869 191588
rect 108803 191523 108869 191524
rect 108435 148748 108501 148749
rect 108435 148684 108436 148748
rect 108500 148684 108501 148748
rect 108435 148683 108501 148684
rect 108438 84210 108498 148683
rect 108619 147252 108685 147253
rect 108619 147188 108620 147252
rect 108684 147188 108685 147252
rect 108619 147187 108685 147188
rect 108254 84150 108498 84210
rect 108254 80341 108314 84150
rect 108251 80340 108317 80341
rect 108251 80276 108252 80340
rect 108316 80276 108317 80340
rect 108251 80275 108317 80276
rect 107515 78572 107581 78573
rect 107515 78508 107516 78572
rect 107580 78508 107581 78572
rect 107515 78507 107581 78508
rect 107331 78028 107397 78029
rect 107331 77964 107332 78028
rect 107396 77964 107397 78028
rect 107331 77963 107397 77964
rect 108254 65517 108314 80275
rect 108251 65516 108317 65517
rect 108251 65452 108252 65516
rect 108316 65452 108317 65516
rect 108251 65451 108317 65452
rect 107147 52460 107213 52461
rect 107147 52396 107148 52460
rect 107212 52396 107213 52460
rect 107147 52395 107213 52396
rect 107150 51781 107210 52395
rect 107147 51780 107213 51781
rect 107147 51716 107148 51780
rect 107212 51716 107213 51780
rect 107147 51715 107213 51716
rect 108622 45525 108682 147187
rect 108806 58581 108866 191523
rect 109542 146301 109602 262515
rect 109794 255454 110414 290898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 111563 265164 111629 265165
rect 111563 265100 111564 265164
rect 111628 265100 111629 265164
rect 111563 265099 111629 265100
rect 111379 265028 111445 265029
rect 111379 264964 111380 265028
rect 111444 264964 111445 265028
rect 111379 264963 111445 264964
rect 111195 259588 111261 259589
rect 111195 259524 111196 259588
rect 111260 259524 111261 259588
rect 111195 259523 111261 259524
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 110827 147116 110893 147117
rect 110827 147052 110828 147116
rect 110892 147052 110893 147116
rect 110827 147051 110893 147052
rect 109539 146300 109605 146301
rect 109539 146236 109540 146300
rect 109604 146236 109605 146300
rect 109539 146235 109605 146236
rect 109539 140044 109605 140045
rect 109539 139980 109540 140044
rect 109604 139980 109605 140044
rect 109539 139979 109605 139980
rect 108803 58580 108869 58581
rect 108803 58516 108804 58580
rect 108868 58516 108869 58580
rect 108803 58515 108869 58516
rect 109542 54637 109602 139979
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 110830 77213 110890 147051
rect 111011 142764 111077 142765
rect 111011 142700 111012 142764
rect 111076 142700 111077 142764
rect 111011 142699 111077 142700
rect 110827 77212 110893 77213
rect 110827 77148 110828 77212
rect 110892 77148 110893 77212
rect 110827 77147 110893 77148
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109539 54636 109605 54637
rect 109539 54572 109540 54636
rect 109604 54572 109605 54636
rect 109539 54571 109605 54572
rect 108619 45524 108685 45525
rect 108619 45460 108620 45524
rect 108684 45460 108685 45524
rect 108619 45459 108685 45460
rect 108622 44845 108682 45459
rect 108619 44844 108685 44845
rect 108619 44780 108620 44844
rect 108684 44780 108685 44844
rect 108619 44779 108685 44780
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 39454 110414 74898
rect 111014 58037 111074 142699
rect 111198 142629 111258 259523
rect 111382 145621 111442 264963
rect 111566 146029 111626 265099
rect 114139 260268 114205 260269
rect 114139 260204 114140 260268
rect 114204 260204 114205 260268
rect 114139 260203 114205 260204
rect 113035 259996 113101 259997
rect 113035 259932 113036 259996
rect 113100 259932 113101 259996
rect 113035 259931 113101 259932
rect 112851 152420 112917 152421
rect 112851 152356 112852 152420
rect 112916 152356 112917 152420
rect 112851 152355 112917 152356
rect 112667 147660 112733 147661
rect 112667 147596 112668 147660
rect 112732 147596 112733 147660
rect 112667 147595 112733 147596
rect 112483 147388 112549 147389
rect 112483 147324 112484 147388
rect 112548 147324 112549 147388
rect 112483 147323 112549 147324
rect 111563 146028 111629 146029
rect 111563 145964 111564 146028
rect 111628 145964 111629 146028
rect 111563 145963 111629 145964
rect 111379 145620 111445 145621
rect 111379 145556 111380 145620
rect 111444 145556 111445 145620
rect 111379 145555 111445 145556
rect 111195 142628 111261 142629
rect 111195 142564 111196 142628
rect 111260 142564 111261 142628
rect 111195 142563 111261 142564
rect 112486 72725 112546 147323
rect 112670 74629 112730 147595
rect 112667 74628 112733 74629
rect 112667 74564 112668 74628
rect 112732 74564 112733 74628
rect 112667 74563 112733 74564
rect 112483 72724 112549 72725
rect 112483 72660 112484 72724
rect 112548 72660 112549 72724
rect 112483 72659 112549 72660
rect 112854 68781 112914 152355
rect 113038 144805 113098 259931
rect 113955 259724 114021 259725
rect 113955 259660 113956 259724
rect 114020 259660 114021 259724
rect 113955 259659 114021 259660
rect 113958 145893 114018 259659
rect 113955 145892 114021 145893
rect 113955 145828 113956 145892
rect 114020 145828 114021 145892
rect 113955 145827 114021 145828
rect 113035 144804 113101 144805
rect 113035 144740 113036 144804
rect 113100 144740 113101 144804
rect 113035 144739 113101 144740
rect 113955 144124 114021 144125
rect 113955 144060 113956 144124
rect 114020 144060 114021 144124
rect 113955 144059 114021 144060
rect 113771 139772 113837 139773
rect 113771 139708 113772 139772
rect 113836 139708 113837 139772
rect 113771 139707 113837 139708
rect 113587 110532 113653 110533
rect 113587 110468 113588 110532
rect 113652 110468 113653 110532
rect 113587 110467 113653 110468
rect 113590 70141 113650 110467
rect 113774 79389 113834 139707
rect 113958 80477 114018 144059
rect 114142 141405 114202 260203
rect 114294 259954 114914 295398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 115795 263804 115861 263805
rect 115795 263740 115796 263804
rect 115860 263740 115861 263804
rect 115795 263739 115861 263740
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 115611 186964 115677 186965
rect 115611 186900 115612 186964
rect 115676 186900 115677 186964
rect 115611 186899 115677 186900
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114139 141404 114205 141405
rect 114139 141340 114140 141404
rect 114204 141340 114205 141404
rect 114139 141339 114205 141340
rect 114139 139092 114205 139093
rect 114139 139028 114140 139092
rect 114204 139028 114205 139092
rect 114139 139027 114205 139028
rect 113955 80476 114021 80477
rect 113955 80412 113956 80476
rect 114020 80412 114021 80476
rect 113955 80411 114021 80412
rect 113771 79388 113837 79389
rect 113771 79324 113772 79388
rect 113836 79324 113837 79388
rect 113771 79323 113837 79324
rect 113587 70140 113653 70141
rect 113587 70076 113588 70140
rect 113652 70076 113653 70140
rect 113587 70075 113653 70076
rect 114142 68917 114202 139027
rect 114294 115954 114914 151398
rect 115243 144260 115309 144261
rect 115243 144196 115244 144260
rect 115308 144196 115309 144260
rect 115243 144195 115309 144196
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 115246 113797 115306 144195
rect 115243 113796 115309 113797
rect 115243 113732 115244 113796
rect 115308 113732 115309 113796
rect 115243 113731 115309 113732
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114139 68916 114205 68917
rect 114139 68852 114140 68916
rect 114204 68852 114205 68916
rect 114139 68851 114205 68852
rect 112851 68780 112917 68781
rect 112851 68716 112852 68780
rect 112916 68716 112917 68780
rect 112851 68715 112917 68716
rect 111011 58036 111077 58037
rect 111011 57972 111012 58036
rect 111076 57972 111077 58036
rect 111011 57971 111077 57972
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 43954 114914 79398
rect 115614 74901 115674 186899
rect 115798 146165 115858 263739
rect 117083 263668 117149 263669
rect 117083 263604 117084 263668
rect 117148 263604 117149 263668
rect 117083 263603 117149 263604
rect 116899 259860 116965 259861
rect 116899 259796 116900 259860
rect 116964 259796 116965 259860
rect 116899 259795 116965 259796
rect 115795 146164 115861 146165
rect 115795 146100 115796 146164
rect 115860 146100 115861 146164
rect 115795 146099 115861 146100
rect 116347 145756 116413 145757
rect 116347 145692 116348 145756
rect 116412 145692 116413 145756
rect 116347 145691 116413 145692
rect 115611 74900 115677 74901
rect 115611 74836 115612 74900
rect 115676 74836 115677 74900
rect 115611 74835 115677 74836
rect 116350 64701 116410 145691
rect 116902 142901 116962 259795
rect 117086 143037 117146 263603
rect 118794 262000 119414 263898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 262000 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 262000 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 262000 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 262000 137414 281898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 262000 141914 286398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 262000 146414 290898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 262000 150914 295398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 262000 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 262000 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 262000 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 262000 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 262000 173414 281898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 262000 177914 286398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 262000 182414 290898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 262000 186914 295398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 189027 289916 189093 289917
rect 189027 289852 189028 289916
rect 189092 289852 189093 289916
rect 189027 289851 189093 289852
rect 187003 281620 187069 281621
rect 187003 281556 187004 281620
rect 187068 281556 187069 281620
rect 187003 281555 187069 281556
rect 118371 260404 118437 260405
rect 118371 260340 118372 260404
rect 118436 260340 118437 260404
rect 118371 260339 118437 260340
rect 118187 194580 118253 194581
rect 118187 194516 118188 194580
rect 118252 194516 118253 194580
rect 118187 194515 118253 194516
rect 118190 144669 118250 194515
rect 118187 144668 118253 144669
rect 118187 144604 118188 144668
rect 118252 144604 118253 144668
rect 118187 144603 118253 144604
rect 118187 144396 118253 144397
rect 118187 144332 118188 144396
rect 118252 144332 118253 144396
rect 118187 144331 118253 144332
rect 117083 143036 117149 143037
rect 117083 142972 117084 143036
rect 117148 142972 117149 143036
rect 117083 142971 117149 142972
rect 116899 142900 116965 142901
rect 116899 142836 116900 142900
rect 116964 142836 116965 142900
rect 116899 142835 116965 142836
rect 116531 141268 116597 141269
rect 116531 141204 116532 141268
rect 116596 141204 116597 141268
rect 116531 141203 116597 141204
rect 116347 64700 116413 64701
rect 116347 64636 116348 64700
rect 116412 64636 116413 64700
rect 116347 64635 116413 64636
rect 116534 44301 116594 141203
rect 118003 140316 118069 140317
rect 118003 140252 118004 140316
rect 118068 140252 118069 140316
rect 118003 140251 118069 140252
rect 116715 139636 116781 139637
rect 116715 139572 116716 139636
rect 116780 139572 116781 139636
rect 116715 139571 116781 139572
rect 116718 96661 116778 139571
rect 116715 96660 116781 96661
rect 116715 96596 116716 96660
rect 116780 96596 116781 96660
rect 116715 96595 116781 96596
rect 118006 77213 118066 140251
rect 118003 77212 118069 77213
rect 118003 77148 118004 77212
rect 118068 77148 118069 77212
rect 118003 77147 118069 77148
rect 118190 77077 118250 144331
rect 118374 143445 118434 260339
rect 118555 260132 118621 260133
rect 118555 260068 118556 260132
rect 118620 260068 118621 260132
rect 118555 260067 118621 260068
rect 118371 143444 118437 143445
rect 118371 143380 118372 143444
rect 118436 143380 118437 143444
rect 118371 143379 118437 143380
rect 118371 143308 118437 143309
rect 118371 143244 118372 143308
rect 118436 143244 118437 143308
rect 118371 143243 118437 143244
rect 118187 77076 118253 77077
rect 118187 77012 118188 77076
rect 118252 77012 118253 77076
rect 118187 77011 118253 77012
rect 118374 74357 118434 143243
rect 118558 143173 118618 260067
rect 186083 259452 186149 259453
rect 186083 259388 186084 259452
rect 186148 259388 186149 259452
rect 186083 259387 186149 259388
rect 124208 255454 124528 255486
rect 124208 255218 124250 255454
rect 124486 255218 124528 255454
rect 124208 255134 124528 255218
rect 124208 254898 124250 255134
rect 124486 254898 124528 255134
rect 124208 254866 124528 254898
rect 154928 255454 155248 255486
rect 154928 255218 154970 255454
rect 155206 255218 155248 255454
rect 154928 255134 155248 255218
rect 154928 254898 154970 255134
rect 155206 254898 155248 255134
rect 154928 254866 155248 254898
rect 185648 255454 185968 255486
rect 185648 255218 185690 255454
rect 185926 255218 185968 255454
rect 185648 255134 185968 255218
rect 185648 254898 185690 255134
rect 185926 254898 185968 255134
rect 185648 254866 185968 254898
rect 139568 223954 139888 223986
rect 139568 223718 139610 223954
rect 139846 223718 139888 223954
rect 139568 223634 139888 223718
rect 139568 223398 139610 223634
rect 139846 223398 139888 223634
rect 139568 223366 139888 223398
rect 170288 223954 170608 223986
rect 170288 223718 170330 223954
rect 170566 223718 170608 223954
rect 170288 223634 170608 223718
rect 170288 223398 170330 223634
rect 170566 223398 170608 223634
rect 170288 223366 170608 223398
rect 124208 219454 124528 219486
rect 124208 219218 124250 219454
rect 124486 219218 124528 219454
rect 124208 219134 124528 219218
rect 124208 218898 124250 219134
rect 124486 218898 124528 219134
rect 124208 218866 124528 218898
rect 154928 219454 155248 219486
rect 154928 219218 154970 219454
rect 155206 219218 155248 219454
rect 154928 219134 155248 219218
rect 154928 218898 154970 219134
rect 155206 218898 155248 219134
rect 154928 218866 155248 218898
rect 185648 219454 185968 219486
rect 185648 219218 185690 219454
rect 185926 219218 185968 219454
rect 185648 219134 185968 219218
rect 185648 218898 185690 219134
rect 185926 218898 185968 219134
rect 185648 218866 185968 218898
rect 186086 212533 186146 259387
rect 186083 212532 186149 212533
rect 186083 212468 186084 212532
rect 186148 212468 186149 212532
rect 186083 212467 186149 212468
rect 137875 200700 137941 200701
rect 137875 200636 137876 200700
rect 137940 200636 137941 200700
rect 137875 200635 137941 200636
rect 136035 200564 136101 200565
rect 136035 200500 136036 200564
rect 136100 200500 136101 200564
rect 136035 200499 136101 200500
rect 134747 199884 134813 199885
rect 134747 199820 134748 199884
rect 134812 199820 134813 199884
rect 134747 199819 134813 199820
rect 135483 199884 135549 199885
rect 135483 199820 135484 199884
rect 135548 199820 135549 199884
rect 135483 199819 135549 199820
rect 134195 199748 134261 199749
rect 134195 199684 134196 199748
rect 134260 199684 134261 199748
rect 134195 199683 134261 199684
rect 124075 198524 124141 198525
rect 124075 198460 124076 198524
rect 124140 198460 124141 198524
rect 124075 198459 124141 198460
rect 118794 192454 119414 198000
rect 123294 196954 123914 198000
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 122971 194444 123037 194445
rect 122971 194380 122972 194444
rect 123036 194380 123037 194444
rect 122971 194379 123037 194380
rect 122419 194308 122485 194309
rect 122419 194244 122420 194308
rect 122484 194244 122485 194308
rect 122419 194243 122485 194244
rect 119843 192812 119909 192813
rect 119843 192748 119844 192812
rect 119908 192748 119909 192812
rect 119843 192747 119909 192748
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118555 143172 118621 143173
rect 118555 143108 118556 143172
rect 118620 143108 118621 143172
rect 118555 143107 118621 143108
rect 118794 142000 119414 155898
rect 119659 146844 119725 146845
rect 119659 146780 119660 146844
rect 119724 146780 119725 146844
rect 119659 146779 119725 146780
rect 118555 140860 118621 140861
rect 118555 140796 118556 140860
rect 118620 140796 118621 140860
rect 118555 140795 118621 140796
rect 118371 74356 118437 74357
rect 118371 74292 118372 74356
rect 118436 74292 118437 74356
rect 118371 74291 118437 74292
rect 118558 70005 118618 140795
rect 119662 138030 119722 146779
rect 119478 137970 119722 138030
rect 119478 112437 119538 137970
rect 119846 135270 119906 192747
rect 120579 187372 120645 187373
rect 120579 187308 120580 187372
rect 120644 187308 120645 187372
rect 120579 187307 120645 187308
rect 120027 140588 120093 140589
rect 120027 140524 120028 140588
rect 120092 140524 120093 140588
rect 120027 140523 120093 140524
rect 119662 135210 119906 135270
rect 119662 130930 119722 135210
rect 119662 130870 119906 130930
rect 119659 130388 119725 130389
rect 119659 130324 119660 130388
rect 119724 130324 119725 130388
rect 119659 130323 119725 130324
rect 119475 112436 119541 112437
rect 119475 112372 119476 112436
rect 119540 112372 119541 112436
rect 119475 112371 119541 112372
rect 119475 111892 119541 111893
rect 119475 111828 119476 111892
rect 119540 111828 119541 111892
rect 119475 111827 119541 111828
rect 119478 79250 119538 111827
rect 119662 84210 119722 130323
rect 119846 93870 119906 130870
rect 120030 130389 120090 140523
rect 120582 137325 120642 187307
rect 121315 148612 121381 148613
rect 121315 148548 121316 148612
rect 121380 148548 121381 148612
rect 121315 148547 121381 148548
rect 120763 140180 120829 140181
rect 120763 140116 120764 140180
rect 120828 140116 120829 140180
rect 120763 140115 120829 140116
rect 120579 137324 120645 137325
rect 120579 137260 120580 137324
rect 120644 137260 120645 137324
rect 120579 137259 120645 137260
rect 120027 130388 120093 130389
rect 120027 130324 120028 130388
rect 120092 130324 120093 130388
rect 120027 130323 120093 130324
rect 120766 110533 120826 140115
rect 121131 138140 121197 138141
rect 121131 138076 121132 138140
rect 121196 138076 121197 138140
rect 121131 138075 121197 138076
rect 120763 110532 120829 110533
rect 120763 110468 120764 110532
rect 120828 110468 120829 110532
rect 120763 110467 120829 110468
rect 119846 93810 120090 93870
rect 119662 84150 119906 84210
rect 119478 79190 119722 79250
rect 118555 70004 118621 70005
rect 118555 69940 118556 70004
rect 118620 69940 118621 70004
rect 118555 69939 118621 69940
rect 118794 48454 119414 78000
rect 119662 67557 119722 79190
rect 119846 74493 119906 84150
rect 120030 78437 120090 93810
rect 120027 78436 120093 78437
rect 120027 78372 120028 78436
rect 120092 78372 120093 78436
rect 120027 78371 120093 78372
rect 119843 74492 119909 74493
rect 119843 74428 119844 74492
rect 119908 74428 119909 74492
rect 119843 74427 119909 74428
rect 119659 67556 119725 67557
rect 119659 67492 119660 67556
rect 119724 67492 119725 67556
rect 119659 67491 119725 67492
rect 121134 64565 121194 138075
rect 121318 69869 121378 148547
rect 122051 148476 122117 148477
rect 122051 148412 122052 148476
rect 122116 148412 122117 148476
rect 122051 148411 122117 148412
rect 122054 111893 122114 148411
rect 122235 122228 122301 122229
rect 122235 122164 122236 122228
rect 122300 122164 122301 122228
rect 122235 122163 122301 122164
rect 122238 113797 122298 122163
rect 122235 113796 122301 113797
rect 122235 113732 122236 113796
rect 122300 113732 122301 113796
rect 122235 113731 122301 113732
rect 122235 112708 122301 112709
rect 122235 112644 122236 112708
rect 122300 112644 122301 112708
rect 122235 112643 122301 112644
rect 122051 111892 122117 111893
rect 122051 111828 122052 111892
rect 122116 111828 122117 111892
rect 122051 111827 122117 111828
rect 122051 110668 122117 110669
rect 122051 110604 122052 110668
rect 122116 110604 122117 110668
rect 122051 110603 122117 110604
rect 121315 69868 121381 69869
rect 121315 69804 121316 69868
rect 121380 69804 121381 69868
rect 121315 69803 121381 69804
rect 122054 68509 122114 110603
rect 122238 103597 122298 112643
rect 122235 103596 122301 103597
rect 122235 103532 122236 103596
rect 122300 103532 122301 103596
rect 122235 103531 122301 103532
rect 122235 103188 122301 103189
rect 122235 103124 122236 103188
rect 122300 103124 122301 103188
rect 122235 103123 122301 103124
rect 122238 94077 122298 103123
rect 122235 94076 122301 94077
rect 122235 94012 122236 94076
rect 122300 94012 122301 94076
rect 122235 94011 122301 94012
rect 122235 93668 122301 93669
rect 122235 93604 122236 93668
rect 122300 93604 122301 93668
rect 122235 93603 122301 93604
rect 122238 84557 122298 93603
rect 122235 84556 122301 84557
rect 122235 84492 122236 84556
rect 122300 84492 122301 84556
rect 122235 84491 122301 84492
rect 122422 71365 122482 194243
rect 122603 194036 122669 194037
rect 122603 193972 122604 194036
rect 122668 193972 122669 194036
rect 122603 193971 122669 193972
rect 122606 122229 122666 193971
rect 122787 138004 122853 138005
rect 122787 137940 122788 138004
rect 122852 137940 122853 138004
rect 122787 137939 122853 137940
rect 122790 128485 122850 137939
rect 122787 128484 122853 128485
rect 122787 128420 122788 128484
rect 122852 128420 122853 128484
rect 122787 128419 122853 128420
rect 122787 123044 122853 123045
rect 122787 122980 122788 123044
rect 122852 122980 122853 123044
rect 122787 122979 122853 122980
rect 122603 122228 122669 122229
rect 122603 122164 122604 122228
rect 122668 122164 122669 122228
rect 122603 122163 122669 122164
rect 122790 122090 122850 122979
rect 122606 122030 122850 122090
rect 122606 113930 122666 122030
rect 122606 113870 122850 113930
rect 122603 113796 122669 113797
rect 122603 113732 122604 113796
rect 122668 113732 122669 113796
rect 122603 113731 122669 113732
rect 122606 112709 122666 113731
rect 122603 112708 122669 112709
rect 122603 112644 122604 112708
rect 122668 112644 122669 112708
rect 122603 112643 122669 112644
rect 122790 112570 122850 113870
rect 122606 112510 122850 112570
rect 122606 103730 122666 112510
rect 122606 103670 122850 103730
rect 122603 103596 122669 103597
rect 122603 103532 122604 103596
rect 122668 103532 122669 103596
rect 122603 103531 122669 103532
rect 122606 103189 122666 103531
rect 122603 103188 122669 103189
rect 122603 103124 122604 103188
rect 122668 103124 122669 103188
rect 122603 103123 122669 103124
rect 122790 103050 122850 103670
rect 122606 102990 122850 103050
rect 122606 94210 122666 102990
rect 122606 94150 122850 94210
rect 122603 94076 122669 94077
rect 122603 94012 122604 94076
rect 122668 94012 122669 94076
rect 122603 94011 122669 94012
rect 122606 93669 122666 94011
rect 122603 93668 122669 93669
rect 122603 93604 122604 93668
rect 122668 93604 122669 93668
rect 122603 93603 122669 93604
rect 122790 93530 122850 94150
rect 122606 93470 122850 93530
rect 122606 84690 122666 93470
rect 122606 84630 122850 84690
rect 122603 84556 122669 84557
rect 122603 84492 122604 84556
rect 122668 84492 122669 84556
rect 122603 84491 122669 84492
rect 122419 71364 122485 71365
rect 122419 71300 122420 71364
rect 122484 71300 122485 71364
rect 122419 71299 122485 71300
rect 122051 68508 122117 68509
rect 122051 68444 122052 68508
rect 122116 68444 122117 68508
rect 122051 68443 122117 68444
rect 122606 66061 122666 84491
rect 122790 84013 122850 84630
rect 122787 84012 122853 84013
rect 122787 83948 122788 84012
rect 122852 83948 122853 84012
rect 122787 83947 122853 83948
rect 122974 78437 123034 194379
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 142000 123914 160398
rect 123155 138140 123221 138141
rect 123155 138076 123156 138140
rect 123220 138076 123221 138140
rect 123155 138075 123221 138076
rect 123158 123453 123218 138075
rect 123155 123452 123221 123453
rect 123155 123388 123156 123452
rect 123220 123388 123221 123452
rect 123155 123387 123221 123388
rect 124078 81293 124138 198459
rect 134198 197845 134258 199683
rect 134195 197844 134261 197845
rect 134195 197780 134196 197844
rect 134260 197780 134261 197844
rect 134195 197779 134261 197780
rect 134750 196893 134810 199819
rect 135486 197029 135546 199819
rect 136038 199749 136098 200499
rect 136403 199884 136469 199885
rect 136403 199820 136404 199884
rect 136468 199820 136469 199884
rect 136403 199819 136469 199820
rect 136771 199884 136837 199885
rect 136771 199820 136772 199884
rect 136836 199820 136837 199884
rect 136771 199819 136837 199820
rect 136035 199748 136101 199749
rect 136035 199684 136036 199748
rect 136100 199684 136101 199748
rect 136035 199683 136101 199684
rect 136406 198389 136466 199819
rect 136403 198388 136469 198389
rect 136403 198324 136404 198388
rect 136468 198324 136469 198388
rect 136403 198323 136469 198324
rect 135483 197028 135549 197029
rect 135483 196964 135484 197028
rect 135548 196964 135549 197028
rect 135483 196963 135549 196964
rect 134011 196892 134077 196893
rect 134011 196828 134012 196892
rect 134076 196828 134077 196892
rect 134011 196827 134077 196828
rect 134747 196892 134813 196893
rect 134747 196828 134748 196892
rect 134812 196828 134813 196892
rect 134747 196827 134813 196828
rect 135483 196892 135549 196893
rect 135483 196828 135484 196892
rect 135548 196828 135549 196892
rect 135483 196827 135549 196828
rect 134014 191045 134074 196827
rect 134195 196484 134261 196485
rect 134195 196420 134196 196484
rect 134260 196420 134261 196484
rect 134195 196419 134261 196420
rect 134011 191044 134077 191045
rect 134011 190980 134012 191044
rect 134076 190980 134077 191044
rect 134011 190979 134077 190980
rect 124811 189548 124877 189549
rect 124811 189484 124812 189548
rect 124876 189484 124877 189548
rect 124811 189483 124877 189484
rect 124814 137869 124874 189483
rect 134198 151061 134258 196419
rect 135299 195940 135365 195941
rect 135299 195876 135300 195940
rect 135364 195876 135365 195940
rect 135299 195875 135365 195876
rect 134195 151060 134261 151061
rect 134195 150996 134196 151060
rect 134260 150996 134261 151060
rect 134195 150995 134261 150996
rect 135302 148341 135362 195875
rect 135486 187101 135546 196827
rect 136587 196756 136653 196757
rect 136587 196692 136588 196756
rect 136652 196692 136653 196756
rect 136587 196691 136653 196692
rect 135667 196076 135733 196077
rect 135667 196012 135668 196076
rect 135732 196012 135733 196076
rect 135667 196011 135733 196012
rect 135670 187509 135730 196011
rect 135667 187508 135733 187509
rect 135667 187444 135668 187508
rect 135732 187444 135733 187508
rect 135667 187443 135733 187444
rect 135483 187100 135549 187101
rect 135483 187036 135484 187100
rect 135548 187036 135549 187100
rect 135483 187035 135549 187036
rect 135299 148340 135365 148341
rect 135299 148276 135300 148340
rect 135364 148276 135365 148340
rect 135299 148275 135365 148276
rect 136590 146845 136650 196691
rect 136774 151197 136834 199819
rect 137878 199613 137938 200635
rect 171363 200428 171429 200429
rect 171363 200364 171364 200428
rect 171428 200364 171429 200428
rect 171363 200363 171429 200364
rect 138982 200230 139410 200290
rect 138243 199884 138309 199885
rect 138243 199820 138244 199884
rect 138308 199820 138309 199884
rect 138243 199819 138309 199820
rect 138059 199748 138125 199749
rect 138059 199684 138060 199748
rect 138124 199684 138125 199748
rect 138059 199683 138125 199684
rect 137875 199612 137941 199613
rect 137875 199548 137876 199612
rect 137940 199548 137941 199612
rect 137875 199547 137941 199548
rect 136771 151196 136837 151197
rect 136771 151132 136772 151196
rect 136836 151132 136837 151196
rect 136771 151131 136837 151132
rect 138062 146981 138122 199683
rect 138246 187645 138306 199819
rect 138427 198932 138493 198933
rect 138427 198868 138428 198932
rect 138492 198868 138493 198932
rect 138427 198867 138493 198868
rect 138430 191317 138490 198867
rect 138982 197370 139042 200230
rect 139350 200021 139410 200230
rect 166211 200156 166277 200157
rect 166211 200092 166212 200156
rect 166276 200092 166277 200156
rect 166211 200091 166277 200092
rect 139347 200020 139413 200021
rect 139347 199956 139348 200020
rect 139412 199956 139413 200020
rect 139347 199955 139413 199956
rect 141463 199918 141529 199919
rect 139163 199884 139229 199885
rect 139163 199820 139164 199884
rect 139228 199820 139229 199884
rect 139163 199819 139229 199820
rect 140635 199884 140701 199885
rect 140635 199820 140636 199884
rect 140700 199820 140701 199884
rect 141463 199882 141464 199918
rect 140635 199819 140701 199820
rect 140822 199854 141464 199882
rect 141528 199854 141529 199918
rect 140822 199853 141529 199854
rect 141923 199884 141989 199885
rect 140822 199822 141526 199853
rect 139166 198661 139226 199819
rect 139163 198660 139229 198661
rect 139163 198596 139164 198660
rect 139228 198596 139229 198660
rect 139163 198595 139229 198596
rect 138982 197310 139410 197370
rect 138427 191316 138493 191317
rect 138427 191252 138428 191316
rect 138492 191252 138493 191316
rect 138427 191251 138493 191252
rect 138243 187644 138309 187645
rect 138243 187580 138244 187644
rect 138308 187580 138309 187644
rect 138243 187579 138309 187580
rect 139350 147253 139410 197310
rect 140638 196893 140698 199819
rect 139531 196892 139597 196893
rect 139531 196828 139532 196892
rect 139596 196828 139597 196892
rect 139531 196827 139597 196828
rect 140635 196892 140701 196893
rect 140635 196828 140636 196892
rect 140700 196828 140701 196892
rect 140635 196827 140701 196828
rect 139534 153781 139594 196827
rect 139531 153780 139597 153781
rect 139531 153716 139532 153780
rect 139596 153716 139597 153780
rect 139531 153715 139597 153716
rect 140822 148885 140882 199822
rect 141923 199820 141924 199884
rect 141988 199820 141989 199884
rect 141923 199819 141989 199820
rect 142107 199884 142173 199885
rect 142107 199820 142108 199884
rect 142172 199820 142173 199884
rect 142107 199819 142173 199820
rect 142843 199884 142909 199885
rect 142843 199820 142844 199884
rect 142908 199820 142909 199884
rect 142843 199819 142909 199820
rect 143211 199884 143277 199885
rect 143211 199820 143212 199884
rect 143276 199820 143277 199884
rect 143211 199819 143277 199820
rect 144131 199884 144197 199885
rect 144131 199820 144132 199884
rect 144196 199820 144197 199884
rect 144131 199819 144197 199820
rect 145419 199884 145485 199885
rect 145419 199820 145420 199884
rect 145484 199820 145485 199884
rect 146523 199884 146589 199885
rect 146523 199882 146524 199884
rect 145419 199819 145485 199820
rect 146342 199822 146524 199882
rect 141926 198253 141986 199819
rect 141923 198252 141989 198253
rect 141923 198188 141924 198252
rect 141988 198188 141989 198252
rect 141923 198187 141989 198188
rect 141294 178954 141914 198000
rect 142110 197029 142170 199819
rect 142659 199748 142725 199749
rect 142659 199684 142660 199748
rect 142724 199684 142725 199748
rect 142659 199683 142725 199684
rect 142107 197028 142173 197029
rect 142107 196964 142108 197028
rect 142172 196964 142173 197028
rect 142107 196963 142173 196964
rect 142291 196892 142357 196893
rect 142291 196828 142292 196892
rect 142356 196828 142357 196892
rect 142291 196827 142357 196828
rect 142294 190093 142354 196827
rect 142475 196484 142541 196485
rect 142475 196420 142476 196484
rect 142540 196420 142541 196484
rect 142475 196419 142541 196420
rect 142291 190092 142357 190093
rect 142291 190028 142292 190092
rect 142356 190028 142357 190092
rect 142291 190027 142357 190028
rect 142478 189957 142538 196419
rect 142475 189956 142541 189957
rect 142475 189892 142476 189956
rect 142540 189892 142541 189956
rect 142475 189891 142541 189892
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 140819 148884 140885 148885
rect 140819 148820 140820 148884
rect 140884 148820 140885 148884
rect 140819 148819 140885 148820
rect 139347 147252 139413 147253
rect 139347 147188 139348 147252
rect 139412 147188 139413 147252
rect 139347 147187 139413 147188
rect 138059 146980 138125 146981
rect 138059 146916 138060 146980
rect 138124 146916 138125 146980
rect 138059 146915 138125 146916
rect 136587 146844 136653 146845
rect 136587 146780 136588 146844
rect 136652 146780 136653 146844
rect 136587 146779 136653 146780
rect 141294 142954 141914 178398
rect 142662 147525 142722 199683
rect 142846 197437 142906 199819
rect 143214 197437 143274 199819
rect 142843 197436 142909 197437
rect 142843 197372 142844 197436
rect 142908 197372 142909 197436
rect 142843 197371 142909 197372
rect 143211 197436 143277 197437
rect 143211 197372 143212 197436
rect 143276 197372 143277 197436
rect 143211 197371 143277 197372
rect 143763 196756 143829 196757
rect 143763 196692 143764 196756
rect 143828 196692 143829 196756
rect 143763 196691 143829 196692
rect 143579 196076 143645 196077
rect 143579 196012 143580 196076
rect 143644 196012 143645 196076
rect 143579 196011 143645 196012
rect 143582 189685 143642 196011
rect 143766 189821 143826 196691
rect 144134 194445 144194 199819
rect 145051 199748 145117 199749
rect 145051 199684 145052 199748
rect 145116 199684 145117 199748
rect 145051 199683 145117 199684
rect 145054 199205 145114 199683
rect 145422 199205 145482 199819
rect 146342 199205 146402 199822
rect 146523 199820 146524 199822
rect 146588 199820 146589 199884
rect 146523 199819 146589 199820
rect 147259 199884 147325 199885
rect 147259 199820 147260 199884
rect 147324 199820 147325 199884
rect 148179 199884 148245 199885
rect 148179 199882 148180 199884
rect 147259 199819 147325 199820
rect 147998 199822 148180 199882
rect 146523 199748 146589 199749
rect 146523 199684 146524 199748
rect 146588 199684 146589 199748
rect 146523 199683 146589 199684
rect 145051 199204 145117 199205
rect 145051 199140 145052 199204
rect 145116 199140 145117 199204
rect 145051 199139 145117 199140
rect 145419 199204 145485 199205
rect 145419 199140 145420 199204
rect 145484 199140 145485 199204
rect 145419 199139 145485 199140
rect 146339 199204 146405 199205
rect 146339 199140 146340 199204
rect 146404 199140 146405 199204
rect 146339 199139 146405 199140
rect 144315 198932 144381 198933
rect 144315 198868 144316 198932
rect 144380 198868 144381 198932
rect 144315 198867 144381 198868
rect 144318 196077 144378 198867
rect 146526 198661 146586 199683
rect 146523 198660 146589 198661
rect 146523 198596 146524 198660
rect 146588 198596 146589 198660
rect 146523 198595 146589 198596
rect 144315 196076 144381 196077
rect 144315 196012 144316 196076
rect 144380 196012 144381 196076
rect 144315 196011 144381 196012
rect 144131 194444 144197 194445
rect 144131 194380 144132 194444
rect 144196 194380 144197 194444
rect 144131 194379 144197 194380
rect 143763 189820 143829 189821
rect 143763 189756 143764 189820
rect 143828 189756 143829 189820
rect 143763 189755 143829 189756
rect 143579 189684 143645 189685
rect 143579 189620 143580 189684
rect 143644 189620 143645 189684
rect 143579 189619 143645 189620
rect 145794 183454 146414 198000
rect 147262 197029 147322 199819
rect 147627 199748 147693 199749
rect 147627 199684 147628 199748
rect 147692 199684 147693 199748
rect 147627 199683 147693 199684
rect 147811 199748 147877 199749
rect 147811 199684 147812 199748
rect 147876 199684 147877 199748
rect 147811 199683 147877 199684
rect 147443 197980 147509 197981
rect 147443 197916 147444 197980
rect 147508 197916 147509 197980
rect 147443 197915 147509 197916
rect 147259 197028 147325 197029
rect 147259 196964 147260 197028
rect 147324 196964 147325 197028
rect 147259 196963 147325 196964
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 142659 147524 142725 147525
rect 142659 147460 142660 147524
rect 142724 147460 142725 147524
rect 142659 147459 142725 147460
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 142000 141914 142398
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 142000 146414 146898
rect 147446 145621 147506 197915
rect 147630 196485 147690 199683
rect 147627 196484 147693 196485
rect 147627 196420 147628 196484
rect 147692 196420 147693 196484
rect 147627 196419 147693 196420
rect 147814 193221 147874 199683
rect 147811 193220 147877 193221
rect 147811 193156 147812 193220
rect 147876 193156 147877 193220
rect 147811 193155 147877 193156
rect 147998 192677 148058 199822
rect 148179 199820 148180 199822
rect 148244 199820 148245 199884
rect 148179 199819 148245 199820
rect 152779 199884 152845 199885
rect 152779 199820 152780 199884
rect 152844 199820 152845 199884
rect 152779 199819 152845 199820
rect 158299 199884 158365 199885
rect 158299 199820 158300 199884
rect 158364 199820 158365 199884
rect 158299 199819 158365 199820
rect 158667 199884 158733 199885
rect 158667 199820 158668 199884
rect 158732 199820 158733 199884
rect 158667 199819 158733 199820
rect 160875 199884 160941 199885
rect 160875 199820 160876 199884
rect 160940 199820 160941 199884
rect 161243 199884 161309 199885
rect 161243 199882 161244 199884
rect 160875 199819 160941 199820
rect 161062 199822 161244 199882
rect 148915 199748 148981 199749
rect 148915 199684 148916 199748
rect 148980 199684 148981 199748
rect 148915 199683 148981 199684
rect 148179 198116 148245 198117
rect 148179 198052 148180 198116
rect 148244 198052 148245 198116
rect 148179 198051 148245 198052
rect 147995 192676 148061 192677
rect 147995 192612 147996 192676
rect 148060 192612 148061 192676
rect 147995 192611 148061 192612
rect 148182 192541 148242 198051
rect 148918 195669 148978 199683
rect 150019 198524 150085 198525
rect 150019 198460 150020 198524
rect 150084 198460 150085 198524
rect 150019 198459 150085 198460
rect 148915 195668 148981 195669
rect 148915 195604 148916 195668
rect 148980 195604 148981 195668
rect 148915 195603 148981 195604
rect 148179 192540 148245 192541
rect 148179 192476 148180 192540
rect 148244 192476 148245 192540
rect 148179 192475 148245 192476
rect 147627 186420 147693 186421
rect 147627 186356 147628 186420
rect 147692 186356 147693 186420
rect 147627 186355 147693 186356
rect 147443 145620 147509 145621
rect 147443 145556 147444 145620
rect 147508 145556 147509 145620
rect 147443 145555 147509 145556
rect 147630 144533 147690 186355
rect 150022 146981 150082 198459
rect 151491 198388 151557 198389
rect 151491 198324 151492 198388
rect 151556 198324 151557 198388
rect 151491 198323 151557 198324
rect 150294 187954 150914 198000
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150019 146980 150085 146981
rect 150019 146916 150020 146980
rect 150084 146916 150085 146980
rect 150019 146915 150085 146916
rect 147627 144532 147693 144533
rect 147627 144468 147628 144532
rect 147692 144468 147693 144532
rect 147627 144467 147693 144468
rect 150294 142000 150914 151398
rect 130331 140316 130397 140317
rect 130331 140252 130332 140316
rect 130396 140252 130397 140316
rect 130331 140251 130397 140252
rect 130334 139093 130394 140251
rect 151494 140045 151554 198323
rect 152782 194309 152842 199819
rect 157011 199748 157077 199749
rect 157011 199684 157012 199748
rect 157076 199684 157077 199748
rect 157011 199683 157077 199684
rect 154067 195940 154133 195941
rect 154067 195876 154068 195940
rect 154132 195876 154133 195940
rect 154067 195875 154133 195876
rect 152779 194308 152845 194309
rect 152779 194244 152780 194308
rect 152844 194244 152845 194308
rect 152779 194243 152845 194244
rect 154070 155685 154130 195875
rect 154251 193356 154317 193357
rect 154251 193292 154252 193356
rect 154316 193292 154317 193356
rect 154251 193291 154317 193292
rect 154254 189685 154314 193291
rect 154794 192454 155414 198000
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154251 189684 154317 189685
rect 154251 189620 154252 189684
rect 154316 189620 154317 189684
rect 154251 189619 154317 189620
rect 154794 156454 155414 191898
rect 157014 189821 157074 199683
rect 157195 198116 157261 198117
rect 157195 198052 157196 198116
rect 157260 198052 157261 198116
rect 157195 198051 157261 198052
rect 157011 189820 157077 189821
rect 157011 189756 157012 189820
rect 157076 189756 157077 189820
rect 157011 189755 157077 189756
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154067 155684 154133 155685
rect 154067 155620 154068 155684
rect 154132 155620 154133 155684
rect 154067 155619 154133 155620
rect 154794 142000 155414 155898
rect 157198 152693 157258 198051
rect 158302 196077 158362 199819
rect 158299 196076 158365 196077
rect 158299 196012 158300 196076
rect 158364 196012 158365 196076
rect 158299 196011 158365 196012
rect 158670 195669 158730 199819
rect 160691 198660 160757 198661
rect 160691 198596 160692 198660
rect 160756 198596 160757 198660
rect 160691 198595 160757 198596
rect 159294 196954 159914 198000
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 158667 195668 158733 195669
rect 158667 195604 158668 195668
rect 158732 195604 158733 195668
rect 158667 195603 158733 195604
rect 159035 193220 159101 193221
rect 159035 193156 159036 193220
rect 159100 193156 159101 193220
rect 159035 193155 159101 193156
rect 159038 189957 159098 193155
rect 159035 189956 159101 189957
rect 159035 189892 159036 189956
rect 159100 189892 159101 189956
rect 159035 189891 159101 189892
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 157195 152692 157261 152693
rect 157195 152628 157196 152692
rect 157260 152628 157261 152692
rect 157195 152627 157261 152628
rect 159294 142000 159914 160398
rect 160694 151061 160754 198595
rect 160878 196757 160938 199819
rect 161062 197029 161122 199822
rect 161243 199820 161244 199822
rect 161308 199820 161309 199884
rect 161243 199819 161309 199820
rect 162531 199884 162597 199885
rect 162531 199820 162532 199884
rect 162596 199820 162597 199884
rect 162531 199819 162597 199820
rect 164739 199884 164805 199885
rect 164739 199820 164740 199884
rect 164804 199820 164805 199884
rect 164739 199819 164805 199820
rect 165107 199884 165173 199885
rect 165107 199820 165108 199884
rect 165172 199820 165173 199884
rect 165475 199884 165541 199885
rect 165475 199882 165476 199884
rect 165107 199819 165173 199820
rect 165294 199822 165476 199882
rect 161243 199748 161309 199749
rect 161243 199684 161244 199748
rect 161308 199684 161309 199748
rect 161243 199683 161309 199684
rect 161246 197370 161306 199683
rect 161246 197310 161490 197370
rect 161059 197028 161125 197029
rect 161059 196964 161060 197028
rect 161124 196964 161125 197028
rect 161059 196963 161125 196964
rect 161059 196892 161125 196893
rect 161059 196828 161060 196892
rect 161124 196828 161125 196892
rect 161059 196827 161125 196828
rect 160875 196756 160941 196757
rect 160875 196692 160876 196756
rect 160940 196692 160941 196756
rect 160875 196691 160941 196692
rect 161062 152557 161122 196827
rect 161430 195941 161490 197310
rect 161427 195940 161493 195941
rect 161427 195876 161428 195940
rect 161492 195876 161493 195940
rect 161427 195875 161493 195876
rect 162534 191850 162594 199819
rect 163819 199612 163885 199613
rect 163819 199548 163820 199612
rect 163884 199548 163885 199612
rect 163819 199547 163885 199548
rect 162350 191790 162594 191850
rect 162350 191181 162410 191790
rect 162347 191180 162413 191181
rect 162347 191116 162348 191180
rect 162412 191116 162413 191180
rect 162347 191115 162413 191116
rect 161059 152556 161125 152557
rect 161059 152492 161060 152556
rect 161124 152492 161125 152556
rect 161059 152491 161125 152492
rect 160691 151060 160757 151061
rect 160691 150996 160692 151060
rect 160756 150996 160757 151060
rect 160691 150995 160757 150996
rect 163822 148477 163882 199547
rect 164742 197709 164802 199819
rect 164739 197708 164805 197709
rect 164739 197644 164740 197708
rect 164804 197644 164805 197708
rect 164739 197643 164805 197644
rect 165110 197301 165170 199819
rect 165107 197300 165173 197301
rect 165107 197236 165108 197300
rect 165172 197236 165173 197300
rect 165107 197235 165173 197236
rect 165294 191045 165354 199822
rect 165475 199820 165476 199822
rect 165540 199820 165541 199884
rect 165475 199819 165541 199820
rect 165843 199884 165909 199885
rect 165843 199820 165844 199884
rect 165908 199820 165909 199884
rect 165843 199819 165909 199820
rect 165475 199748 165541 199749
rect 165475 199684 165476 199748
rect 165540 199684 165541 199748
rect 165475 199683 165541 199684
rect 165291 191044 165357 191045
rect 165291 190980 165292 191044
rect 165356 190980 165357 191044
rect 165291 190979 165357 190980
rect 165478 155821 165538 199683
rect 165846 196757 165906 199819
rect 166027 199612 166093 199613
rect 166027 199548 166028 199612
rect 166092 199548 166093 199612
rect 166027 199547 166093 199548
rect 165843 196756 165909 196757
rect 165843 196692 165844 196756
rect 165908 196692 165909 196756
rect 165843 196691 165909 196692
rect 166030 196349 166090 199547
rect 166027 196348 166093 196349
rect 166027 196284 166028 196348
rect 166092 196284 166093 196348
rect 166027 196283 166093 196284
rect 165475 155820 165541 155821
rect 165475 155756 165476 155820
rect 165540 155756 165541 155820
rect 165475 155755 165541 155756
rect 163819 148476 163885 148477
rect 163819 148412 163820 148476
rect 163884 148412 163885 148476
rect 163819 148411 163885 148412
rect 166214 147253 166274 200091
rect 166579 199884 166645 199885
rect 166579 199820 166580 199884
rect 166644 199820 166645 199884
rect 166579 199819 166645 199820
rect 168603 199884 168669 199885
rect 168603 199820 168604 199884
rect 168668 199820 168669 199884
rect 168603 199819 168669 199820
rect 169155 199884 169221 199885
rect 169155 199820 169156 199884
rect 169220 199820 169221 199884
rect 169155 199819 169221 199820
rect 169891 199884 169957 199885
rect 169891 199820 169892 199884
rect 169956 199820 169957 199884
rect 169891 199819 169957 199820
rect 170995 199884 171061 199885
rect 170995 199820 170996 199884
rect 171060 199820 171061 199884
rect 170995 199819 171061 199820
rect 166582 151333 166642 199819
rect 168051 199612 168117 199613
rect 168051 199548 168052 199612
rect 168116 199548 168117 199612
rect 168051 199547 168117 199548
rect 167867 198660 167933 198661
rect 167867 198596 167868 198660
rect 167932 198596 167933 198660
rect 167867 198595 167933 198596
rect 167870 186965 167930 198595
rect 168054 197370 168114 199547
rect 168606 199205 168666 199819
rect 168603 199204 168669 199205
rect 168603 199140 168604 199204
rect 168668 199140 168669 199204
rect 168603 199139 168669 199140
rect 169158 198661 169218 199819
rect 169339 199612 169405 199613
rect 169339 199548 169340 199612
rect 169404 199548 169405 199612
rect 169339 199547 169405 199548
rect 169155 198660 169221 198661
rect 169155 198596 169156 198660
rect 169220 198596 169221 198660
rect 169155 198595 169221 198596
rect 168054 197310 168298 197370
rect 168051 195940 168117 195941
rect 168051 195876 168052 195940
rect 168116 195876 168117 195940
rect 168051 195875 168117 195876
rect 167867 186964 167933 186965
rect 167867 186900 167868 186964
rect 167932 186900 167933 186964
rect 167867 186899 167933 186900
rect 168054 158133 168114 195875
rect 168051 158132 168117 158133
rect 168051 158068 168052 158132
rect 168116 158068 168117 158132
rect 168051 158067 168117 158068
rect 168238 155277 168298 197310
rect 169342 155549 169402 199547
rect 169523 198660 169589 198661
rect 169523 198596 169524 198660
rect 169588 198596 169589 198660
rect 169523 198595 169589 198596
rect 169339 155548 169405 155549
rect 169339 155484 169340 155548
rect 169404 155484 169405 155548
rect 169339 155483 169405 155484
rect 168235 155276 168301 155277
rect 168235 155212 168236 155276
rect 168300 155212 168301 155276
rect 168235 155211 168301 155212
rect 166579 151332 166645 151333
rect 166579 151268 166580 151332
rect 166644 151268 166645 151332
rect 166579 151267 166645 151268
rect 169526 148341 169586 198595
rect 169894 196485 169954 199819
rect 169891 196484 169957 196485
rect 169891 196420 169892 196484
rect 169956 196420 169957 196484
rect 169891 196419 169957 196420
rect 170998 196077 171058 199819
rect 171366 199477 171426 200363
rect 171915 199884 171981 199885
rect 171915 199820 171916 199884
rect 171980 199820 171981 199884
rect 171915 199819 171981 199820
rect 172651 199884 172717 199885
rect 172651 199820 172652 199884
rect 172716 199820 172717 199884
rect 172651 199819 172717 199820
rect 173571 199884 173637 199885
rect 173571 199820 173572 199884
rect 173636 199820 173637 199884
rect 173571 199819 173637 199820
rect 174859 199884 174925 199885
rect 174859 199820 174860 199884
rect 174924 199820 174925 199884
rect 174859 199819 174925 199820
rect 176331 199884 176397 199885
rect 176331 199820 176332 199884
rect 176396 199820 176397 199884
rect 176331 199819 176397 199820
rect 171547 199612 171613 199613
rect 171547 199548 171548 199612
rect 171612 199548 171613 199612
rect 171547 199547 171613 199548
rect 171363 199476 171429 199477
rect 171363 199412 171364 199476
rect 171428 199412 171429 199476
rect 171363 199411 171429 199412
rect 171550 197981 171610 199547
rect 171918 198525 171978 199819
rect 171915 198524 171981 198525
rect 171915 198460 171916 198524
rect 171980 198460 171981 198524
rect 171915 198459 171981 198460
rect 171547 197980 171613 197981
rect 171547 197916 171548 197980
rect 171612 197916 171613 197980
rect 171547 197915 171613 197916
rect 170995 196076 171061 196077
rect 170995 196012 170996 196076
rect 171060 196012 171061 196076
rect 170995 196011 171061 196012
rect 170995 195940 171061 195941
rect 170995 195876 170996 195940
rect 171060 195876 171061 195940
rect 170995 195875 171061 195876
rect 169523 148340 169589 148341
rect 169523 148276 169524 148340
rect 169588 148276 169589 148340
rect 169523 148275 169589 148276
rect 166211 147252 166277 147253
rect 166211 147188 166212 147252
rect 166276 147188 166277 147252
rect 166211 147187 166277 147188
rect 170998 147117 171058 195875
rect 172654 194309 172714 199819
rect 173574 198389 173634 199819
rect 173755 199748 173821 199749
rect 173755 199684 173756 199748
rect 173820 199684 173821 199748
rect 173755 199683 173821 199684
rect 173758 199205 173818 199683
rect 173755 199204 173821 199205
rect 173755 199140 173756 199204
rect 173820 199140 173821 199204
rect 173755 199139 173821 199140
rect 173571 198388 173637 198389
rect 173571 198324 173572 198388
rect 173636 198324 173637 198388
rect 173571 198323 173637 198324
rect 172651 194308 172717 194309
rect 172651 194244 172652 194308
rect 172716 194244 172717 194308
rect 172651 194243 172717 194244
rect 174862 191850 174922 199819
rect 174678 191790 174922 191850
rect 174678 190093 174738 191790
rect 176334 190229 176394 199819
rect 176331 190228 176397 190229
rect 176331 190164 176332 190228
rect 176396 190164 176397 190228
rect 176331 190163 176397 190164
rect 174675 190092 174741 190093
rect 174675 190028 174676 190092
rect 174740 190028 174741 190092
rect 174675 190027 174741 190028
rect 177294 178954 177914 198000
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 170995 147116 171061 147117
rect 170995 147052 170996 147116
rect 171060 147052 171061 147116
rect 170995 147051 171061 147052
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 142000 177914 142398
rect 181794 183454 182414 198000
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 142000 182414 146898
rect 186294 187954 186914 198000
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 142000 186914 151398
rect 187006 144125 187066 281555
rect 187739 192948 187805 192949
rect 187739 192884 187740 192948
rect 187804 192884 187805 192948
rect 187739 192883 187805 192884
rect 187187 187100 187253 187101
rect 187187 187036 187188 187100
rect 187252 187036 187253 187100
rect 187187 187035 187253 187036
rect 187003 144124 187069 144125
rect 187003 144060 187004 144124
rect 187068 144060 187069 144124
rect 187003 144059 187069 144060
rect 151491 140044 151557 140045
rect 151491 139980 151492 140044
rect 151556 139980 151557 140044
rect 151491 139979 151557 139980
rect 130331 139092 130397 139093
rect 130331 139028 130332 139092
rect 130396 139028 130397 139092
rect 130331 139027 130397 139028
rect 187190 137869 187250 187035
rect 124811 137868 124877 137869
rect 124811 137804 124812 137868
rect 124876 137804 124877 137868
rect 124811 137803 124877 137804
rect 187187 137868 187253 137869
rect 187187 137804 187188 137868
rect 187252 137804 187253 137868
rect 187187 137803 187253 137804
rect 139568 115954 139888 115986
rect 139568 115718 139610 115954
rect 139846 115718 139888 115954
rect 139568 115634 139888 115718
rect 139568 115398 139610 115634
rect 139846 115398 139888 115634
rect 139568 115366 139888 115398
rect 170288 115954 170608 115986
rect 170288 115718 170330 115954
rect 170566 115718 170608 115954
rect 170288 115634 170608 115718
rect 170288 115398 170330 115634
rect 170566 115398 170608 115634
rect 170288 115366 170608 115398
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 185648 111454 185968 111486
rect 185648 111218 185690 111454
rect 185926 111218 185968 111454
rect 185648 111134 185968 111218
rect 185648 110898 185690 111134
rect 185926 110898 185968 111134
rect 185648 110866 185968 110898
rect 187742 109850 187802 192883
rect 187923 147660 187989 147661
rect 187923 147596 187924 147660
rect 187988 147596 187989 147660
rect 187923 147595 187989 147596
rect 187926 138005 187986 147595
rect 189030 144397 189090 289851
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 262000 191414 263898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 193443 262580 193509 262581
rect 193443 262516 193444 262580
rect 193508 262516 193509 262580
rect 193443 262515 193509 262516
rect 193259 262444 193325 262445
rect 193259 262380 193260 262444
rect 193324 262380 193325 262444
rect 193259 262379 193325 262380
rect 190794 192454 191414 198000
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 189211 146028 189277 146029
rect 189211 145964 189212 146028
rect 189276 145964 189277 146028
rect 189211 145963 189277 145964
rect 189027 144396 189093 144397
rect 189027 144332 189028 144396
rect 189092 144332 189093 144396
rect 189027 144331 189093 144332
rect 188291 140452 188357 140453
rect 188291 140388 188292 140452
rect 188356 140388 188357 140452
rect 188291 140387 188357 140388
rect 187923 138004 187989 138005
rect 187923 137940 187924 138004
rect 187988 137940 187989 138004
rect 187923 137939 187989 137940
rect 188294 137869 188354 140387
rect 188291 137868 188357 137869
rect 188291 137804 188292 137868
rect 188356 137804 188357 137868
rect 188291 137803 188357 137804
rect 189214 115950 189274 145963
rect 189763 144804 189829 144805
rect 189763 144740 189764 144804
rect 189828 144740 189829 144804
rect 189763 144739 189829 144740
rect 189579 141540 189645 141541
rect 189579 141476 189580 141540
rect 189644 141476 189645 141540
rect 189579 141475 189645 141476
rect 189395 139500 189461 139501
rect 189395 139436 189396 139500
rect 189460 139436 189461 139500
rect 189395 139435 189461 139436
rect 188478 115890 189274 115950
rect 188478 113190 188538 115890
rect 189398 113389 189458 139435
rect 189582 113933 189642 141475
rect 189579 113932 189645 113933
rect 189579 113868 189580 113932
rect 189644 113868 189645 113932
rect 189579 113867 189645 113868
rect 189395 113388 189461 113389
rect 189395 113324 189396 113388
rect 189460 113324 189461 113388
rect 189395 113323 189461 113324
rect 189579 113388 189645 113389
rect 189579 113324 189580 113388
rect 189644 113324 189645 113388
rect 189579 113323 189645 113324
rect 188478 113130 189458 113190
rect 189398 110669 189458 113130
rect 189395 110668 189461 110669
rect 189395 110604 189396 110668
rect 189460 110604 189461 110668
rect 189395 110603 189461 110604
rect 188478 110470 189458 110530
rect 188478 109850 188538 110470
rect 187742 109790 188538 109850
rect 189398 109309 189458 110470
rect 189395 109308 189461 109309
rect 189395 109244 189396 109308
rect 189460 109244 189461 109308
rect 189395 109243 189461 109244
rect 189395 107132 189461 107133
rect 189395 107130 189396 107132
rect 189214 107070 189396 107130
rect 124075 81292 124141 81293
rect 124075 81228 124076 81292
rect 124140 81228 124141 81292
rect 124075 81227 124141 81228
rect 147811 81292 147877 81293
rect 147811 81228 147812 81292
rect 147876 81228 147877 81292
rect 147811 81227 147877 81228
rect 164003 81292 164069 81293
rect 164003 81228 164004 81292
rect 164068 81228 164069 81292
rect 164003 81227 164069 81228
rect 146339 80748 146405 80749
rect 146339 80684 146340 80748
rect 146404 80684 146405 80748
rect 146339 80683 146405 80684
rect 139347 80204 139413 80205
rect 139347 80140 139348 80204
rect 139412 80140 139413 80204
rect 139347 80139 139413 80140
rect 143395 80204 143461 80205
rect 143395 80140 143396 80204
rect 143460 80140 143461 80204
rect 143395 80139 143461 80140
rect 135299 80068 135365 80069
rect 135299 80004 135300 80068
rect 135364 80004 135365 80068
rect 135299 80003 135365 80004
rect 134195 79932 134261 79933
rect 134195 79868 134196 79932
rect 134260 79868 134261 79932
rect 134195 79867 134261 79868
rect 134563 79932 134629 79933
rect 134563 79868 134564 79932
rect 134628 79868 134629 79932
rect 134563 79867 134629 79868
rect 122971 78436 123037 78437
rect 122971 78372 122972 78436
rect 123036 78372 123037 78436
rect 122971 78371 123037 78372
rect 134011 78028 134077 78029
rect 122603 66060 122669 66061
rect 122603 65996 122604 66060
rect 122668 65996 122669 66060
rect 122603 65995 122669 65996
rect 121131 64564 121197 64565
rect 121131 64500 121132 64564
rect 121196 64500 121197 64564
rect 121131 64499 121197 64500
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 116531 44300 116597 44301
rect 116531 44236 116532 44300
rect 116596 44236 116597 44300
rect 116531 44235 116597 44236
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 78000
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 78000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 78000
rect 134011 77964 134012 78028
rect 134076 77964 134077 78028
rect 134011 77963 134077 77964
rect 133459 77620 133525 77621
rect 133459 77556 133460 77620
rect 133524 77556 133525 77620
rect 133459 77555 133525 77556
rect 133275 77484 133341 77485
rect 133275 77420 133276 77484
rect 133340 77420 133341 77484
rect 133275 77419 133341 77420
rect 133091 77348 133157 77349
rect 133091 77284 133092 77348
rect 133156 77284 133157 77348
rect 133091 77283 133157 77284
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 133094 53685 133154 77283
rect 133278 56541 133338 77419
rect 133462 67421 133522 77555
rect 133827 76668 133893 76669
rect 133827 76604 133828 76668
rect 133892 76604 133893 76668
rect 133827 76603 133893 76604
rect 133459 67420 133525 67421
rect 133459 67356 133460 67420
rect 133524 67356 133525 67420
rect 133459 67355 133525 67356
rect 133275 56540 133341 56541
rect 133275 56476 133276 56540
rect 133340 56476 133341 56540
rect 133275 56475 133341 56476
rect 133091 53684 133157 53685
rect 133091 53620 133092 53684
rect 133156 53620 133157 53684
rect 133091 53619 133157 53620
rect 133830 50965 133890 76603
rect 134014 57765 134074 77963
rect 134198 62117 134258 79867
rect 134566 77349 134626 79867
rect 134563 77348 134629 77349
rect 134563 77284 134564 77348
rect 134628 77284 134629 77348
rect 134563 77283 134629 77284
rect 134195 62116 134261 62117
rect 134195 62052 134196 62116
rect 134260 62052 134261 62116
rect 134195 62051 134261 62052
rect 134011 57764 134077 57765
rect 134011 57700 134012 57764
rect 134076 57700 134077 57764
rect 134011 57699 134077 57700
rect 133827 50964 133893 50965
rect 133827 50900 133828 50964
rect 133892 50900 133893 50964
rect 133827 50899 133893 50900
rect 135302 46885 135362 80003
rect 135851 79932 135917 79933
rect 135851 79868 135852 79932
rect 135916 79868 135917 79932
rect 135851 79867 135917 79868
rect 136955 79932 137021 79933
rect 136955 79868 136956 79932
rect 137020 79868 137021 79932
rect 136955 79867 137021 79868
rect 137875 79932 137941 79933
rect 137875 79868 137876 79932
rect 137940 79868 137941 79932
rect 137875 79867 137941 79868
rect 138611 79932 138677 79933
rect 138611 79868 138612 79932
rect 138676 79868 138677 79932
rect 138611 79867 138677 79868
rect 138979 79932 139045 79933
rect 138979 79868 138980 79932
rect 139044 79868 139045 79932
rect 138979 79867 139045 79868
rect 135667 79796 135733 79797
rect 135667 79732 135668 79796
rect 135732 79732 135733 79796
rect 135667 79731 135733 79732
rect 135483 77484 135549 77485
rect 135483 77420 135484 77484
rect 135548 77420 135549 77484
rect 135483 77419 135549 77420
rect 135486 48245 135546 77419
rect 135670 49605 135730 79731
rect 135854 55181 135914 79867
rect 136587 79388 136653 79389
rect 136587 79324 136588 79388
rect 136652 79324 136653 79388
rect 136587 79323 136653 79324
rect 135851 55180 135917 55181
rect 135851 55116 135852 55180
rect 135916 55116 135917 55180
rect 135851 55115 135917 55116
rect 135667 49604 135733 49605
rect 135667 49540 135668 49604
rect 135732 49540 135733 49604
rect 135667 49539 135733 49540
rect 135483 48244 135549 48245
rect 135483 48180 135484 48244
rect 135548 48180 135549 48244
rect 135483 48179 135549 48180
rect 135299 46884 135365 46885
rect 135299 46820 135300 46884
rect 135364 46820 135365 46884
rect 135299 46819 135365 46820
rect 136590 44165 136650 79323
rect 136958 78165 137018 79867
rect 137878 78709 137938 79867
rect 137875 78708 137941 78709
rect 137875 78644 137876 78708
rect 137940 78644 137941 78708
rect 137875 78643 137941 78644
rect 137507 78300 137573 78301
rect 137507 78236 137508 78300
rect 137572 78236 137573 78300
rect 137507 78235 137573 78236
rect 136955 78164 137021 78165
rect 136955 78100 136956 78164
rect 137020 78100 137021 78164
rect 136955 78099 137021 78100
rect 136794 66454 137414 78000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136587 44164 136653 44165
rect 136587 44100 136588 44164
rect 136652 44100 136653 44164
rect 136587 44099 136653 44100
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 30454 137414 65898
rect 137510 56405 137570 78235
rect 138059 76124 138125 76125
rect 138059 76060 138060 76124
rect 138124 76060 138125 76124
rect 138059 76059 138125 76060
rect 138243 76124 138309 76125
rect 138243 76060 138244 76124
rect 138308 76060 138309 76124
rect 138243 76059 138309 76060
rect 137507 56404 137573 56405
rect 137507 56340 137508 56404
rect 137572 56340 137573 56404
rect 137507 56339 137573 56340
rect 138062 41309 138122 76059
rect 138246 52461 138306 76059
rect 138614 75986 138674 79867
rect 138430 75926 138674 75986
rect 138430 57901 138490 75926
rect 138982 75853 139042 79867
rect 138979 75852 139045 75853
rect 138979 75788 138980 75852
rect 139044 75788 139045 75852
rect 138979 75787 139045 75788
rect 138611 75172 138677 75173
rect 138611 75108 138612 75172
rect 138676 75108 138677 75172
rect 138611 75107 138677 75108
rect 138614 61981 138674 75107
rect 138611 61980 138677 61981
rect 138611 61916 138612 61980
rect 138676 61916 138677 61980
rect 138611 61915 138677 61916
rect 138427 57900 138493 57901
rect 138427 57836 138428 57900
rect 138492 57836 138493 57900
rect 138427 57835 138493 57836
rect 138243 52460 138309 52461
rect 138243 52396 138244 52460
rect 138308 52396 138309 52460
rect 138243 52395 138309 52396
rect 138059 41308 138125 41309
rect 138059 41244 138060 41308
rect 138124 41244 138125 41308
rect 138059 41243 138125 41244
rect 139350 36549 139410 80139
rect 139715 79932 139781 79933
rect 139715 79868 139716 79932
rect 139780 79868 139781 79932
rect 139715 79867 139781 79868
rect 139899 79932 139965 79933
rect 139899 79868 139900 79932
rect 139964 79868 139965 79932
rect 139899 79867 139965 79868
rect 140635 79932 140701 79933
rect 140635 79868 140636 79932
rect 140700 79868 140701 79932
rect 141187 79932 141253 79933
rect 141187 79930 141188 79932
rect 140635 79867 140701 79868
rect 141006 79870 141188 79930
rect 139531 78300 139597 78301
rect 139531 78236 139532 78300
rect 139596 78236 139597 78300
rect 139531 78235 139597 78236
rect 139534 45525 139594 78235
rect 139718 53821 139778 79867
rect 139902 79389 139962 79867
rect 139899 79388 139965 79389
rect 139899 79324 139900 79388
rect 139964 79324 139965 79388
rect 139899 79323 139965 79324
rect 140638 78709 140698 79867
rect 140819 79524 140885 79525
rect 140819 79460 140820 79524
rect 140884 79460 140885 79524
rect 140819 79459 140885 79460
rect 140635 78708 140701 78709
rect 140635 78644 140636 78708
rect 140700 78644 140701 78708
rect 140635 78643 140701 78644
rect 139899 78028 139965 78029
rect 139899 77964 139900 78028
rect 139964 77964 139965 78028
rect 139899 77963 139965 77964
rect 139902 59261 139962 77963
rect 140822 77310 140882 79459
rect 140638 77250 140882 77310
rect 140638 76261 140698 77250
rect 140635 76260 140701 76261
rect 140635 76196 140636 76260
rect 140700 76196 140701 76260
rect 140635 76195 140701 76196
rect 140819 75172 140885 75173
rect 140819 75108 140820 75172
rect 140884 75108 140885 75172
rect 140819 75107 140885 75108
rect 140822 61845 140882 75107
rect 141006 65517 141066 79870
rect 141187 79868 141188 79870
rect 141252 79868 141253 79932
rect 141187 79867 141253 79868
rect 142291 79932 142357 79933
rect 142291 79868 142292 79932
rect 142356 79868 142357 79932
rect 142291 79867 142357 79868
rect 142659 79932 142725 79933
rect 142659 79868 142660 79932
rect 142724 79868 142725 79932
rect 143027 79932 143093 79933
rect 143027 79930 143028 79932
rect 142659 79867 142725 79868
rect 142846 79870 143028 79930
rect 142294 78301 142354 79867
rect 142662 79525 142722 79867
rect 142659 79524 142725 79525
rect 142659 79460 142660 79524
rect 142724 79460 142725 79524
rect 142659 79459 142725 79460
rect 142291 78300 142357 78301
rect 142291 78236 142292 78300
rect 142356 78236 142357 78300
rect 142291 78235 142357 78236
rect 141294 70954 141914 78000
rect 142846 77349 142906 79870
rect 143027 79868 143028 79870
rect 143092 79868 143093 79932
rect 143027 79867 143093 79868
rect 143211 79932 143277 79933
rect 143211 79868 143212 79932
rect 143276 79868 143277 79932
rect 143211 79867 143277 79868
rect 143027 79660 143093 79661
rect 143027 79596 143028 79660
rect 143092 79596 143093 79660
rect 143027 79595 143093 79596
rect 142843 77348 142909 77349
rect 142843 77284 142844 77348
rect 142908 77284 142909 77348
rect 142843 77283 142909 77284
rect 143030 73813 143090 79595
rect 143214 77349 143274 79867
rect 143398 79525 143458 80139
rect 143763 79932 143829 79933
rect 143763 79868 143764 79932
rect 143828 79868 143829 79932
rect 143763 79867 143829 79868
rect 144315 79932 144381 79933
rect 144315 79868 144316 79932
rect 144380 79868 144381 79932
rect 144315 79867 144381 79868
rect 144683 79932 144749 79933
rect 144683 79868 144684 79932
rect 144748 79868 144749 79932
rect 144683 79867 144749 79868
rect 145051 79932 145117 79933
rect 145051 79868 145052 79932
rect 145116 79868 145117 79932
rect 145051 79867 145117 79868
rect 145419 79932 145485 79933
rect 145419 79868 145420 79932
rect 145484 79868 145485 79932
rect 145419 79867 145485 79868
rect 145603 79932 145669 79933
rect 145603 79868 145604 79932
rect 145668 79868 145669 79932
rect 145603 79867 145669 79868
rect 143395 79524 143461 79525
rect 143395 79460 143396 79524
rect 143460 79460 143461 79524
rect 143395 79459 143461 79460
rect 143579 77484 143645 77485
rect 143579 77420 143580 77484
rect 143644 77420 143645 77484
rect 143579 77419 143645 77420
rect 143211 77348 143277 77349
rect 143211 77284 143212 77348
rect 143276 77284 143277 77348
rect 143211 77283 143277 77284
rect 143027 73812 143093 73813
rect 143027 73748 143028 73812
rect 143092 73748 143093 73812
rect 143027 73747 143093 73748
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141003 65516 141069 65517
rect 141003 65452 141004 65516
rect 141068 65452 141069 65516
rect 141003 65451 141069 65452
rect 140819 61844 140885 61845
rect 140819 61780 140820 61844
rect 140884 61780 140885 61844
rect 140819 61779 140885 61780
rect 139899 59260 139965 59261
rect 139899 59196 139900 59260
rect 139964 59196 139965 59260
rect 139899 59195 139965 59196
rect 139715 53820 139781 53821
rect 139715 53756 139716 53820
rect 139780 53756 139781 53820
rect 139715 53755 139781 53756
rect 139531 45524 139597 45525
rect 139531 45460 139532 45524
rect 139596 45460 139597 45524
rect 139531 45459 139597 45460
rect 139347 36548 139413 36549
rect 139347 36484 139348 36548
rect 139412 36484 139413 36548
rect 139347 36483 139413 36484
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 34954 141914 70398
rect 143582 64837 143642 77419
rect 143766 77077 143826 79867
rect 144131 77620 144197 77621
rect 144131 77556 144132 77620
rect 144196 77556 144197 77620
rect 144131 77555 144197 77556
rect 143763 77076 143829 77077
rect 143763 77012 143764 77076
rect 143828 77012 143829 77076
rect 143763 77011 143829 77012
rect 143763 76940 143829 76941
rect 143763 76876 143764 76940
rect 143828 76876 143829 76940
rect 143763 76875 143829 76876
rect 143766 65925 143826 76875
rect 144134 70410 144194 77555
rect 144318 77349 144378 79867
rect 144686 79525 144746 79867
rect 145054 79525 145114 79867
rect 144683 79524 144749 79525
rect 144683 79460 144684 79524
rect 144748 79460 144749 79524
rect 144683 79459 144749 79460
rect 145051 79524 145117 79525
rect 145051 79460 145052 79524
rect 145116 79460 145117 79524
rect 145051 79459 145117 79460
rect 145422 78709 145482 79867
rect 145419 78708 145485 78709
rect 145419 78644 145420 78708
rect 145484 78644 145485 78708
rect 145419 78643 145485 78644
rect 144315 77348 144381 77349
rect 144315 77284 144316 77348
rect 144380 77284 144381 77348
rect 144315 77283 144381 77284
rect 145606 76261 145666 79867
rect 146342 79661 146402 80683
rect 147075 80204 147141 80205
rect 147075 80140 147076 80204
rect 147140 80140 147141 80204
rect 147075 80139 147141 80140
rect 146523 79932 146589 79933
rect 146523 79868 146524 79932
rect 146588 79868 146589 79932
rect 146523 79867 146589 79868
rect 146339 79660 146405 79661
rect 146339 79596 146340 79660
rect 146404 79596 146405 79660
rect 146339 79595 146405 79596
rect 145603 76260 145669 76261
rect 145603 76196 145604 76260
rect 145668 76196 145669 76260
rect 145603 76195 145669 76196
rect 145419 75580 145485 75581
rect 145419 75516 145420 75580
rect 145484 75516 145485 75580
rect 145419 75515 145485 75516
rect 145422 75173 145482 75515
rect 145794 75454 146414 78000
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145419 75172 145485 75173
rect 145419 75108 145420 75172
rect 145484 75108 145485 75172
rect 145419 75107 145485 75108
rect 145794 75134 146414 75218
rect 144315 75036 144381 75037
rect 144315 74972 144316 75036
rect 144380 74972 144381 75036
rect 144315 74971 144381 74972
rect 143950 70350 144194 70410
rect 143950 66197 144010 70350
rect 144318 70277 144378 74971
rect 144315 70276 144381 70277
rect 144315 70212 144316 70276
rect 144380 70212 144381 70276
rect 144315 70211 144381 70212
rect 143947 66196 144013 66197
rect 143947 66132 143948 66196
rect 144012 66132 144013 66196
rect 143947 66131 144013 66132
rect 143763 65924 143829 65925
rect 143763 65860 143764 65924
rect 143828 65860 143829 65924
rect 143763 65859 143829 65860
rect 143579 64836 143645 64837
rect 143579 64772 143580 64836
rect 143644 64772 143645 64836
rect 143579 64771 143645 64772
rect 143582 63613 143642 64771
rect 143579 63612 143645 63613
rect 143579 63548 143580 63612
rect 143644 63548 143645 63612
rect 143579 63547 143645 63548
rect 143766 55230 143826 65859
rect 143766 55170 144194 55230
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 144134 7581 144194 55170
rect 144318 15877 144378 70211
rect 144683 66196 144749 66197
rect 144683 66132 144684 66196
rect 144748 66132 144749 66196
rect 144683 66131 144749 66132
rect 144499 63612 144565 63613
rect 144499 63548 144500 63612
rect 144564 63548 144565 63612
rect 144499 63547 144565 63548
rect 144502 46205 144562 63547
rect 144686 56541 144746 66131
rect 144683 56540 144749 56541
rect 144683 56476 144684 56540
rect 144748 56476 144749 56540
rect 144683 56475 144749 56476
rect 144499 46204 144565 46205
rect 144499 46140 144500 46204
rect 144564 46140 144565 46204
rect 144499 46139 144565 46140
rect 145422 22677 145482 75107
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 146526 68781 146586 79867
rect 146891 79252 146957 79253
rect 146891 79188 146892 79252
rect 146956 79188 146957 79252
rect 146891 79187 146957 79188
rect 146894 76261 146954 79187
rect 146891 76260 146957 76261
rect 146891 76196 146892 76260
rect 146956 76196 146957 76260
rect 146891 76195 146957 76196
rect 147078 71773 147138 80139
rect 147627 79932 147693 79933
rect 147627 79868 147628 79932
rect 147692 79868 147693 79932
rect 147627 79867 147693 79868
rect 147259 79660 147325 79661
rect 147259 79596 147260 79660
rect 147324 79596 147325 79660
rect 147259 79595 147325 79596
rect 147262 75717 147322 79595
rect 147630 79253 147690 79867
rect 147814 79661 147874 81227
rect 151307 81020 151373 81021
rect 151307 80956 151308 81020
rect 151372 80956 151373 81020
rect 151307 80955 151373 80956
rect 148915 80884 148981 80885
rect 148915 80820 148916 80884
rect 148980 80820 148981 80884
rect 148915 80819 148981 80820
rect 147995 79932 148061 79933
rect 147995 79868 147996 79932
rect 148060 79868 148061 79932
rect 147995 79867 148061 79868
rect 148363 79932 148429 79933
rect 148363 79868 148364 79932
rect 148428 79868 148429 79932
rect 148363 79867 148429 79868
rect 147811 79660 147877 79661
rect 147811 79596 147812 79660
rect 147876 79596 147877 79660
rect 147811 79595 147877 79596
rect 147811 79524 147877 79525
rect 147811 79460 147812 79524
rect 147876 79460 147877 79524
rect 147811 79459 147877 79460
rect 147627 79252 147693 79253
rect 147627 79188 147628 79252
rect 147692 79188 147693 79252
rect 147627 79187 147693 79188
rect 147259 75716 147325 75717
rect 147259 75652 147260 75716
rect 147324 75652 147325 75716
rect 147259 75651 147325 75652
rect 147075 71772 147141 71773
rect 147075 71708 147076 71772
rect 147140 71708 147141 71772
rect 147075 71707 147141 71708
rect 146523 68780 146589 68781
rect 146523 68716 146524 68780
rect 146588 68716 146589 68780
rect 146523 68715 146589 68716
rect 146526 64890 146586 68715
rect 146526 64830 146954 64890
rect 146894 43485 146954 64830
rect 147078 50285 147138 71707
rect 147262 65517 147322 75651
rect 147814 68509 147874 79459
rect 147998 77485 148058 79867
rect 147995 77484 148061 77485
rect 147995 77420 147996 77484
rect 148060 77420 148061 77484
rect 147995 77419 148061 77420
rect 148179 77484 148245 77485
rect 148179 77420 148180 77484
rect 148244 77420 148245 77484
rect 148179 77419 148245 77420
rect 147995 77348 148061 77349
rect 147995 77284 147996 77348
rect 148060 77284 148061 77348
rect 147995 77283 148061 77284
rect 147998 68917 148058 77283
rect 148182 71229 148242 77419
rect 148366 72725 148426 79867
rect 148918 79661 148978 80819
rect 151310 79933 151370 80955
rect 158115 80204 158181 80205
rect 158115 80140 158116 80204
rect 158180 80140 158181 80204
rect 158115 80139 158181 80140
rect 151675 80068 151741 80069
rect 151675 80004 151676 80068
rect 151740 80004 151741 80068
rect 151675 80003 151741 80004
rect 149467 79932 149533 79933
rect 149467 79868 149468 79932
rect 149532 79868 149533 79932
rect 149467 79867 149533 79868
rect 149651 79932 149717 79933
rect 149651 79868 149652 79932
rect 149716 79868 149717 79932
rect 149651 79867 149717 79868
rect 151123 79932 151189 79933
rect 151123 79868 151124 79932
rect 151188 79868 151189 79932
rect 151123 79867 151189 79868
rect 151307 79932 151373 79933
rect 151307 79868 151308 79932
rect 151372 79868 151373 79932
rect 151307 79867 151373 79868
rect 148915 79660 148981 79661
rect 148915 79596 148916 79660
rect 148980 79596 148981 79660
rect 148915 79595 148981 79596
rect 149470 78845 149530 79867
rect 149467 78844 149533 78845
rect 149467 78780 149468 78844
rect 149532 78780 149533 78844
rect 149467 78779 149533 78780
rect 149467 78708 149533 78709
rect 149467 78644 149468 78708
rect 149532 78644 149533 78708
rect 149467 78643 149533 78644
rect 149099 78572 149165 78573
rect 149099 78508 149100 78572
rect 149164 78508 149165 78572
rect 149099 78507 149165 78508
rect 148363 72724 148429 72725
rect 148363 72660 148364 72724
rect 148428 72660 148429 72724
rect 148363 72659 148429 72660
rect 148731 72724 148797 72725
rect 148731 72660 148732 72724
rect 148796 72660 148797 72724
rect 148731 72659 148797 72660
rect 148179 71228 148245 71229
rect 148179 71164 148180 71228
rect 148244 71164 148245 71228
rect 148179 71163 148245 71164
rect 148182 70410 148242 71163
rect 148182 70350 148426 70410
rect 147995 68916 148061 68917
rect 147995 68852 147996 68916
rect 148060 68852 148061 68916
rect 147995 68851 148061 68852
rect 147811 68508 147877 68509
rect 147811 68444 147812 68508
rect 147876 68444 147877 68508
rect 147811 68443 147877 68444
rect 148179 68508 148245 68509
rect 148179 68444 148180 68508
rect 148244 68444 148245 68508
rect 148179 68443 148245 68444
rect 147259 65516 147325 65517
rect 147259 65452 147260 65516
rect 147324 65452 147325 65516
rect 147259 65451 147325 65452
rect 147075 50284 147141 50285
rect 147075 50220 147076 50284
rect 147140 50220 147141 50284
rect 147075 50219 147141 50220
rect 146891 43484 146957 43485
rect 146891 43420 146892 43484
rect 146956 43420 146957 43484
rect 146891 43419 146957 43420
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145419 22676 145485 22677
rect 145419 22612 145420 22676
rect 145484 22612 145485 22676
rect 145419 22611 145485 22612
rect 144315 15876 144381 15877
rect 144315 15812 144316 15876
rect 144380 15812 144381 15876
rect 144315 15811 144381 15812
rect 144131 7580 144197 7581
rect 144131 7516 144132 7580
rect 144196 7516 144197 7580
rect 144131 7515 144197 7516
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 3454 146414 38898
rect 148182 28253 148242 68443
rect 148366 30973 148426 70350
rect 148547 68916 148613 68917
rect 148547 68852 148548 68916
rect 148612 68852 148613 68916
rect 148547 68851 148613 68852
rect 148550 54501 148610 68851
rect 148734 62797 148794 72659
rect 149102 68645 149162 78507
rect 149283 78436 149349 78437
rect 149283 78372 149284 78436
rect 149348 78372 149349 78436
rect 149283 78371 149349 78372
rect 149286 73949 149346 78371
rect 149470 74221 149530 78643
rect 149467 74220 149533 74221
rect 149467 74156 149468 74220
rect 149532 74156 149533 74220
rect 149467 74155 149533 74156
rect 149283 73948 149349 73949
rect 149283 73884 149284 73948
rect 149348 73884 149349 73948
rect 149283 73883 149349 73884
rect 149286 73810 149346 73883
rect 149286 73750 149530 73810
rect 149283 71500 149349 71501
rect 149283 71436 149284 71500
rect 149348 71436 149349 71500
rect 149283 71435 149349 71436
rect 149099 68644 149165 68645
rect 149099 68580 149100 68644
rect 149164 68580 149165 68644
rect 149099 68579 149165 68580
rect 148731 62796 148797 62797
rect 148731 62732 148732 62796
rect 148796 62732 148797 62796
rect 148731 62731 148797 62732
rect 149286 60750 149346 71435
rect 149470 66877 149530 73750
rect 149654 71501 149714 79867
rect 149835 74220 149901 74221
rect 149835 74156 149836 74220
rect 149900 74156 149901 74220
rect 149835 74155 149901 74156
rect 149651 71500 149717 71501
rect 149651 71436 149652 71500
rect 149716 71436 149717 71500
rect 149651 71435 149717 71436
rect 149467 66876 149533 66877
rect 149467 66812 149468 66876
rect 149532 66812 149533 66876
rect 149467 66811 149533 66812
rect 149286 60690 149714 60750
rect 148547 54500 148613 54501
rect 148547 54436 148548 54500
rect 148612 54436 148613 54500
rect 148547 54435 148613 54436
rect 149654 40765 149714 60690
rect 149838 45253 149898 74155
rect 150019 68644 150085 68645
rect 150019 68580 150020 68644
rect 150084 68580 150085 68644
rect 150019 68579 150085 68580
rect 150022 61709 150082 68579
rect 150019 61708 150085 61709
rect 150019 61644 150020 61708
rect 150084 61644 150085 61708
rect 150019 61643 150085 61644
rect 149835 45252 149901 45253
rect 149835 45188 149836 45252
rect 149900 45188 149901 45252
rect 149835 45187 149901 45188
rect 150294 43954 150914 78000
rect 151126 74221 151186 79867
rect 151310 79389 151370 79867
rect 151491 79796 151557 79797
rect 151491 79732 151492 79796
rect 151556 79732 151557 79796
rect 151491 79731 151557 79732
rect 151307 79388 151373 79389
rect 151307 79324 151308 79388
rect 151372 79324 151373 79388
rect 151307 79323 151373 79324
rect 151123 74220 151189 74221
rect 151123 74156 151124 74220
rect 151188 74156 151189 74220
rect 151123 74155 151189 74156
rect 151494 63477 151554 79731
rect 151491 63476 151557 63477
rect 151491 63412 151492 63476
rect 151556 63412 151557 63476
rect 151491 63411 151557 63412
rect 151678 59261 151738 80003
rect 153883 79932 153949 79933
rect 153883 79868 153884 79932
rect 153948 79868 153949 79932
rect 154251 79932 154317 79933
rect 154251 79930 154252 79932
rect 153883 79867 153949 79868
rect 154070 79870 154252 79930
rect 152411 79524 152477 79525
rect 152411 79460 152412 79524
rect 152476 79460 152477 79524
rect 152411 79459 152477 79460
rect 152414 71365 152474 79459
rect 152595 77756 152661 77757
rect 152595 77692 152596 77756
rect 152660 77692 152661 77756
rect 152595 77691 152661 77692
rect 152411 71364 152477 71365
rect 152411 71300 152412 71364
rect 152476 71300 152477 71364
rect 152411 71299 152477 71300
rect 151675 59260 151741 59261
rect 151675 59196 151676 59260
rect 151740 59196 151741 59260
rect 151675 59195 151741 59196
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 149651 40764 149717 40765
rect 149651 40700 149652 40764
rect 149716 40700 149717 40764
rect 149651 40699 149717 40700
rect 148363 30972 148429 30973
rect 148363 30908 148364 30972
rect 148428 30908 148429 30972
rect 148363 30907 148429 30908
rect 148179 28252 148245 28253
rect 148179 28188 148180 28252
rect 148244 28188 148245 28252
rect 148179 28187 148245 28188
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 7954 150914 43398
rect 152414 18597 152474 71299
rect 152598 46885 152658 77691
rect 152779 77212 152845 77213
rect 152779 77148 152780 77212
rect 152844 77148 152845 77212
rect 152779 77147 152845 77148
rect 152782 74357 152842 77147
rect 152779 74356 152845 74357
rect 152779 74292 152780 74356
rect 152844 74292 152845 74356
rect 152779 74291 152845 74292
rect 152595 46884 152661 46885
rect 152595 46820 152596 46884
rect 152660 46820 152661 46884
rect 152595 46819 152661 46820
rect 153886 39949 153946 79867
rect 154070 59125 154130 79870
rect 154251 79868 154252 79870
rect 154316 79868 154317 79932
rect 154251 79867 154317 79868
rect 155723 79932 155789 79933
rect 155723 79868 155724 79932
rect 155788 79868 155789 79932
rect 155723 79867 155789 79868
rect 156827 79932 156893 79933
rect 156827 79868 156828 79932
rect 156892 79868 156893 79932
rect 156827 79867 156893 79868
rect 157195 79932 157261 79933
rect 157195 79868 157196 79932
rect 157260 79868 157261 79932
rect 157195 79867 157261 79868
rect 154435 79796 154501 79797
rect 154435 79732 154436 79796
rect 154500 79732 154501 79796
rect 154435 79731 154501 79732
rect 155539 79796 155605 79797
rect 155539 79732 155540 79796
rect 155604 79732 155605 79796
rect 155539 79731 155605 79732
rect 154251 77212 154317 77213
rect 154251 77148 154252 77212
rect 154316 77148 154317 77212
rect 154251 77147 154317 77148
rect 154067 59124 154133 59125
rect 154067 59060 154068 59124
rect 154132 59060 154133 59124
rect 154067 59059 154133 59060
rect 154254 53821 154314 77147
rect 154438 73677 154498 79731
rect 154435 73676 154501 73677
rect 154435 73612 154436 73676
rect 154500 73612 154501 73676
rect 154435 73611 154501 73612
rect 154251 53820 154317 53821
rect 154251 53756 154252 53820
rect 154316 53756 154317 53820
rect 154251 53755 154317 53756
rect 154794 48454 155414 78000
rect 155542 66197 155602 79731
rect 155539 66196 155605 66197
rect 155539 66132 155540 66196
rect 155604 66132 155605 66196
rect 155539 66131 155605 66132
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 153883 39948 153949 39949
rect 153883 39884 153884 39948
rect 153948 39884 153949 39948
rect 153883 39883 153949 39884
rect 152411 18596 152477 18597
rect 152411 18532 152412 18596
rect 152476 18532 152477 18596
rect 152411 18531 152477 18532
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 12454 155414 47898
rect 155726 38589 155786 79867
rect 156643 78572 156709 78573
rect 156643 78508 156644 78572
rect 156708 78508 156709 78572
rect 156643 78507 156709 78508
rect 155723 38588 155789 38589
rect 155723 38524 155724 38588
rect 155788 38524 155789 38588
rect 155723 38523 155789 38524
rect 156646 17917 156706 78507
rect 156830 55181 156890 79867
rect 157011 78980 157077 78981
rect 157011 78916 157012 78980
rect 157076 78916 157077 78980
rect 157011 78915 157077 78916
rect 156827 55180 156893 55181
rect 156827 55116 156828 55180
rect 156892 55116 156893 55180
rect 156827 55115 156893 55116
rect 157014 35869 157074 78915
rect 157198 73133 157258 79867
rect 157931 78572 157997 78573
rect 157931 78508 157932 78572
rect 157996 78508 157997 78572
rect 157931 78507 157997 78508
rect 157195 73132 157261 73133
rect 157195 73068 157196 73132
rect 157260 73068 157261 73132
rect 157195 73067 157261 73068
rect 157011 35868 157077 35869
rect 157011 35804 157012 35868
rect 157076 35804 157077 35868
rect 157011 35803 157077 35804
rect 157934 21997 157994 78507
rect 158118 41309 158178 80139
rect 158851 80068 158917 80069
rect 158851 80004 158852 80068
rect 158916 80004 158917 80068
rect 158851 80003 158917 80004
rect 158299 79932 158365 79933
rect 158299 79868 158300 79932
rect 158364 79868 158365 79932
rect 158299 79867 158365 79868
rect 158115 41308 158181 41309
rect 158115 41244 158116 41308
rect 158180 41244 158181 41308
rect 158115 41243 158181 41244
rect 158302 30293 158362 79867
rect 158483 79796 158549 79797
rect 158483 79732 158484 79796
rect 158548 79732 158549 79796
rect 158483 79731 158549 79732
rect 158486 72997 158546 79731
rect 158483 72996 158549 72997
rect 158483 72932 158484 72996
rect 158548 72932 158549 72996
rect 158483 72931 158549 72932
rect 158854 49333 158914 80003
rect 164006 79933 164066 81227
rect 175411 81156 175477 81157
rect 175411 81092 175412 81156
rect 175476 81092 175477 81156
rect 175411 81091 175477 81092
rect 174307 81020 174373 81021
rect 174307 80956 174308 81020
rect 174372 80956 174373 81020
rect 174307 80955 174373 80956
rect 172283 80884 172349 80885
rect 172283 80820 172284 80884
rect 172348 80820 172349 80884
rect 172283 80819 172349 80820
rect 165107 80204 165173 80205
rect 165107 80140 165108 80204
rect 165172 80140 165173 80204
rect 165107 80139 165173 80140
rect 160875 79932 160941 79933
rect 160875 79868 160876 79932
rect 160940 79868 160941 79932
rect 160875 79867 160941 79868
rect 163267 79932 163333 79933
rect 163267 79868 163268 79932
rect 163332 79868 163333 79932
rect 163267 79867 163333 79868
rect 164003 79932 164069 79933
rect 164003 79868 164004 79932
rect 164068 79868 164069 79932
rect 164003 79867 164069 79868
rect 164187 79932 164253 79933
rect 164187 79868 164188 79932
rect 164252 79868 164253 79932
rect 164187 79867 164253 79868
rect 159035 78572 159101 78573
rect 159035 78508 159036 78572
rect 159100 78508 159101 78572
rect 159035 78507 159101 78508
rect 160691 78572 160757 78573
rect 160691 78508 160692 78572
rect 160756 78508 160757 78572
rect 160691 78507 160757 78508
rect 158851 49332 158917 49333
rect 158851 49268 158852 49332
rect 158916 49268 158917 49332
rect 158851 49267 158917 49268
rect 158299 30292 158365 30293
rect 158299 30228 158300 30292
rect 158364 30228 158365 30292
rect 158299 30227 158365 30228
rect 157931 21996 157997 21997
rect 157931 21932 157932 21996
rect 157996 21932 157997 21996
rect 157931 21931 157997 21932
rect 159038 21861 159098 78507
rect 159294 52954 159914 78000
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159035 21860 159101 21861
rect 159035 21796 159036 21860
rect 159100 21796 159101 21860
rect 159035 21795 159101 21796
rect 156643 17916 156709 17917
rect 156643 17852 156644 17916
rect 156708 17852 156709 17916
rect 156643 17851 156709 17852
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 16954 159914 52398
rect 160694 50965 160754 78507
rect 160878 54909 160938 79867
rect 162163 79660 162229 79661
rect 162163 79596 162164 79660
rect 162228 79596 162229 79660
rect 162163 79595 162229 79596
rect 162347 79660 162413 79661
rect 162347 79596 162348 79660
rect 162412 79596 162413 79660
rect 162347 79595 162413 79596
rect 161059 77484 161125 77485
rect 161059 77420 161060 77484
rect 161124 77420 161125 77484
rect 161059 77419 161125 77420
rect 160875 54908 160941 54909
rect 160875 54844 160876 54908
rect 160940 54844 160941 54908
rect 160875 54843 160941 54844
rect 161062 52189 161122 77419
rect 162166 53685 162226 79595
rect 162163 53684 162229 53685
rect 162163 53620 162164 53684
rect 162228 53620 162229 53684
rect 162163 53619 162229 53620
rect 161059 52188 161125 52189
rect 161059 52124 161060 52188
rect 161124 52124 161125 52188
rect 161059 52123 161125 52124
rect 160691 50964 160757 50965
rect 160691 50900 160692 50964
rect 160756 50900 160757 50964
rect 160691 50899 160757 50900
rect 162350 49469 162410 79595
rect 162531 77212 162597 77213
rect 162531 77148 162532 77212
rect 162596 77148 162597 77212
rect 162531 77147 162597 77148
rect 162347 49468 162413 49469
rect 162347 49404 162348 49468
rect 162412 49404 162413 49468
rect 162347 49403 162413 49404
rect 162534 45525 162594 77147
rect 162715 76532 162781 76533
rect 162715 76468 162716 76532
rect 162780 76468 162781 76532
rect 162715 76467 162781 76468
rect 162531 45524 162597 45525
rect 162531 45460 162532 45524
rect 162596 45460 162597 45524
rect 162531 45459 162597 45460
rect 162718 33013 162778 76467
rect 163270 52461 163330 79867
rect 163451 79388 163517 79389
rect 163451 79324 163452 79388
rect 163516 79324 163517 79388
rect 163451 79323 163517 79324
rect 163267 52460 163333 52461
rect 163267 52396 163268 52460
rect 163332 52396 163333 52460
rect 163267 52395 163333 52396
rect 162715 33012 162781 33013
rect 162715 32948 162716 33012
rect 162780 32948 162781 33012
rect 162715 32947 162781 32948
rect 163454 21725 163514 79323
rect 164006 79253 164066 79867
rect 164003 79252 164069 79253
rect 164003 79188 164004 79252
rect 164068 79188 164069 79252
rect 164003 79187 164069 79188
rect 164190 78165 164250 79867
rect 164923 78980 164989 78981
rect 164923 78916 164924 78980
rect 164988 78916 164989 78980
rect 164923 78915 164989 78916
rect 164187 78164 164253 78165
rect 164187 78100 164188 78164
rect 164252 78100 164253 78164
rect 164187 78099 164253 78100
rect 163635 75988 163701 75989
rect 163635 75924 163636 75988
rect 163700 75924 163701 75988
rect 163635 75923 163701 75924
rect 163638 48109 163698 75923
rect 163794 57454 164414 78000
rect 164926 62117 164986 78915
rect 164923 62116 164989 62117
rect 164923 62052 164924 62116
rect 164988 62052 164989 62116
rect 164923 62051 164989 62052
rect 165110 60349 165170 80139
rect 165291 79932 165357 79933
rect 165291 79868 165292 79932
rect 165356 79868 165357 79932
rect 165291 79867 165357 79868
rect 165659 79932 165725 79933
rect 165659 79868 165660 79932
rect 165724 79868 165725 79932
rect 165659 79867 165725 79868
rect 165843 79932 165909 79933
rect 165843 79868 165844 79932
rect 165908 79868 165909 79932
rect 165843 79867 165909 79868
rect 166395 79932 166461 79933
rect 166395 79868 166396 79932
rect 166460 79868 166461 79932
rect 166395 79867 166461 79868
rect 167867 79932 167933 79933
rect 167867 79868 167868 79932
rect 167932 79868 167933 79932
rect 167867 79867 167933 79868
rect 168971 79932 169037 79933
rect 168971 79868 168972 79932
rect 169036 79868 169037 79932
rect 168971 79867 169037 79868
rect 170259 79932 170325 79933
rect 170259 79868 170260 79932
rect 170324 79868 170325 79932
rect 170259 79867 170325 79868
rect 170627 79932 170693 79933
rect 170627 79868 170628 79932
rect 170692 79868 170693 79932
rect 170627 79867 170693 79868
rect 165294 76941 165354 79867
rect 165475 78300 165541 78301
rect 165475 78236 165476 78300
rect 165540 78236 165541 78300
rect 165475 78235 165541 78236
rect 165291 76940 165357 76941
rect 165291 76876 165292 76940
rect 165356 76876 165357 76940
rect 165291 76875 165357 76876
rect 165291 75988 165357 75989
rect 165291 75924 165292 75988
rect 165356 75924 165357 75988
rect 165291 75923 165357 75924
rect 165107 60348 165173 60349
rect 165107 60284 165108 60348
rect 165172 60284 165173 60348
rect 165107 60283 165173 60284
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163635 48108 163701 48109
rect 163635 48044 163636 48108
rect 163700 48044 163701 48108
rect 163635 48043 163701 48044
rect 163451 21724 163517 21725
rect 163451 21660 163452 21724
rect 163516 21660 163517 21724
rect 163451 21659 163517 21660
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 21454 164414 56898
rect 165294 50693 165354 75923
rect 165291 50692 165357 50693
rect 165291 50628 165292 50692
rect 165356 50628 165357 50692
rect 165291 50627 165357 50628
rect 165478 46749 165538 78235
rect 165662 75989 165722 79867
rect 165659 75988 165725 75989
rect 165659 75924 165660 75988
rect 165724 75924 165725 75988
rect 165659 75923 165725 75924
rect 165846 71790 165906 79867
rect 165846 71730 166274 71790
rect 166214 63205 166274 71730
rect 166211 63204 166277 63205
rect 166211 63140 166212 63204
rect 166276 63140 166277 63204
rect 166211 63139 166277 63140
rect 166398 57765 166458 79867
rect 166763 79796 166829 79797
rect 166763 79732 166764 79796
rect 166828 79732 166829 79796
rect 166763 79731 166829 79732
rect 166579 78572 166645 78573
rect 166579 78508 166580 78572
rect 166644 78508 166645 78572
rect 166579 78507 166645 78508
rect 166395 57764 166461 57765
rect 166395 57700 166396 57764
rect 166460 57700 166461 57764
rect 166395 57699 166461 57700
rect 166582 53549 166642 78507
rect 166579 53548 166645 53549
rect 166579 53484 166580 53548
rect 166644 53484 166645 53548
rect 166579 53483 166645 53484
rect 165475 46748 165541 46749
rect 165475 46684 165476 46748
rect 165540 46684 165541 46748
rect 165475 46683 165541 46684
rect 166766 45389 166826 79731
rect 167499 78572 167565 78573
rect 167499 78508 167500 78572
rect 167564 78508 167565 78572
rect 167499 78507 167565 78508
rect 167315 78436 167381 78437
rect 167315 78372 167316 78436
rect 167380 78372 167381 78436
rect 167315 78371 167381 78372
rect 167318 75989 167378 78371
rect 167315 75988 167381 75989
rect 167315 75924 167316 75988
rect 167380 75924 167381 75988
rect 167315 75923 167381 75924
rect 167502 52325 167562 78507
rect 167683 75988 167749 75989
rect 167683 75924 167684 75988
rect 167748 75924 167749 75988
rect 167683 75923 167749 75924
rect 167499 52324 167565 52325
rect 167499 52260 167500 52324
rect 167564 52260 167565 52324
rect 167499 52259 167565 52260
rect 167686 49605 167746 75923
rect 167683 49604 167749 49605
rect 167683 49540 167684 49604
rect 167748 49540 167749 49604
rect 167683 49539 167749 49540
rect 166763 45388 166829 45389
rect 166763 45324 166764 45388
rect 166828 45324 166829 45388
rect 166763 45323 166829 45324
rect 167870 35733 167930 79867
rect 168051 79796 168117 79797
rect 168051 79732 168052 79796
rect 168116 79732 168117 79796
rect 168051 79731 168117 79732
rect 167867 35732 167933 35733
rect 167867 35668 167868 35732
rect 167932 35668 167933 35732
rect 167867 35667 167933 35668
rect 168054 33149 168114 79731
rect 168974 78301 169034 79867
rect 170075 79796 170141 79797
rect 170075 79732 170076 79796
rect 170140 79732 170141 79796
rect 170075 79731 170141 79732
rect 169339 78980 169405 78981
rect 169339 78916 169340 78980
rect 169404 78916 169405 78980
rect 169339 78915 169405 78916
rect 168971 78300 169037 78301
rect 168971 78236 168972 78300
rect 169036 78236 169037 78300
rect 168971 78235 169037 78236
rect 168294 61954 168914 78000
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168051 33148 168117 33149
rect 168051 33084 168052 33148
rect 168116 33084 168117 33148
rect 168051 33083 168117 33084
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 25954 168914 61398
rect 169342 48245 169402 78915
rect 169523 78436 169589 78437
rect 169523 78372 169524 78436
rect 169588 78372 169589 78436
rect 169523 78371 169589 78372
rect 169339 48244 169405 48245
rect 169339 48180 169340 48244
rect 169404 48180 169405 48244
rect 169339 48179 169405 48180
rect 169526 47973 169586 78371
rect 170078 76941 170138 79731
rect 170075 76940 170141 76941
rect 170075 76876 170076 76940
rect 170140 76876 170141 76940
rect 170075 76875 170141 76876
rect 170262 76533 170322 79867
rect 170630 78573 170690 79867
rect 172286 79797 172346 80819
rect 173019 80476 173085 80477
rect 173019 80412 173020 80476
rect 173084 80412 173085 80476
rect 173019 80411 173085 80412
rect 171547 79796 171613 79797
rect 171547 79732 171548 79796
rect 171612 79732 171613 79796
rect 171547 79731 171613 79732
rect 172283 79796 172349 79797
rect 172283 79732 172284 79796
rect 172348 79732 172349 79796
rect 172283 79731 172349 79732
rect 172835 79796 172901 79797
rect 172835 79732 172836 79796
rect 172900 79732 172901 79796
rect 172835 79731 172901 79732
rect 170627 78572 170693 78573
rect 170627 78508 170628 78572
rect 170692 78508 170693 78572
rect 170627 78507 170693 78508
rect 170811 78436 170877 78437
rect 170811 78372 170812 78436
rect 170876 78372 170877 78436
rect 170811 78371 170877 78372
rect 170259 76532 170325 76533
rect 170259 76468 170260 76532
rect 170324 76468 170325 76532
rect 170259 76467 170325 76468
rect 170627 76532 170693 76533
rect 170627 76468 170628 76532
rect 170692 76468 170693 76532
rect 170627 76467 170693 76468
rect 170443 76124 170509 76125
rect 170443 76060 170444 76124
rect 170508 76060 170509 76124
rect 170443 76059 170509 76060
rect 170446 66061 170506 76059
rect 170443 66060 170509 66061
rect 170443 65996 170444 66060
rect 170508 65996 170509 66060
rect 170443 65995 170509 65996
rect 170630 58989 170690 76467
rect 170627 58988 170693 58989
rect 170627 58924 170628 58988
rect 170692 58924 170693 58988
rect 170627 58923 170693 58924
rect 170814 55045 170874 78371
rect 170995 76940 171061 76941
rect 170995 76876 170996 76940
rect 171060 76876 171061 76940
rect 170995 76875 171061 76876
rect 170811 55044 170877 55045
rect 170811 54980 170812 55044
rect 170876 54980 170877 55044
rect 170811 54979 170877 54980
rect 169523 47972 169589 47973
rect 169523 47908 169524 47972
rect 169588 47908 169589 47972
rect 169523 47907 169589 47908
rect 170998 46613 171058 76875
rect 171550 75853 171610 79731
rect 172838 78437 172898 79731
rect 173022 78981 173082 80411
rect 173387 79932 173453 79933
rect 173387 79868 173388 79932
rect 173452 79868 173453 79932
rect 173387 79867 173453 79868
rect 173019 78980 173085 78981
rect 173019 78916 173020 78980
rect 173084 78916 173085 78980
rect 173019 78915 173085 78916
rect 173390 78437 173450 79867
rect 173571 79796 173637 79797
rect 173571 79732 173572 79796
rect 173636 79732 173637 79796
rect 173571 79731 173637 79732
rect 172835 78436 172901 78437
rect 172835 78372 172836 78436
rect 172900 78372 172901 78436
rect 172835 78371 172901 78372
rect 173387 78436 173453 78437
rect 173387 78372 173388 78436
rect 173452 78372 173453 78436
rect 173387 78371 173453 78372
rect 171915 77756 171981 77757
rect 171915 77692 171916 77756
rect 171980 77692 171981 77756
rect 171915 77691 171981 77692
rect 171731 76532 171797 76533
rect 171731 76468 171732 76532
rect 171796 76468 171797 76532
rect 171731 76467 171797 76468
rect 171547 75852 171613 75853
rect 171547 75788 171548 75852
rect 171612 75788 171613 75852
rect 171547 75787 171613 75788
rect 171734 70277 171794 76467
rect 171731 70276 171797 70277
rect 171731 70212 171732 70276
rect 171796 70212 171797 70276
rect 171731 70211 171797 70212
rect 171918 65925 171978 77691
rect 172099 76532 172165 76533
rect 172099 76468 172100 76532
rect 172164 76468 172165 76532
rect 172099 76467 172165 76468
rect 172283 76532 172349 76533
rect 172283 76468 172284 76532
rect 172348 76468 172349 76532
rect 172283 76467 172349 76468
rect 171915 65924 171981 65925
rect 171915 65860 171916 65924
rect 171980 65860 171981 65924
rect 171915 65859 171981 65860
rect 172102 64837 172162 76467
rect 172099 64836 172165 64837
rect 172099 64772 172100 64836
rect 172164 64772 172165 64836
rect 172099 64771 172165 64772
rect 172286 62933 172346 76467
rect 172794 66454 173414 78000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172283 62932 172349 62933
rect 172283 62868 172284 62932
rect 172348 62868 172349 62932
rect 172283 62867 172349 62868
rect 170995 46612 171061 46613
rect 170995 46548 170996 46612
rect 171060 46548 171061 46612
rect 170995 46547 171061 46548
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 30454 173414 65898
rect 173574 60485 173634 79731
rect 174310 78981 174370 80955
rect 175227 80068 175293 80069
rect 175227 80004 175228 80068
rect 175292 80004 175293 80068
rect 175227 80003 175293 80004
rect 174675 79796 174741 79797
rect 174675 79732 174676 79796
rect 174740 79732 174741 79796
rect 174675 79731 174741 79732
rect 174307 78980 174373 78981
rect 174307 78916 174308 78980
rect 174372 78916 174373 78980
rect 174307 78915 174373 78916
rect 173755 77756 173821 77757
rect 173755 77692 173756 77756
rect 173820 77692 173821 77756
rect 173755 77691 173821 77692
rect 173571 60484 173637 60485
rect 173571 60420 173572 60484
rect 173636 60420 173637 60484
rect 173571 60419 173637 60420
rect 173758 44845 173818 77691
rect 174491 76940 174557 76941
rect 174491 76876 174492 76940
rect 174556 76876 174557 76940
rect 174491 76875 174557 76876
rect 174494 58853 174554 76875
rect 174491 58852 174557 58853
rect 174491 58788 174492 58852
rect 174556 58788 174557 58852
rect 174491 58787 174557 58788
rect 174678 57901 174738 79731
rect 174859 76532 174925 76533
rect 174859 76468 174860 76532
rect 174924 76468 174925 76532
rect 174859 76467 174925 76468
rect 175043 76532 175109 76533
rect 175043 76468 175044 76532
rect 175108 76468 175109 76532
rect 175043 76467 175109 76468
rect 174675 57900 174741 57901
rect 174675 57836 174676 57900
rect 174740 57836 174741 57900
rect 174675 57835 174741 57836
rect 174862 51781 174922 76467
rect 174859 51780 174925 51781
rect 174859 51716 174860 51780
rect 174924 51716 174925 51780
rect 174859 51715 174925 51716
rect 173755 44844 173821 44845
rect 173755 44780 173756 44844
rect 173820 44780 173821 44844
rect 173755 44779 173821 44780
rect 175046 44165 175106 76467
rect 175230 75581 175290 80003
rect 175414 79933 175474 81091
rect 181667 80748 181733 80749
rect 181667 80684 181668 80748
rect 181732 80684 181733 80748
rect 181667 80683 181733 80684
rect 181670 80205 181730 80683
rect 187739 80340 187805 80341
rect 187739 80276 187740 80340
rect 187804 80276 187805 80340
rect 187739 80275 187805 80276
rect 181667 80204 181733 80205
rect 181667 80140 181668 80204
rect 181732 80140 181733 80204
rect 181667 80139 181733 80140
rect 175411 79932 175477 79933
rect 175411 79868 175412 79932
rect 175476 79868 175477 79932
rect 176515 79932 176581 79933
rect 176515 79930 176516 79932
rect 175411 79867 175477 79868
rect 176334 79870 176516 79930
rect 175414 78437 175474 79867
rect 175963 79796 176029 79797
rect 175963 79732 175964 79796
rect 176028 79732 176029 79796
rect 175963 79731 176029 79732
rect 175411 78436 175477 78437
rect 175411 78372 175412 78436
rect 175476 78372 175477 78436
rect 175411 78371 175477 78372
rect 175227 75580 175293 75581
rect 175227 75516 175228 75580
rect 175292 75516 175293 75580
rect 175227 75515 175293 75516
rect 175966 63341 176026 79731
rect 176147 76940 176213 76941
rect 176147 76876 176148 76940
rect 176212 76876 176213 76940
rect 176147 76875 176213 76876
rect 175963 63340 176029 63341
rect 175963 63276 175964 63340
rect 176028 63276 176029 63340
rect 175963 63275 176029 63276
rect 176150 61981 176210 76875
rect 176147 61980 176213 61981
rect 176147 61916 176148 61980
rect 176212 61916 176213 61980
rect 176147 61915 176213 61916
rect 176334 50829 176394 79870
rect 176515 79868 176516 79870
rect 176580 79868 176581 79932
rect 176515 79867 176581 79868
rect 176515 76260 176581 76261
rect 176515 76196 176516 76260
rect 176580 76196 176581 76260
rect 176515 76195 176581 76196
rect 176331 50828 176397 50829
rect 176331 50764 176332 50828
rect 176396 50764 176397 50828
rect 176331 50763 176397 50764
rect 176518 48925 176578 76195
rect 177294 70954 177914 78000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 176515 48924 176581 48925
rect 176515 48860 176516 48924
rect 176580 48860 176581 48924
rect 176515 48859 176581 48860
rect 175043 44164 175109 44165
rect 175043 44100 175044 44164
rect 175108 44100 175109 44164
rect 175043 44099 175109 44100
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 75454 182414 78000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 78000
rect 187742 67421 187802 80275
rect 189214 67557 189274 107070
rect 189395 107068 189396 107070
rect 189460 107068 189461 107132
rect 189395 107067 189461 107068
rect 189582 103530 189642 113323
rect 189398 103470 189642 103530
rect 189398 79253 189458 103470
rect 189395 79252 189461 79253
rect 189395 79188 189396 79252
rect 189460 79188 189461 79252
rect 189395 79187 189461 79188
rect 189211 67556 189277 67557
rect 189211 67492 189212 67556
rect 189276 67492 189277 67556
rect 189211 67491 189277 67492
rect 187739 67420 187805 67421
rect 187739 67356 187740 67420
rect 187804 67356 187805 67420
rect 187739 67355 187805 67356
rect 189766 52053 189826 144739
rect 190794 142000 191414 155898
rect 191603 148476 191669 148477
rect 191603 148412 191604 148476
rect 191668 148412 191669 148476
rect 191603 148411 191669 148412
rect 190683 140316 190749 140317
rect 190683 140252 190684 140316
rect 190748 140252 190749 140316
rect 190683 140251 190749 140252
rect 190499 139908 190565 139909
rect 190499 139844 190500 139908
rect 190564 139844 190565 139908
rect 190499 139843 190565 139844
rect 190502 79525 190562 139843
rect 190499 79524 190565 79525
rect 190499 79460 190500 79524
rect 190564 79460 190565 79524
rect 190499 79459 190565 79460
rect 190686 79117 190746 140251
rect 191606 114477 191666 148411
rect 191787 146164 191853 146165
rect 191787 146100 191788 146164
rect 191852 146100 191853 146164
rect 191787 146099 191853 146100
rect 191603 114476 191669 114477
rect 191603 114412 191604 114476
rect 191668 114412 191669 114476
rect 191603 114411 191669 114412
rect 191603 81564 191669 81565
rect 191603 81500 191604 81564
rect 191668 81500 191669 81564
rect 191603 81499 191669 81500
rect 190683 79116 190749 79117
rect 190683 79052 190684 79116
rect 190748 79052 190749 79116
rect 190683 79051 190749 79052
rect 189763 52052 189829 52053
rect 189763 51988 189764 52052
rect 189828 51988 189829 52052
rect 189763 51987 189829 51988
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 48454 191414 78000
rect 191606 70005 191666 81499
rect 191603 70004 191669 70005
rect 191603 69940 191604 70004
rect 191668 69940 191669 70004
rect 191603 69939 191669 69940
rect 191790 49333 191850 146099
rect 191971 145892 192037 145893
rect 191971 145828 191972 145892
rect 192036 145828 192037 145892
rect 191971 145827 192037 145828
rect 191974 81293 192034 145827
rect 193262 144669 193322 262379
rect 193259 144668 193325 144669
rect 193259 144604 193260 144668
rect 193324 144604 193325 144668
rect 193259 144603 193325 144604
rect 193446 144533 193506 262515
rect 195294 232954 195914 268398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 198779 265028 198845 265029
rect 198779 264964 198780 265028
rect 198844 264964 198845 265028
rect 198779 264963 198845 264964
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 196019 196892 196085 196893
rect 196019 196828 196020 196892
rect 196084 196828 196085 196892
rect 196019 196827 196085 196828
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 193627 148612 193693 148613
rect 193627 148548 193628 148612
rect 193692 148548 193693 148612
rect 193627 148547 193693 148548
rect 193443 144532 193509 144533
rect 193443 144468 193444 144532
rect 193508 144468 193509 144532
rect 193443 144467 193509 144468
rect 193443 140724 193509 140725
rect 193443 140660 193444 140724
rect 193508 140660 193509 140724
rect 193443 140659 193509 140660
rect 192155 139772 192221 139773
rect 192155 139708 192156 139772
rect 192220 139708 192221 139772
rect 192155 139707 192221 139708
rect 191971 81292 192037 81293
rect 191971 81228 191972 81292
rect 192036 81228 192037 81292
rect 191971 81227 192037 81228
rect 192158 79389 192218 139707
rect 193446 80477 193506 140659
rect 193443 80476 193509 80477
rect 193443 80412 193444 80476
rect 193508 80412 193509 80476
rect 193443 80411 193509 80412
rect 192155 79388 192221 79389
rect 192155 79324 192156 79388
rect 192220 79324 192221 79388
rect 192155 79323 192221 79324
rect 193630 60621 193690 148547
rect 194547 140180 194613 140181
rect 194547 140116 194548 140180
rect 194612 140116 194613 140180
rect 194547 140115 194613 140116
rect 193627 60620 193693 60621
rect 193627 60556 193628 60620
rect 193692 60556 193693 60620
rect 193627 60555 193693 60556
rect 194550 53549 194610 140115
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 194547 53548 194613 53549
rect 194547 53484 194548 53548
rect 194612 53484 194613 53548
rect 194547 53483 194613 53484
rect 194550 53141 194610 53483
rect 194547 53140 194613 53141
rect 194547 53076 194548 53140
rect 194612 53076 194613 53140
rect 194547 53075 194613 53076
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 191787 49332 191853 49333
rect 191787 49268 191788 49332
rect 191852 49268 191853 49332
rect 191787 49267 191853 49268
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 16954 195914 52398
rect 196022 45525 196082 196827
rect 196203 193084 196269 193085
rect 196203 193020 196204 193084
rect 196268 193020 196269 193084
rect 196203 193019 196269 193020
rect 196206 75445 196266 193019
rect 196387 151332 196453 151333
rect 196387 151268 196388 151332
rect 196452 151268 196453 151332
rect 196387 151267 196453 151268
rect 196390 82245 196450 151267
rect 197307 151196 197373 151197
rect 197307 151132 197308 151196
rect 197372 151132 197373 151196
rect 197307 151131 197373 151132
rect 196387 82244 196453 82245
rect 196387 82180 196388 82244
rect 196452 82180 196453 82244
rect 196387 82179 196453 82180
rect 197310 78573 197370 151131
rect 197675 147524 197741 147525
rect 197675 147460 197676 147524
rect 197740 147460 197741 147524
rect 197675 147459 197741 147460
rect 197491 147388 197557 147389
rect 197491 147324 197492 147388
rect 197556 147324 197557 147388
rect 197491 147323 197557 147324
rect 197307 78572 197373 78573
rect 197307 78508 197308 78572
rect 197372 78508 197373 78572
rect 197307 78507 197373 78508
rect 197494 76669 197554 147323
rect 197678 80613 197738 147459
rect 198782 145757 198842 264963
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 203011 199340 203077 199341
rect 203011 199276 203012 199340
rect 203076 199276 203077 199340
rect 203011 199275 203077 199276
rect 200803 199204 200869 199205
rect 200803 199140 200804 199204
rect 200868 199140 200869 199204
rect 200803 199139 200869 199140
rect 200619 197436 200685 197437
rect 200619 197372 200620 197436
rect 200684 197372 200685 197436
rect 200619 197371 200685 197372
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199147 147252 199213 147253
rect 199147 147188 199148 147252
rect 199212 147188 199213 147252
rect 199147 147187 199213 147188
rect 198779 145756 198845 145757
rect 198779 145692 198780 145756
rect 198844 145692 198845 145756
rect 198779 145691 198845 145692
rect 198963 138140 199029 138141
rect 198963 138076 198964 138140
rect 199028 138076 199029 138140
rect 198963 138075 199029 138076
rect 197675 80612 197741 80613
rect 197675 80548 197676 80612
rect 197740 80548 197741 80612
rect 197675 80547 197741 80548
rect 198966 78573 199026 138075
rect 198963 78572 199029 78573
rect 198963 78508 198964 78572
rect 199028 78508 199029 78572
rect 198963 78507 199029 78508
rect 197491 76668 197557 76669
rect 197491 76604 197492 76668
rect 197556 76604 197557 76668
rect 197491 76603 197557 76604
rect 196203 75444 196269 75445
rect 196203 75380 196204 75444
rect 196268 75380 196269 75444
rect 196203 75379 196269 75380
rect 199150 75309 199210 147187
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199147 75308 199213 75309
rect 199147 75244 199148 75308
rect 199212 75244 199213 75308
rect 199147 75243 199213 75244
rect 199794 57454 200414 92898
rect 200622 64837 200682 197371
rect 200806 80069 200866 199139
rect 201539 198524 201605 198525
rect 201539 198460 201540 198524
rect 201604 198460 201605 198524
rect 201539 198459 201605 198460
rect 200987 150108 201053 150109
rect 200987 150044 200988 150108
rect 201052 150044 201053 150108
rect 200987 150043 201053 150044
rect 200803 80068 200869 80069
rect 200803 80004 200804 80068
rect 200868 80004 200869 80068
rect 200803 80003 200869 80004
rect 200990 76533 201050 150043
rect 200987 76532 201053 76533
rect 200987 76468 200988 76532
rect 201052 76468 201053 76532
rect 200987 76467 201053 76468
rect 200619 64836 200685 64837
rect 200619 64772 200620 64836
rect 200684 64772 200685 64836
rect 200619 64771 200685 64772
rect 201542 62933 201602 198459
rect 202827 197844 202893 197845
rect 202827 197780 202828 197844
rect 202892 197780 202893 197844
rect 202827 197779 202893 197780
rect 201723 195940 201789 195941
rect 201723 195876 201724 195940
rect 201788 195876 201789 195940
rect 201723 195875 201789 195876
rect 201726 71093 201786 195875
rect 202830 74550 202890 197779
rect 203014 79250 203074 199275
rect 204294 169954 204914 205398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 205035 199068 205101 199069
rect 205035 199004 205036 199068
rect 205100 199004 205101 199068
rect 205035 199003 205101 199004
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 203195 152828 203261 152829
rect 203195 152764 203196 152828
rect 203260 152764 203261 152828
rect 203195 152763 203261 152764
rect 203198 93870 203258 152763
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 203198 93810 203442 93870
rect 203014 79190 203258 79250
rect 202830 74490 203074 74550
rect 201723 71092 201789 71093
rect 201723 71028 201724 71092
rect 201788 71028 201789 71092
rect 201723 71027 201789 71028
rect 201539 62932 201605 62933
rect 201539 62868 201540 62932
rect 201604 62868 201605 62932
rect 201539 62867 201605 62868
rect 203014 61981 203074 74490
rect 203198 68237 203258 79190
rect 203382 75581 203442 93810
rect 203379 75580 203445 75581
rect 203379 75516 203380 75580
rect 203444 75516 203445 75580
rect 203379 75515 203445 75516
rect 203195 68236 203261 68237
rect 203195 68172 203196 68236
rect 203260 68172 203261 68236
rect 203195 68171 203261 68172
rect 203011 61980 203077 61981
rect 203011 61916 203012 61980
rect 203076 61916 203077 61980
rect 203011 61915 203077 61916
rect 204115 61980 204181 61981
rect 204115 61916 204116 61980
rect 204180 61916 204181 61980
rect 204115 61915 204181 61916
rect 204294 61954 204914 97398
rect 205038 67557 205098 199003
rect 205219 198932 205285 198933
rect 205219 198868 205220 198932
rect 205284 198868 205285 198932
rect 205219 198867 205285 198868
rect 205222 70141 205282 198867
rect 207059 194444 207125 194445
rect 207059 194380 207060 194444
rect 207124 194380 207125 194444
rect 207059 194379 207125 194380
rect 205587 194308 205653 194309
rect 205587 194244 205588 194308
rect 205652 194244 205653 194308
rect 205587 194243 205653 194244
rect 205590 75853 205650 194243
rect 205771 194172 205837 194173
rect 205771 194108 205772 194172
rect 205836 194108 205837 194172
rect 205771 194107 205837 194108
rect 205774 75853 205834 194107
rect 206139 149972 206205 149973
rect 206139 149908 206140 149972
rect 206204 149908 206205 149972
rect 206139 149907 206205 149908
rect 205955 149836 206021 149837
rect 205955 149772 205956 149836
rect 206020 149772 206021 149836
rect 205955 149771 206021 149772
rect 205587 75852 205653 75853
rect 205587 75788 205588 75852
rect 205652 75788 205653 75852
rect 205587 75787 205653 75788
rect 205771 75852 205837 75853
rect 205771 75788 205772 75852
rect 205836 75788 205837 75852
rect 205771 75787 205837 75788
rect 205219 70140 205285 70141
rect 205219 70076 205220 70140
rect 205284 70076 205285 70140
rect 205219 70075 205285 70076
rect 205222 69597 205282 70075
rect 205219 69596 205285 69597
rect 205219 69532 205220 69596
rect 205284 69532 205285 69596
rect 205219 69531 205285 69532
rect 205035 67556 205101 67557
rect 205035 67492 205036 67556
rect 205100 67492 205101 67556
rect 205035 67491 205101 67492
rect 204118 61437 204178 61915
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204115 61436 204181 61437
rect 204115 61372 204116 61436
rect 204180 61372 204181 61436
rect 204115 61371 204181 61372
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 196019 45524 196085 45525
rect 196019 45460 196020 45524
rect 196084 45460 196085 45524
rect 196019 45459 196085 45460
rect 196022 45117 196082 45459
rect 196019 45116 196085 45117
rect 196019 45052 196020 45116
rect 196084 45052 196085 45116
rect 196019 45051 196085 45052
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 25954 204914 61398
rect 205958 45525 206018 149771
rect 206142 78981 206202 149907
rect 206139 78980 206205 78981
rect 206139 78916 206140 78980
rect 206204 78916 206205 78980
rect 206139 78915 206205 78916
rect 205955 45524 206021 45525
rect 205955 45460 205956 45524
rect 206020 45460 206021 45524
rect 205955 45459 206021 45460
rect 207062 44845 207122 194379
rect 208794 174454 209414 209898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 209819 190228 209885 190229
rect 209819 190164 209820 190228
rect 209884 190164 209885 190228
rect 209819 190163 209885 190164
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 207243 149700 207309 149701
rect 207243 149636 207244 149700
rect 207308 149636 207309 149700
rect 207243 149635 207309 149636
rect 207246 71637 207306 149635
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 207243 71636 207309 71637
rect 207243 71572 207244 71636
rect 207308 71572 207309 71636
rect 207243 71571 207309 71572
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 207059 44844 207125 44845
rect 207059 44780 207060 44844
rect 207124 44780 207125 44844
rect 207059 44779 207125 44780
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 30454 209414 65898
rect 209822 50829 209882 190163
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 211107 157996 211173 157997
rect 211107 157932 211108 157996
rect 211172 157932 211173 157996
rect 211107 157931 211173 157932
rect 210003 152420 210069 152421
rect 210003 152356 210004 152420
rect 210068 152356 210069 152420
rect 210003 152355 210069 152356
rect 209819 50828 209885 50829
rect 209819 50764 209820 50828
rect 209884 50764 209885 50828
rect 209819 50763 209885 50764
rect 210006 44165 210066 152355
rect 211110 77893 211170 157931
rect 211291 155412 211357 155413
rect 211291 155348 211292 155412
rect 211356 155348 211357 155412
rect 211291 155347 211357 155348
rect 211294 78165 211354 155347
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 211291 78164 211357 78165
rect 211291 78100 211292 78164
rect 211356 78100 211357 78164
rect 211291 78099 211357 78100
rect 211107 77892 211173 77893
rect 211107 77828 211108 77892
rect 211172 77828 211173 77892
rect 211107 77827 211173 77828
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 211107 50828 211173 50829
rect 211107 50764 211108 50828
rect 211172 50764 211173 50828
rect 211107 50763 211173 50764
rect 211110 50285 211170 50763
rect 211107 50284 211173 50285
rect 211107 50220 211108 50284
rect 211172 50220 211173 50284
rect 211107 50219 211173 50220
rect 210003 44164 210069 44165
rect 210003 44100 210004 44164
rect 210068 44100 210069 44164
rect 210003 44099 210069 44100
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 124250 255218 124486 255454
rect 124250 254898 124486 255134
rect 154970 255218 155206 255454
rect 154970 254898 155206 255134
rect 185690 255218 185926 255454
rect 185690 254898 185926 255134
rect 139610 223718 139846 223954
rect 139610 223398 139846 223634
rect 170330 223718 170566 223954
rect 170330 223398 170566 223634
rect 124250 219218 124486 219454
rect 124250 218898 124486 219134
rect 154970 219218 155206 219454
rect 154970 218898 155206 219134
rect 185690 219218 185926 219454
rect 185690 218898 185926 219134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 139610 115718 139846 115954
rect 139610 115398 139846 115634
rect 170330 115718 170566 115954
rect 170330 115398 170566 115634
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 185690 111218 185926 111454
rect 185690 110898 185926 111134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 124250 255454
rect 124486 255218 154970 255454
rect 155206 255218 185690 255454
rect 185926 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 124250 255134
rect 124486 254898 154970 255134
rect 155206 254898 185690 255134
rect 185926 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 139610 223954
rect 139846 223718 170330 223954
rect 170566 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 139610 223634
rect 139846 223398 170330 223634
rect 170566 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 124250 219454
rect 124486 219218 154970 219454
rect 155206 219218 185690 219454
rect 185926 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 124250 219134
rect 124486 218898 154970 219134
rect 155206 218898 185690 219134
rect 185926 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 139610 115954
rect 139846 115718 170330 115954
rect 170566 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 139610 115634
rect 139846 115398 170330 115634
rect 170566 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 154970 111454
rect 155206 111218 185690 111454
rect 185926 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 154970 111134
rect 155206 110898 185690 111134
rect 185926 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use pixel_macro  pixel_macro0
timestamp 0
transform 1 0 120000 0 1 200000
box 1066 0 68854 60000
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 120000 0 1 80000
box 1066 0 70000 60000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 142000 146414 198000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 262000 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 142000 182414 198000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 262000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 142000 119414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 262000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 142000 155414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 262000 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 142000 191414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 262000 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 262000 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 262000 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 262000 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 262000 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 262000 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 262000 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 142000 141914 198000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 262000 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 142000 177914 198000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 262000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 142000 150914 198000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 262000 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 142000 186914 198000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 262000 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 142000 123914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 262000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 142000 159914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 262000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
