VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO SystemLevel
  CLASS BLOCK ;
  FOREIGN SystemLevel ;
  ORIGIN 65.000 72.400 ;
  SIZE 150.600 BY 162.400 ;
  PIN Aout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.350000 ;
    PORT
      LAYER li1 ;
        RECT 21.750 11.730 21.920 12.770 ;
        RECT 23.030 11.730 23.200 12.770 ;
        RECT 27.000 11.730 27.170 12.770 ;
        RECT 28.280 11.730 28.450 12.770 ;
        RECT 32.250 11.730 32.420 12.770 ;
        RECT 33.530 11.730 33.700 12.770 ;
        RECT 37.450 11.730 37.620 12.770 ;
        RECT 38.730 11.730 38.900 12.770 ;
        RECT 42.700 11.730 42.870 12.770 ;
        RECT 43.980 11.730 44.150 12.770 ;
        RECT 22.440 8.570 22.610 9.610 ;
        RECT 27.690 8.570 27.860 9.610 ;
        RECT 32.940 8.570 33.110 9.610 ;
        RECT 38.140 8.570 38.310 9.610 ;
        RECT 43.390 8.570 43.560 9.610 ;
      LAYER mcon ;
        RECT 21.750 11.810 21.920 12.690 ;
        RECT 23.030 11.810 23.200 12.690 ;
        RECT 27.000 11.810 27.170 12.690 ;
        RECT 28.280 11.810 28.450 12.690 ;
        RECT 32.250 11.810 32.420 12.690 ;
        RECT 33.530 11.810 33.700 12.690 ;
        RECT 37.450 11.810 37.620 12.690 ;
        RECT 38.730 11.810 38.900 12.690 ;
        RECT 42.700 11.810 42.870 12.690 ;
        RECT 43.980 11.810 44.150 12.690 ;
        RECT 22.440 8.650 22.610 9.530 ;
        RECT 27.690 8.650 27.860 9.530 ;
        RECT 32.940 8.650 33.110 9.530 ;
        RECT 38.140 8.650 38.310 9.530 ;
        RECT 43.390 8.650 43.560 9.530 ;
      LAYER met1 ;
        RECT 41.695 13.950 42.145 14.495 ;
        RECT 20.800 13.600 42.150 13.950 ;
        RECT 20.800 13.350 21.200 13.600 ;
        RECT 26.050 13.350 26.450 13.600 ;
        RECT 31.300 13.350 31.700 13.600 ;
        RECT 36.500 13.350 36.900 13.600 ;
        RECT 41.750 13.350 42.150 13.600 ;
        RECT 20.800 13.050 23.300 13.350 ;
        RECT 26.050 13.050 28.550 13.350 ;
        RECT 31.300 13.050 33.800 13.350 ;
        RECT 36.500 13.050 39.000 13.350 ;
        RECT 41.750 13.050 44.250 13.350 ;
        RECT 21.600 12.750 21.900 13.050 ;
        RECT 21.600 11.750 21.950 12.750 ;
        RECT 23.000 11.750 23.300 13.050 ;
        RECT 26.850 12.750 27.150 13.050 ;
        RECT 26.850 11.750 27.200 12.750 ;
        RECT 28.250 11.750 28.550 13.050 ;
        RECT 32.100 12.750 32.400 13.050 ;
        RECT 32.100 11.750 32.450 12.750 ;
        RECT 33.500 11.750 33.800 13.050 ;
        RECT 37.300 12.750 37.600 13.050 ;
        RECT 37.300 11.750 37.650 12.750 ;
        RECT 38.700 11.750 39.000 13.050 ;
        RECT 42.550 12.750 42.850 13.050 ;
        RECT 42.550 11.750 42.900 12.750 ;
        RECT 43.950 11.750 44.250 13.050 ;
        RECT 21.600 10.650 21.900 11.750 ;
        RECT 26.850 10.650 27.150 11.750 ;
        RECT 32.100 10.650 32.400 11.750 ;
        RECT 37.300 10.650 37.600 11.750 ;
        RECT 42.550 10.650 42.850 11.750 ;
        RECT 21.600 10.450 22.600 10.650 ;
        RECT 26.850 10.450 27.850 10.650 ;
        RECT 32.100 10.450 33.100 10.650 ;
        RECT 37.300 10.450 38.300 10.650 ;
        RECT 42.550 10.450 43.550 10.650 ;
        RECT 22.400 9.590 22.600 10.450 ;
        RECT 27.650 9.590 27.850 10.450 ;
        RECT 32.900 9.590 33.100 10.450 ;
        RECT 38.100 9.590 38.300 10.450 ;
        RECT 43.350 9.590 43.550 10.450 ;
        RECT 22.400 9.350 22.640 9.590 ;
        RECT 27.650 9.350 27.890 9.590 ;
        RECT 32.900 9.350 33.140 9.590 ;
        RECT 38.100 9.350 38.340 9.590 ;
        RECT 43.350 9.350 43.590 9.590 ;
        RECT 22.410 8.590 22.640 9.350 ;
        RECT 27.660 8.590 27.890 9.350 ;
        RECT 32.910 8.590 33.140 9.350 ;
        RECT 38.110 8.590 38.340 9.350 ;
        RECT 43.360 8.590 43.590 9.350 ;
      LAYER via ;
        RECT 41.695 14.015 42.145 14.465 ;
      LAYER met2 ;
        RECT 41.665 14.015 52.465 14.465 ;
        RECT 52.015 7.025 52.465 14.015 ;
        RECT 78.550 7.025 82.500 7.100 ;
        RECT 52.015 6.575 82.500 7.025 ;
        RECT 78.550 6.500 82.500 6.575 ;
    END
  END Aout
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 44.900 13.490 47.500 13.500 ;
        RECT 18.700 12.500 47.500 13.490 ;
        RECT 18.700 10.650 47.480 12.500 ;
        RECT -20.000 6.200 0.850 9.040 ;
        RECT -20.000 -3.150 -1.600 -0.200 ;
        RECT 3.500 -3.150 21.900 -0.200 ;
        RECT 23.750 -3.150 42.150 -0.200 ;
        RECT -20.000 -4.600 -1.680 -3.150 ;
        RECT 3.500 -4.600 21.820 -3.150 ;
        RECT 23.750 -4.600 42.070 -3.150 ;
        RECT -20.000 -5.400 -14.000 -4.600 ;
        RECT -20.000 -7.400 -14.040 -5.400 ;
        RECT -20.000 -8.400 -17.040 -7.400 ;
        RECT -7.300 -8.100 -1.760 -4.600 ;
        RECT 3.500 -5.400 9.500 -4.600 ;
        RECT 3.500 -7.400 9.460 -5.400 ;
        RECT 3.500 -8.400 6.460 -7.400 ;
        RECT 16.200 -8.100 21.740 -4.600 ;
        RECT 23.750 -5.400 29.750 -4.600 ;
        RECT 23.750 -7.400 29.710 -5.400 ;
        RECT 23.750 -8.400 26.710 -7.400 ;
        RECT 36.450 -8.100 41.990 -4.600 ;
        RECT 61.850 -16.510 62.900 -16.450 ;
        RECT 59.820 -19.350 72.850 -16.510 ;
        RECT 33.000 -22.450 35.960 -19.610 ;
        RECT 42.400 -26.650 60.800 -23.700 ;
        RECT 62.250 -26.650 80.650 -23.700 ;
        RECT 22.200 -29.160 38.060 -27.960 ;
        RECT 42.480 -28.100 60.800 -26.650 ;
        RECT 62.330 -28.100 80.650 -26.650 ;
        RECT 22.200 -32.000 40.960 -29.160 ;
        RECT 42.560 -31.600 48.100 -28.100 ;
        RECT 54.800 -28.900 60.800 -28.100 ;
        RECT 54.840 -30.900 60.800 -28.900 ;
        RECT 57.840 -31.900 60.800 -30.900 ;
        RECT 62.410 -31.600 67.950 -28.100 ;
        RECT 74.650 -28.900 80.650 -28.100 ;
        RECT 74.690 -30.900 80.650 -28.900 ;
        RECT 77.690 -31.900 80.650 -30.900 ;
      LAYER li1 ;
        RECT 17.150 13.530 45.450 13.550 ;
        RECT 17.150 13.130 47.530 13.530 ;
        RECT 17.150 13.100 45.530 13.130 ;
        RECT 17.150 13.050 44.850 13.100 ;
        RECT 17.150 13.000 19.100 13.050 ;
        RECT -21.925 9.000 0.800 9.100 ;
        RECT -22.000 8.600 0.800 9.000 ;
        RECT -22.000 8.550 -19.600 8.600 ;
        RECT -22.000 7.250 -20.750 8.550 ;
        RECT -19.900 8.200 -19.600 8.550 ;
        RECT -18.610 8.300 -18.440 8.320 ;
        RECT -18.100 8.300 -17.800 8.600 ;
        RECT -21.925 0.450 -20.875 7.250 ;
        RECT -19.820 6.785 -19.650 8.200 ;
        RECT -18.610 7.400 -17.800 8.300 ;
        RECT -17.600 8.200 -17.300 8.600 ;
        RECT -15.200 8.200 -14.900 8.600 ;
        RECT -14.700 8.200 -14.400 8.600 ;
        RECT -13.410 8.300 -13.240 8.320 ;
        RECT -12.900 8.300 -12.600 8.600 ;
        RECT -18.610 7.280 -18.440 7.400 ;
        RECT -18.040 6.785 -17.870 7.400 ;
        RECT -17.520 6.785 -17.350 8.200 ;
        RECT -15.100 6.785 -14.930 8.200 ;
        RECT -14.620 6.785 -14.450 8.200 ;
        RECT -13.410 7.400 -12.600 8.300 ;
        RECT -12.400 8.200 -12.100 8.600 ;
        RECT -10.000 8.200 -9.700 8.600 ;
        RECT -9.500 8.200 -9.200 8.600 ;
        RECT -8.210 8.300 -8.040 8.320 ;
        RECT -7.700 8.300 -7.400 8.600 ;
        RECT -13.410 7.280 -13.240 7.400 ;
        RECT -12.840 6.785 -12.670 7.400 ;
        RECT -12.320 6.785 -12.150 8.200 ;
        RECT -9.900 6.785 -9.730 8.200 ;
        RECT -9.420 6.785 -9.250 8.200 ;
        RECT -8.210 7.400 -7.400 8.300 ;
        RECT -7.200 8.200 -6.900 8.600 ;
        RECT -4.800 8.200 -4.500 8.600 ;
        RECT -4.300 8.200 -4.000 8.600 ;
        RECT -3.010 8.300 -2.840 8.320 ;
        RECT -2.500 8.300 -2.200 8.600 ;
        RECT -8.210 7.280 -8.040 7.400 ;
        RECT -7.640 6.785 -7.470 7.400 ;
        RECT -7.120 6.785 -6.950 8.200 ;
        RECT -4.700 6.785 -4.530 8.200 ;
        RECT -4.220 6.785 -4.050 8.200 ;
        RECT -3.010 7.400 -2.200 8.300 ;
        RECT -2.000 8.200 -1.700 8.600 ;
        RECT 0.400 8.200 0.700 8.600 ;
        RECT -3.010 7.280 -2.840 7.400 ;
        RECT -2.440 6.785 -2.270 7.400 ;
        RECT -1.920 6.785 -1.750 8.200 ;
        RECT 0.500 6.785 0.670 8.200 ;
        RECT 17.200 0.450 18.050 13.000 ;
        RECT 18.800 12.650 19.100 13.000 ;
        RECT 20.090 12.750 20.260 12.770 ;
        RECT 20.600 12.750 20.900 13.050 ;
        RECT 18.880 11.235 19.050 12.650 ;
        RECT 20.090 11.850 20.900 12.750 ;
        RECT 21.100 12.650 21.400 13.050 ;
        RECT 23.500 12.650 23.800 13.050 ;
        RECT 24.050 12.650 24.350 13.050 ;
        RECT 25.340 12.750 25.510 12.770 ;
        RECT 25.850 12.750 26.150 13.050 ;
        RECT 20.090 11.730 20.260 11.850 ;
        RECT 20.660 11.235 20.830 11.850 ;
        RECT 21.180 11.235 21.350 12.650 ;
        RECT 23.600 11.235 23.770 12.650 ;
        RECT 24.130 11.235 24.300 12.650 ;
        RECT 25.340 11.850 26.150 12.750 ;
        RECT 26.350 12.650 26.650 13.050 ;
        RECT 28.750 12.650 29.050 13.050 ;
        RECT 29.300 12.650 29.600 13.050 ;
        RECT 30.590 12.750 30.760 12.770 ;
        RECT 31.100 12.750 31.400 13.050 ;
        RECT 25.340 11.730 25.510 11.850 ;
        RECT 25.910 11.235 26.080 11.850 ;
        RECT 26.430 11.235 26.600 12.650 ;
        RECT 28.850 11.235 29.020 12.650 ;
        RECT 29.380 11.235 29.550 12.650 ;
        RECT 30.590 11.850 31.400 12.750 ;
        RECT 31.600 12.650 31.900 13.050 ;
        RECT 34.000 12.650 34.300 13.050 ;
        RECT 34.500 12.650 34.800 13.050 ;
        RECT 35.790 12.750 35.960 12.770 ;
        RECT 36.300 12.750 36.600 13.050 ;
        RECT 30.590 11.730 30.760 11.850 ;
        RECT 31.160 11.235 31.330 11.850 ;
        RECT 31.680 11.235 31.850 12.650 ;
        RECT 34.100 11.235 34.270 12.650 ;
        RECT 34.580 11.235 34.750 12.650 ;
        RECT 35.790 11.850 36.600 12.750 ;
        RECT 36.800 12.650 37.100 13.050 ;
        RECT 39.200 12.650 39.500 13.050 ;
        RECT 39.750 12.650 40.050 13.050 ;
        RECT 41.040 12.750 41.210 12.770 ;
        RECT 41.550 12.750 41.850 13.050 ;
        RECT 35.790 11.730 35.960 11.850 ;
        RECT 36.360 11.235 36.530 11.850 ;
        RECT 36.880 11.235 37.050 12.650 ;
        RECT 39.300 11.235 39.470 12.650 ;
        RECT 39.830 11.235 40.000 12.650 ;
        RECT 41.040 11.850 41.850 12.750 ;
        RECT 42.050 12.650 42.350 13.050 ;
        RECT 44.450 12.650 44.750 13.050 ;
        RECT 45.130 12.650 45.530 13.100 ;
        RECT 45.920 12.650 46.090 12.770 ;
        RECT 41.040 11.730 41.210 11.850 ;
        RECT 41.610 11.235 41.780 11.850 ;
        RECT 42.130 11.235 42.300 12.650 ;
        RECT 44.550 11.235 44.720 12.650 ;
        RECT 45.130 11.770 46.090 12.650 ;
        RECT 45.130 11.530 45.530 11.770 ;
        RECT 45.920 11.730 46.090 11.770 ;
        RECT 45.350 11.235 45.520 11.530 ;
        RECT 47.130 11.235 47.300 12.905 ;
        RECT 41.050 0.450 41.950 3.800 ;
        RECT -21.925 -0.450 42.000 0.450 ;
        RECT -21.925 -0.600 41.910 -0.450 ;
        RECT -20.000 -0.710 41.910 -0.600 ;
        RECT -20.000 -0.800 -19.300 -0.710 ;
        RECT -20.000 -4.250 -19.440 -0.800 ;
        RECT -11.230 -4.250 -10.450 -0.710 ;
        RECT -2.250 -0.750 4.250 -0.710 ;
        RECT -2.200 -3.150 -1.840 -0.750 ;
        RECT 3.500 -0.800 4.200 -0.750 ;
        RECT -2.200 -4.200 -1.850 -3.150 ;
        RECT -6.700 -4.250 -1.850 -4.200 ;
        RECT -20.000 -4.350 -1.850 -4.250 ;
        RECT -20.000 -4.420 -11.060 -4.350 ;
        RECT -10.620 -4.420 -1.850 -4.350 ;
        RECT -20.000 -4.600 -14.250 -4.420 ;
        RECT -20.000 -4.740 -14.240 -4.600 ;
        RECT -6.700 -4.730 -1.850 -4.420 ;
        RECT -20.000 -5.000 -14.220 -4.740 ;
        RECT -19.820 -5.040 -14.220 -5.000 ;
        RECT -19.820 -8.050 -19.650 -5.040 ;
        RECT -17.880 -5.280 -17.200 -5.040 ;
        RECT -17.960 -7.280 -17.200 -5.280 ;
        RECT -16.820 -7.050 -16.650 -5.040 ;
        RECT -14.880 -5.280 -14.220 -5.040 ;
        RECT -14.960 -6.280 -14.220 -5.280 ;
        RECT -14.960 -6.320 -14.790 -6.280 ;
        RECT -14.390 -7.050 -14.220 -6.280 ;
        RECT -16.820 -7.220 -14.220 -7.050 ;
        RECT -7.120 -4.900 -1.850 -4.730 ;
        RECT 3.500 -4.250 4.060 -0.800 ;
        RECT 12.270 -4.250 13.050 -0.710 ;
        RECT 21.250 -0.800 24.450 -0.710 ;
        RECT 21.300 -3.150 21.660 -0.800 ;
        RECT 21.300 -4.200 21.650 -3.150 ;
        RECT 16.800 -4.250 21.650 -4.200 ;
        RECT 3.500 -4.350 21.650 -4.250 ;
        RECT 3.500 -4.420 12.440 -4.350 ;
        RECT 12.880 -4.420 21.650 -4.350 ;
        RECT 3.500 -4.600 9.250 -4.420 ;
        RECT 3.500 -4.740 9.260 -4.600 ;
        RECT 16.800 -4.730 21.650 -4.420 ;
        RECT -17.960 -7.320 -17.790 -7.280 ;
        RECT -17.390 -8.050 -17.220 -7.280 ;
        RECT -7.120 -7.750 -6.950 -4.900 ;
        RECT -6.700 -5.600 -6.300 -4.900 ;
        RECT -4.100 -5.600 -3.700 -4.900 ;
        RECT -6.550 -7.020 -6.380 -5.600 ;
        RECT -3.970 -7.020 -3.800 -5.600 ;
        RECT -2.110 -7.750 -1.940 -4.900 ;
        RECT 3.500 -5.000 9.280 -4.740 ;
        RECT -7.120 -7.920 -1.940 -7.750 ;
        RECT 3.680 -5.040 9.280 -5.000 ;
        RECT -19.820 -8.220 -17.220 -8.050 ;
        RECT 3.680 -8.050 3.850 -5.040 ;
        RECT 5.620 -5.280 6.300 -5.040 ;
        RECT 5.540 -7.280 6.300 -5.280 ;
        RECT 6.680 -7.050 6.850 -5.040 ;
        RECT 8.620 -5.280 9.280 -5.040 ;
        RECT 8.540 -6.280 9.280 -5.280 ;
        RECT 8.540 -6.320 8.710 -6.280 ;
        RECT 9.110 -7.050 9.280 -6.280 ;
        RECT 6.680 -7.220 9.280 -7.050 ;
        RECT 16.380 -4.900 21.650 -4.730 ;
        RECT 23.750 -4.250 24.310 -0.800 ;
        RECT 32.520 -4.250 33.300 -0.710 ;
        RECT 41.550 -3.150 41.910 -0.710 ;
        RECT 41.550 -4.200 41.900 -3.150 ;
        RECT 37.050 -4.250 41.900 -4.200 ;
        RECT 23.750 -4.350 41.900 -4.250 ;
        RECT 23.750 -4.420 32.690 -4.350 ;
        RECT 33.130 -4.420 41.900 -4.350 ;
        RECT 23.750 -4.600 29.500 -4.420 ;
        RECT 23.750 -4.740 29.510 -4.600 ;
        RECT 37.050 -4.730 41.900 -4.420 ;
        RECT 5.540 -7.320 5.710 -7.280 ;
        RECT 6.110 -8.050 6.280 -7.280 ;
        RECT 16.380 -7.750 16.550 -4.900 ;
        RECT 16.800 -5.600 17.200 -4.900 ;
        RECT 19.400 -5.600 19.800 -4.900 ;
        RECT 16.950 -7.020 17.120 -5.600 ;
        RECT 19.530 -7.020 19.700 -5.600 ;
        RECT 21.390 -7.750 21.560 -4.900 ;
        RECT 23.750 -5.000 29.530 -4.740 ;
        RECT 16.380 -7.920 21.560 -7.750 ;
        RECT 23.930 -5.040 29.530 -5.000 ;
        RECT 3.680 -8.220 6.280 -8.050 ;
        RECT 23.930 -8.050 24.100 -5.040 ;
        RECT 25.870 -5.280 26.550 -5.040 ;
        RECT 25.790 -7.280 26.550 -5.280 ;
        RECT 26.930 -7.050 27.100 -5.040 ;
        RECT 28.870 -5.280 29.530 -5.040 ;
        RECT 28.790 -6.280 29.530 -5.280 ;
        RECT 28.790 -6.320 28.960 -6.280 ;
        RECT 29.360 -7.050 29.530 -6.280 ;
        RECT 26.930 -7.220 29.530 -7.050 ;
        RECT 36.630 -4.900 41.900 -4.730 ;
        RECT 25.790 -7.320 25.960 -7.280 ;
        RECT 26.360 -8.050 26.530 -7.280 ;
        RECT 36.630 -7.750 36.800 -4.900 ;
        RECT 37.050 -5.600 37.450 -4.900 ;
        RECT 39.650 -5.600 40.050 -4.900 ;
        RECT 37.200 -7.020 37.370 -5.600 ;
        RECT 39.780 -7.020 39.950 -5.600 ;
        RECT 41.640 -7.750 41.810 -4.900 ;
        RECT 36.630 -7.920 41.810 -7.750 ;
        RECT 23.930 -8.220 26.530 -8.050 ;
        RECT 33.100 -20.050 35.900 -19.750 ;
        RECT 33.100 -21.850 33.400 -20.050 ;
        RECT 35.040 -20.850 35.210 -20.690 ;
        RECT 35.600 -20.850 35.900 -20.050 ;
        RECT 36.100 -20.850 36.600 -15.600 ;
        RECT 62.050 -16.470 72.800 -16.450 ;
        RECT 59.700 -16.500 72.800 -16.470 ;
        RECT 55.800 -16.800 72.800 -16.500 ;
        RECT 55.800 -20.450 56.100 -16.800 ;
        RECT 59.700 -16.870 72.800 -16.800 ;
        RECT 59.780 -17.350 60.180 -16.870 ;
        RECT 62.050 -16.950 72.800 -16.870 ;
        RECT 60.570 -17.350 60.740 -17.230 ;
        RECT 59.780 -18.230 60.740 -17.350 ;
        RECT 59.780 -18.470 60.180 -18.230 ;
        RECT 60.570 -18.270 60.740 -18.230 ;
        RECT 60.000 -18.765 60.170 -18.470 ;
        RECT 61.780 -18.765 61.950 -17.095 ;
        RECT 62.450 -17.350 62.750 -16.950 ;
        RECT 63.740 -17.250 63.910 -17.230 ;
        RECT 64.250 -17.250 64.550 -16.950 ;
        RECT 62.530 -18.765 62.700 -17.350 ;
        RECT 63.740 -18.150 64.550 -17.250 ;
        RECT 64.750 -17.350 65.050 -16.950 ;
        RECT 67.150 -17.350 67.450 -16.950 ;
        RECT 67.700 -17.350 68.000 -16.950 ;
        RECT 68.990 -17.250 69.160 -17.230 ;
        RECT 69.500 -17.250 69.800 -16.950 ;
        RECT 63.740 -18.270 63.910 -18.150 ;
        RECT 64.310 -18.765 64.480 -18.150 ;
        RECT 64.830 -18.765 65.000 -17.350 ;
        RECT 67.250 -18.765 67.420 -17.350 ;
        RECT 67.780 -18.765 67.950 -17.350 ;
        RECT 68.990 -18.150 69.800 -17.250 ;
        RECT 70.000 -17.350 70.300 -16.950 ;
        RECT 72.400 -17.350 72.700 -16.950 ;
        RECT 68.990 -18.270 69.160 -18.150 ;
        RECT 69.560 -18.765 69.730 -18.150 ;
        RECT 70.080 -18.765 70.250 -17.350 ;
        RECT 72.500 -18.765 72.670 -17.350 ;
        RECT 35.040 -21.450 36.600 -20.850 ;
        RECT 35.040 -21.550 36.300 -21.450 ;
        RECT 35.040 -21.730 35.210 -21.550 ;
        RECT 33.180 -21.865 33.350 -21.850 ;
        RECT 35.610 -21.865 35.780 -21.550 ;
        RECT 55.500 -22.950 56.400 -20.450 ;
        RECT 51.150 -23.780 80.650 -22.950 ;
        RECT 42.640 -24.210 80.650 -23.780 ;
        RECT 42.640 -26.650 43.000 -24.210 ;
        RECT 29.900 -28.000 30.600 -27.050 ;
        RECT 42.650 -27.700 43.000 -26.650 ;
        RECT 42.650 -27.750 47.500 -27.700 ;
        RECT 51.250 -27.750 52.030 -24.210 ;
        RECT 60.100 -24.300 62.850 -24.210 ;
        RECT 60.240 -24.400 62.850 -24.300 ;
        RECT 60.240 -27.750 60.800 -24.400 ;
        RECT 62.490 -26.650 62.850 -24.400 ;
        RECT 42.650 -27.850 60.800 -27.750 ;
        RECT 42.650 -27.920 51.420 -27.850 ;
        RECT 51.860 -27.920 60.800 -27.850 ;
        RECT 22.300 -28.500 38.400 -28.000 ;
        RECT 42.650 -28.230 47.500 -27.920 ;
        RECT 55.050 -28.100 60.800 -27.920 ;
        RECT 42.650 -28.400 47.920 -28.230 ;
        RECT 55.040 -28.240 60.800 -28.100 ;
        RECT 22.380 -31.650 22.550 -28.500 ;
        RECT 24.200 -28.900 24.500 -28.500 ;
        RECT 26.700 -28.900 27.000 -28.500 ;
        RECT 29.300 -28.900 29.600 -28.500 ;
        RECT 31.900 -28.900 32.200 -28.500 ;
        RECT 34.500 -28.900 34.800 -28.500 ;
        RECT 37.100 -28.900 37.400 -28.500 ;
        RECT 24.240 -30.920 24.410 -28.900 ;
        RECT 26.820 -30.920 26.990 -28.900 ;
        RECT 29.400 -30.920 29.570 -28.900 ;
        RECT 31.980 -30.920 32.150 -28.900 ;
        RECT 34.560 -30.920 34.730 -28.900 ;
        RECT 37.140 -30.920 37.310 -28.900 ;
        RECT 37.710 -29.200 38.400 -28.500 ;
        RECT 37.710 -29.600 41.000 -29.200 ;
        RECT 37.710 -30.500 39.000 -29.600 ;
        RECT 37.710 -30.900 38.920 -30.500 ;
        RECT 37.710 -31.650 37.880 -30.900 ;
        RECT 22.380 -31.820 37.880 -31.650 ;
        RECT 38.180 -31.650 38.350 -30.900 ;
        RECT 38.750 -30.920 38.920 -30.900 ;
        RECT 40.610 -31.650 40.780 -29.600 ;
        RECT 42.740 -31.250 42.910 -28.400 ;
        RECT 44.500 -29.100 44.900 -28.400 ;
        RECT 47.100 -29.100 47.500 -28.400 ;
        RECT 44.600 -30.520 44.770 -29.100 ;
        RECT 47.180 -30.520 47.350 -29.100 ;
        RECT 47.750 -31.250 47.920 -28.400 ;
        RECT 55.020 -28.500 60.800 -28.240 ;
        RECT 62.500 -27.700 62.850 -26.650 ;
        RECT 62.500 -27.750 67.350 -27.700 ;
        RECT 71.100 -27.750 71.880 -24.210 ;
        RECT 79.950 -24.300 80.650 -24.210 ;
        RECT 80.090 -27.750 80.650 -24.300 ;
        RECT 62.500 -27.850 80.650 -27.750 ;
        RECT 62.500 -27.920 71.270 -27.850 ;
        RECT 71.710 -27.920 80.650 -27.850 ;
        RECT 62.500 -28.230 67.350 -27.920 ;
        RECT 74.900 -28.100 80.650 -27.920 ;
        RECT 62.500 -28.400 67.770 -28.230 ;
        RECT 74.890 -28.240 80.650 -28.100 ;
        RECT 55.020 -28.540 60.620 -28.500 ;
        RECT 55.020 -28.780 55.680 -28.540 ;
        RECT 55.020 -29.780 55.760 -28.780 ;
        RECT 55.020 -30.550 55.190 -29.780 ;
        RECT 55.590 -29.820 55.760 -29.780 ;
        RECT 57.450 -30.550 57.620 -28.540 ;
        RECT 55.020 -30.720 57.620 -30.550 ;
        RECT 58.000 -28.780 58.680 -28.540 ;
        RECT 58.000 -30.780 58.760 -28.780 ;
        RECT 42.740 -31.420 47.920 -31.250 ;
        RECT 38.180 -31.820 40.780 -31.650 ;
        RECT 58.020 -31.550 58.190 -30.780 ;
        RECT 58.590 -30.820 58.760 -30.780 ;
        RECT 60.450 -31.550 60.620 -28.540 ;
        RECT 62.590 -31.250 62.760 -28.400 ;
        RECT 64.350 -29.100 64.750 -28.400 ;
        RECT 66.950 -29.100 67.350 -28.400 ;
        RECT 64.450 -30.520 64.620 -29.100 ;
        RECT 67.030 -30.520 67.200 -29.100 ;
        RECT 67.600 -31.250 67.770 -28.400 ;
        RECT 74.870 -28.500 80.650 -28.240 ;
        RECT 74.870 -28.540 80.470 -28.500 ;
        RECT 74.870 -28.780 75.530 -28.540 ;
        RECT 74.870 -29.780 75.610 -28.780 ;
        RECT 74.870 -30.550 75.040 -29.780 ;
        RECT 75.440 -29.820 75.610 -29.780 ;
        RECT 77.300 -30.550 77.470 -28.540 ;
        RECT 74.870 -30.720 77.470 -30.550 ;
        RECT 77.850 -28.780 78.530 -28.540 ;
        RECT 77.850 -30.780 78.610 -28.780 ;
        RECT 62.590 -31.420 67.770 -31.250 ;
        RECT 58.020 -31.720 60.620 -31.550 ;
        RECT 77.870 -31.550 78.040 -30.780 ;
        RECT 78.440 -30.820 78.610 -30.780 ;
        RECT 80.300 -31.550 80.470 -28.540 ;
        RECT 77.870 -31.720 80.470 -31.550 ;
      LAYER mcon ;
        RECT -21.750 7.500 -21.000 8.750 ;
        RECT -18.610 7.360 -18.440 8.240 ;
        RECT -13.410 7.360 -13.240 8.240 ;
        RECT -8.210 7.360 -8.040 8.240 ;
        RECT -3.010 7.360 -2.840 8.240 ;
        RECT 20.090 11.810 20.260 12.690 ;
        RECT 25.340 11.810 25.510 12.690 ;
        RECT 30.590 11.810 30.760 12.690 ;
        RECT 35.790 11.810 35.960 12.690 ;
        RECT 41.040 11.810 41.210 12.690 ;
        RECT 45.920 11.810 46.090 12.690 ;
        RECT 41.050 2.900 41.950 3.800 ;
        RECT -17.960 -7.240 -17.790 -5.360 ;
        RECT -14.960 -6.240 -14.790 -5.360 ;
        RECT -6.550 -6.940 -6.380 -5.350 ;
        RECT -3.970 -6.940 -3.800 -5.350 ;
        RECT 5.540 -7.240 5.710 -5.360 ;
        RECT 8.540 -6.240 8.710 -5.360 ;
        RECT 16.950 -6.940 17.120 -5.350 ;
        RECT 19.530 -6.940 19.700 -5.350 ;
        RECT 25.790 -7.240 25.960 -5.360 ;
        RECT 28.790 -6.240 28.960 -5.360 ;
        RECT 37.200 -6.940 37.370 -5.350 ;
        RECT 39.780 -6.940 39.950 -5.350 ;
        RECT 36.100 -16.100 36.600 -15.600 ;
        RECT 35.040 -21.650 35.210 -20.770 ;
        RECT 60.570 -18.190 60.740 -17.310 ;
        RECT 63.740 -18.190 63.910 -17.310 ;
        RECT 68.990 -18.190 69.160 -17.310 ;
        RECT 55.530 -21.320 56.370 -20.480 ;
        RECT 29.900 -27.750 30.600 -27.050 ;
        RECT 24.240 -30.840 24.410 -28.760 ;
        RECT 26.820 -30.840 26.990 -28.760 ;
        RECT 29.400 -30.840 29.570 -28.760 ;
        RECT 31.980 -30.840 32.150 -28.760 ;
        RECT 34.560 -30.840 34.730 -28.760 ;
        RECT 37.140 -30.840 37.310 -28.760 ;
        RECT 38.750 -30.840 38.920 -29.960 ;
        RECT 44.600 -30.440 44.770 -28.850 ;
        RECT 47.180 -30.440 47.350 -28.850 ;
        RECT 55.590 -29.740 55.760 -28.860 ;
        RECT 58.590 -30.740 58.760 -28.860 ;
        RECT 64.450 -30.440 64.620 -28.850 ;
        RECT 67.030 -30.440 67.200 -28.850 ;
        RECT 75.440 -29.740 75.610 -28.860 ;
        RECT 78.440 -30.740 78.610 -28.860 ;
      LAYER met1 ;
        RECT 20.060 11.750 20.290 12.750 ;
        RECT 25.310 11.750 25.540 12.750 ;
        RECT 30.560 11.750 30.790 12.750 ;
        RECT 35.760 11.750 35.990 12.750 ;
        RECT 41.010 11.750 41.240 12.750 ;
        RECT 45.890 11.750 46.120 12.750 ;
        RECT -51.000 9.000 -48.000 9.030 ;
        RECT -51.000 6.000 -20.500 9.000 ;
        RECT -18.640 7.300 -18.410 8.300 ;
        RECT -13.440 7.300 -13.210 8.300 ;
        RECT -8.240 7.300 -8.010 8.300 ;
        RECT -3.040 7.300 -2.810 8.300 ;
        RECT -51.000 5.970 -48.000 6.000 ;
        RECT 40.990 3.800 42.010 3.830 ;
        RECT 44.250 3.800 45.350 3.900 ;
        RECT 40.990 2.900 45.350 3.800 ;
        RECT 40.990 2.870 42.010 2.900 ;
        RECT 44.250 2.800 45.350 2.900 ;
        RECT -17.990 -7.300 -17.760 -5.300 ;
        RECT -14.990 -6.300 -14.760 -5.300 ;
        RECT -6.580 -7.000 -6.350 -5.290 ;
        RECT -4.000 -7.000 -3.770 -5.290 ;
        RECT 5.510 -7.300 5.740 -5.300 ;
        RECT 8.510 -6.300 8.740 -5.300 ;
        RECT 16.920 -7.000 17.150 -5.290 ;
        RECT 19.500 -7.000 19.730 -5.290 ;
        RECT 25.760 -7.300 25.990 -5.300 ;
        RECT 28.760 -6.300 28.990 -5.300 ;
        RECT 37.170 -7.000 37.400 -5.290 ;
        RECT 39.750 -7.000 39.980 -5.290 ;
        RECT 35.150 -15.550 35.850 -15.520 ;
        RECT 35.150 -15.570 36.650 -15.550 ;
        RECT 35.150 -15.600 36.660 -15.570 ;
        RECT 44.450 -15.600 45.050 -15.550 ;
        RECT 35.150 -16.100 45.050 -15.600 ;
        RECT 35.150 -16.130 36.660 -16.100 ;
        RECT 35.150 -16.250 36.650 -16.130 ;
        RECT 44.450 -16.150 45.050 -16.100 ;
        RECT 35.150 -16.280 35.850 -16.250 ;
        RECT 60.540 -18.250 60.770 -17.250 ;
        RECT 63.710 -18.250 63.940 -17.250 ;
        RECT 68.960 -18.250 69.190 -17.250 ;
        RECT 35.010 -21.710 35.240 -20.710 ;
        RECT 55.400 -21.450 56.500 -20.350 ;
        RECT 29.800 -27.800 30.700 -27.000 ;
        RECT 24.210 -30.900 24.440 -28.700 ;
        RECT 26.790 -30.900 27.020 -28.700 ;
        RECT 29.370 -30.900 29.600 -28.700 ;
        RECT 31.950 -30.900 32.180 -28.700 ;
        RECT 34.530 -30.900 34.760 -28.700 ;
        RECT 37.110 -30.900 37.340 -28.700 ;
        RECT 38.720 -30.900 38.950 -29.900 ;
        RECT 44.570 -30.500 44.800 -28.790 ;
        RECT 47.150 -30.500 47.380 -28.790 ;
        RECT 55.560 -29.800 55.790 -28.800 ;
        RECT 58.560 -30.800 58.790 -28.800 ;
        RECT 64.420 -30.500 64.650 -28.790 ;
        RECT 67.000 -30.500 67.230 -28.790 ;
        RECT 75.410 -29.800 75.640 -28.800 ;
        RECT 78.410 -30.800 78.640 -28.800 ;
      LAYER via ;
        RECT 44.350 2.900 45.250 3.800 ;
        RECT 44.500 -16.100 45.000 -15.600 ;
        RECT 55.500 -21.350 56.400 -20.450 ;
        RECT 29.870 -27.780 30.630 -27.020 ;
      LAYER met2 ;
        RECT -57.500 9.000 -54.500 9.545 ;
        RECT -57.500 6.000 -47.970 9.000 ;
        RECT -57.500 5.500 -54.500 6.000 ;
        RECT 44.250 2.800 45.350 3.900 ;
        RECT 29.900 -16.250 35.880 -15.550 ;
        RECT 44.450 -16.150 45.050 -15.550 ;
        RECT 29.900 -27.000 30.600 -16.250 ;
        RECT 55.400 -21.450 56.500 -20.350 ;
        RECT 29.800 -27.800 30.700 -27.000 ;
      LAYER via2 ;
        RECT -57.500 6.500 -54.500 9.500 ;
        RECT 44.350 2.900 45.250 3.800 ;
        RECT 44.500 -16.100 45.000 -15.600 ;
        RECT 55.525 -21.325 56.375 -20.475 ;
      LAYER met3 ;
        RECT -57.525 64.505 -54.475 67.495 ;
        RECT -57.495 62.900 -54.505 64.505 ;
        RECT -57.500 9.525 -54.500 62.900 ;
        RECT -57.525 6.475 -54.475 9.525 ;
        RECT 44.250 2.800 45.350 3.900 ;
        RECT 44.350 -20.450 45.250 2.800 ;
        RECT 55.400 -20.450 56.500 -20.350 ;
        RECT 44.350 -21.350 56.500 -20.450 ;
        RECT 55.400 -21.450 56.500 -21.350 ;
      LAYER via3 ;
        RECT -57.495 64.505 -54.505 67.495 ;
      LAYER met4 ;
        RECT -58.000 64.000 83.000 68.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -24.700 23.700 -21.910 26.550 ;
        RECT -18.250 23.700 -15.460 26.550 ;
        RECT -11.800 23.700 -9.010 26.550 ;
        RECT -5.350 23.700 -2.560 26.550 ;
        RECT 1.100 23.700 3.890 26.550 ;
        RECT 7.550 23.700 10.340 26.550 ;
        RECT 14.000 23.700 16.790 26.550 ;
        RECT 20.450 23.700 23.240 26.550 ;
        RECT 26.900 23.700 29.690 26.550 ;
        RECT 33.350 23.700 36.140 26.550 ;
        RECT 39.800 23.700 42.590 26.550 ;
        RECT 46.250 23.700 49.040 26.550 ;
        RECT -24.700 20.500 -21.910 23.350 ;
        RECT -18.300 20.500 -15.510 23.350 ;
        RECT -11.800 20.500 -9.010 23.350 ;
        RECT -5.400 20.500 -2.610 23.350 ;
        RECT 1.100 20.500 3.890 23.350 ;
        RECT 7.500 20.500 10.290 23.350 ;
        RECT 14.000 20.500 16.790 23.350 ;
        RECT 20.400 20.500 23.190 23.350 ;
        RECT 26.900 20.500 29.690 23.350 ;
        RECT 33.300 20.500 36.090 23.350 ;
        RECT 39.800 20.500 42.590 23.350 ;
        RECT 46.200 20.500 48.990 23.350 ;
        RECT -1.400 12.000 4.250 14.790 ;
        RECT 18.700 7.850 20.810 10.640 ;
        RECT 21.100 7.850 26.060 10.640 ;
        RECT 26.350 7.850 31.310 10.640 ;
        RECT 31.600 7.850 36.510 10.640 ;
        RECT 36.800 7.850 41.760 10.640 ;
        RECT 42.050 7.850 44.900 10.640 ;
        RECT 45.170 7.850 47.280 10.640 ;
        RECT -20.000 3.400 -17.890 6.190 ;
        RECT -17.600 3.400 -12.690 6.190 ;
        RECT -12.400 3.400 -7.490 6.190 ;
        RECT -7.200 3.400 -2.290 6.190 ;
        RECT -2.000 3.400 0.850 6.190 ;
        RECT -13.600 -7.400 -11.140 -4.610 ;
        RECT -10.600 -7.400 -8.140 -4.610 ;
        RECT -17.000 -12.450 -2.430 -8.160 ;
        RECT 0.000 -9.600 2.850 -6.810 ;
        RECT 9.900 -7.400 12.360 -4.610 ;
        RECT 12.900 -7.400 15.360 -4.610 ;
        RECT 30.150 -7.400 32.610 -4.610 ;
        RECT 33.150 -7.400 35.610 -4.610 ;
        RECT 6.500 -12.450 21.070 -8.160 ;
        RECT 26.750 -12.450 41.320 -8.160 ;
        RECT -18.870 -28.530 15.050 -21.340 ;
        RECT 15.100 -24.200 18.060 -21.410 ;
        RECT 59.820 -22.150 61.930 -19.360 ;
        RECT 62.350 -22.150 64.460 -19.360 ;
        RECT 64.750 -22.150 69.710 -19.360 ;
        RECT 70.000 -22.150 72.850 -19.360 ;
        RECT 15.100 -28.600 18.060 -25.810 ;
        RECT 18.105 -28.595 21.065 -25.805 ;
        RECT -18.870 -35.930 15.050 -28.740 ;
        RECT 15.100 -31.600 18.060 -28.810 ;
        RECT 48.940 -30.900 51.400 -28.110 ;
        RECT 51.940 -30.900 54.400 -28.110 ;
        RECT 68.790 -30.900 71.250 -28.110 ;
        RECT 71.790 -30.900 74.250 -28.110 ;
        RECT 15.100 -36.000 18.060 -33.210 ;
        RECT 18.105 -35.995 21.065 -33.205 ;
        RECT 22.200 -33.210 38.060 -32.010 ;
        RECT 22.200 -36.000 40.960 -33.210 ;
        RECT 43.230 -35.910 57.800 -31.660 ;
        RECT 43.200 -35.950 57.800 -35.910 ;
        RECT 63.080 -35.950 77.650 -31.660 ;
        RECT 43.200 -38.700 48.900 -35.950 ;
      LAYER li1 ;
        RECT -24.520 26.200 -22.090 26.370 ;
        RECT -24.520 24.100 -24.350 26.200 ;
        RECT -22.260 24.100 -22.090 26.200 ;
        RECT -18.070 26.200 -15.640 26.370 ;
        RECT -18.070 24.100 -17.900 26.200 ;
        RECT -15.810 24.100 -15.640 26.200 ;
        RECT -11.620 26.200 -9.190 26.370 ;
        RECT -11.620 24.100 -11.450 26.200 ;
        RECT -9.360 24.100 -9.190 26.200 ;
        RECT -5.170 26.200 -2.740 26.370 ;
        RECT -5.170 24.100 -5.000 26.200 ;
        RECT -2.910 24.100 -2.740 26.200 ;
        RECT 1.280 26.200 3.710 26.370 ;
        RECT 1.280 24.100 1.450 26.200 ;
        RECT 3.540 24.100 3.710 26.200 ;
        RECT 7.730 26.200 10.160 26.370 ;
        RECT 7.730 24.100 7.900 26.200 ;
        RECT 9.990 24.100 10.160 26.200 ;
        RECT 14.180 26.200 16.610 26.370 ;
        RECT 14.180 24.100 14.350 26.200 ;
        RECT 16.440 24.100 16.610 26.200 ;
        RECT 20.630 26.200 23.060 26.370 ;
        RECT 20.630 24.100 20.800 26.200 ;
        RECT 22.890 24.100 23.060 26.200 ;
        RECT 27.080 26.200 29.510 26.370 ;
        RECT 27.080 24.100 27.250 26.200 ;
        RECT 29.340 24.100 29.510 26.200 ;
        RECT 33.530 26.200 35.960 26.370 ;
        RECT 33.530 24.100 33.700 26.200 ;
        RECT 35.790 24.100 35.960 26.200 ;
        RECT 39.980 26.200 42.410 26.370 ;
        RECT 39.980 24.100 40.150 26.200 ;
        RECT 42.240 24.100 42.410 26.200 ;
        RECT 46.430 26.200 48.860 26.370 ;
        RECT 46.430 24.100 46.600 26.200 ;
        RECT 48.690 24.100 48.860 26.200 ;
        RECT -24.700 23.700 49.100 24.100 ;
        RECT -24.700 23.170 -24.400 23.700 ;
        RECT -24.700 23.000 -22.090 23.170 ;
        RECT -24.700 20.900 -24.350 23.000 ;
        RECT -22.260 20.900 -22.090 23.000 ;
        RECT -18.120 23.000 -15.690 23.170 ;
        RECT -18.120 20.900 -17.950 23.000 ;
        RECT -15.860 20.900 -15.690 23.000 ;
        RECT -11.620 23.000 -9.190 23.170 ;
        RECT -11.620 20.900 -11.450 23.000 ;
        RECT -9.360 20.900 -9.190 23.000 ;
        RECT -5.220 23.000 -2.790 23.170 ;
        RECT -5.220 20.900 -5.050 23.000 ;
        RECT -2.960 20.900 -2.790 23.000 ;
        RECT 1.280 23.000 3.710 23.170 ;
        RECT 1.280 20.900 1.450 23.000 ;
        RECT 3.540 20.900 3.710 23.000 ;
        RECT 7.680 23.000 10.110 23.170 ;
        RECT 7.680 20.900 7.850 23.000 ;
        RECT 9.940 20.900 10.110 23.000 ;
        RECT 14.180 23.000 16.610 23.170 ;
        RECT 14.180 20.900 14.350 23.000 ;
        RECT 16.440 20.900 16.610 23.000 ;
        RECT 20.580 23.000 23.010 23.170 ;
        RECT 20.580 20.900 20.750 23.000 ;
        RECT 22.840 20.900 23.010 23.000 ;
        RECT 27.080 23.000 29.510 23.170 ;
        RECT 27.080 20.900 27.250 23.000 ;
        RECT 29.340 20.900 29.510 23.000 ;
        RECT 33.480 23.000 35.910 23.170 ;
        RECT 33.480 20.900 33.650 23.000 ;
        RECT 35.740 20.900 35.910 23.000 ;
        RECT 39.980 23.000 42.410 23.170 ;
        RECT 39.980 20.900 40.150 23.000 ;
        RECT 42.240 20.900 42.410 23.000 ;
        RECT 46.380 23.000 48.810 23.170 ;
        RECT 46.380 20.900 46.550 23.000 ;
        RECT 48.640 20.900 48.810 23.000 ;
        RECT -24.900 20.500 49.000 20.900 ;
        RECT -24.900 1.825 -24.000 20.500 ;
        RECT 1.100 14.610 1.800 20.500 ;
        RECT -1.220 14.440 4.070 14.610 ;
        RECT -1.220 12.350 -1.050 14.440 ;
        RECT 1.100 12.600 1.800 14.440 ;
        RECT 1.100 12.350 1.270 12.600 ;
        RECT -1.220 12.180 1.270 12.350 ;
        RECT 1.580 12.350 1.750 12.600 ;
        RECT 3.900 12.350 4.070 14.440 ;
        RECT 1.580 12.180 4.070 12.350 ;
        RECT 18.880 8.550 19.050 10.060 ;
        RECT 19.890 9.550 20.060 9.610 ;
        RECT 20.460 9.550 20.630 10.060 ;
        RECT 19.890 8.650 20.700 9.550 ;
        RECT 19.890 8.570 20.060 8.650 ;
        RECT 18.800 8.350 19.100 8.550 ;
        RECT 20.400 8.350 20.700 8.650 ;
        RECT 21.280 8.550 21.450 10.060 ;
        RECT 23.600 8.550 23.770 10.060 ;
        RECT 24.130 8.550 24.300 10.060 ;
        RECT 25.140 9.550 25.310 9.610 ;
        RECT 25.710 9.550 25.880 10.060 ;
        RECT 25.140 8.650 25.950 9.550 ;
        RECT 25.140 8.570 25.310 8.650 ;
        RECT 21.200 8.350 21.500 8.550 ;
        RECT 23.500 8.350 23.800 8.550 ;
        RECT 24.050 8.350 24.350 8.550 ;
        RECT 25.650 8.350 25.950 8.650 ;
        RECT 26.530 8.550 26.700 10.060 ;
        RECT 28.850 8.550 29.020 10.060 ;
        RECT 29.380 8.550 29.550 10.060 ;
        RECT 30.390 9.550 30.560 9.610 ;
        RECT 30.960 9.550 31.130 10.060 ;
        RECT 30.390 8.650 31.200 9.550 ;
        RECT 30.390 8.570 30.560 8.650 ;
        RECT 26.450 8.350 26.750 8.550 ;
        RECT 28.750 8.350 29.050 8.550 ;
        RECT 29.300 8.350 29.600 8.550 ;
        RECT 30.900 8.350 31.200 8.650 ;
        RECT 31.780 8.550 31.950 10.060 ;
        RECT 34.100 8.550 34.270 10.060 ;
        RECT 34.580 8.550 34.750 10.060 ;
        RECT 35.590 9.550 35.760 9.610 ;
        RECT 36.160 9.550 36.330 10.060 ;
        RECT 35.590 8.650 36.400 9.550 ;
        RECT 35.590 8.570 35.760 8.650 ;
        RECT 31.700 8.350 32.000 8.550 ;
        RECT 34.000 8.350 34.300 8.550 ;
        RECT 34.500 8.350 34.800 8.550 ;
        RECT 36.100 8.350 36.400 8.650 ;
        RECT 36.980 8.550 37.150 10.060 ;
        RECT 39.300 8.550 39.470 10.060 ;
        RECT 39.830 8.550 40.000 10.060 ;
        RECT 40.840 9.550 41.010 9.610 ;
        RECT 41.410 9.550 41.580 10.060 ;
        RECT 40.840 8.650 41.650 9.550 ;
        RECT 40.840 8.570 41.010 8.650 ;
        RECT 36.900 8.350 37.200 8.550 ;
        RECT 39.200 8.350 39.500 8.550 ;
        RECT 39.750 8.350 40.050 8.550 ;
        RECT 41.350 8.350 41.650 8.650 ;
        RECT 42.230 8.550 42.400 10.060 ;
        RECT 44.550 8.550 44.720 10.060 ;
        RECT 45.350 9.530 45.520 10.060 ;
        RECT 45.920 9.530 46.090 9.610 ;
        RECT 45.130 8.650 46.090 9.530 ;
        RECT 42.150 8.350 42.450 8.550 ;
        RECT 44.450 8.350 44.750 8.550 ;
        RECT 18.600 8.250 44.850 8.350 ;
        RECT 45.130 8.250 45.530 8.650 ;
        RECT 45.920 8.570 46.090 8.650 ;
        RECT 46.930 8.430 47.100 10.060 ;
        RECT 18.600 7.850 47.530 8.250 ;
        RECT -19.820 4.100 -19.650 5.610 ;
        RECT -18.810 5.100 -18.640 5.160 ;
        RECT -18.240 5.100 -18.070 5.610 ;
        RECT -18.810 4.200 -18.000 5.100 ;
        RECT -18.810 4.120 -18.640 4.200 ;
        RECT -19.900 3.900 -19.600 4.100 ;
        RECT -18.300 3.900 -18.000 4.200 ;
        RECT -17.420 4.100 -17.250 5.610 ;
        RECT -15.100 4.100 -14.930 5.610 ;
        RECT -14.620 4.100 -14.450 5.610 ;
        RECT -13.610 5.100 -13.440 5.160 ;
        RECT -13.040 5.100 -12.870 5.610 ;
        RECT -13.610 4.200 -12.800 5.100 ;
        RECT -13.610 4.120 -13.440 4.200 ;
        RECT -17.500 3.900 -17.200 4.100 ;
        RECT -15.200 3.900 -14.900 4.100 ;
        RECT -14.700 3.900 -14.400 4.100 ;
        RECT -13.100 3.900 -12.800 4.200 ;
        RECT -12.220 4.100 -12.050 5.610 ;
        RECT -9.900 4.100 -9.730 5.610 ;
        RECT -9.420 4.100 -9.250 5.610 ;
        RECT -8.410 5.100 -8.240 5.160 ;
        RECT -7.840 5.100 -7.670 5.610 ;
        RECT -8.410 4.200 -7.600 5.100 ;
        RECT -8.410 4.120 -8.240 4.200 ;
        RECT -12.300 3.900 -12.000 4.100 ;
        RECT -10.000 3.900 -9.700 4.100 ;
        RECT -9.500 3.900 -9.200 4.100 ;
        RECT -7.900 3.900 -7.600 4.200 ;
        RECT -7.020 4.100 -6.850 5.610 ;
        RECT -4.700 4.100 -4.530 5.610 ;
        RECT -4.220 4.100 -4.050 5.610 ;
        RECT -3.210 5.100 -3.040 5.160 ;
        RECT -2.640 5.100 -2.470 5.610 ;
        RECT -3.210 4.200 -2.400 5.100 ;
        RECT -3.210 4.120 -3.040 4.200 ;
        RECT -7.100 3.900 -6.800 4.100 ;
        RECT -4.800 3.900 -4.500 4.100 ;
        RECT -4.300 3.900 -4.000 4.100 ;
        RECT -2.700 3.900 -2.400 4.200 ;
        RECT -1.820 4.100 -1.650 5.610 ;
        RECT 0.500 4.100 0.670 5.610 ;
        RECT -1.900 3.900 -1.600 4.100 ;
        RECT 0.400 3.950 0.700 4.100 ;
        RECT 0.400 3.900 2.475 3.950 ;
        RECT -20.100 3.575 2.475 3.900 ;
        RECT -20.325 3.400 2.475 3.575 ;
        RECT -25.325 -11.925 -23.775 1.825 ;
        RECT -20.325 1.225 -18.775 3.400 ;
        RECT 0.450 3.300 1.000 3.400 ;
        RECT -13.420 -4.960 -11.320 -4.790 ;
        RECT -13.420 -7.050 -13.250 -4.960 ;
        RECT -12.060 -5.400 -11.890 -5.330 ;
        RECT -11.490 -5.400 -11.320 -4.960 ;
        RECT -10.420 -4.960 -8.320 -4.790 ;
        RECT -10.420 -5.400 -10.250 -4.960 ;
        RECT -9.850 -5.400 -9.680 -5.330 ;
        RECT -12.060 -6.360 -9.680 -5.400 ;
        RECT -12.060 -6.370 -10.250 -6.360 ;
        RECT -9.850 -6.370 -9.680 -6.360 ;
        RECT -11.900 -7.000 -10.250 -6.370 ;
        RECT -8.490 -7.000 -8.320 -4.960 ;
        RECT 10.080 -4.960 12.180 -4.790 ;
        RECT -13.050 -7.050 -8.320 -7.000 ;
        RECT -13.420 -7.220 -8.320 -7.050 ;
        RECT 0.180 -7.160 2.670 -6.990 ;
        RECT -13.050 -8.050 -8.350 -7.220 ;
        RECT -17.050 -8.340 -8.350 -8.050 ;
        RECT -17.050 -8.510 -2.610 -8.340 ;
        RECT -17.050 -8.600 -8.350 -8.510 ;
        RECT -17.050 -11.850 -16.550 -8.600 ;
        RECT -16.250 -10.950 -16.080 -9.190 ;
        RECT -13.670 -10.900 -13.500 -9.190 ;
        RECT -11.090 -10.900 -10.920 -9.190 ;
        RECT -8.510 -10.850 -8.340 -9.190 ;
        RECT -5.930 -10.800 -5.760 -9.190 ;
        RECT -16.350 -11.850 -16.050 -10.950 ;
        RECT -20.000 -11.925 -16.050 -11.850 ;
        RECT -25.325 -12.000 -16.050 -11.925 ;
        RECT -13.750 -12.000 -13.450 -10.900 ;
        RECT -11.150 -12.000 -10.850 -10.900 ;
        RECT -8.550 -12.000 -8.250 -10.850 ;
        RECT -6.000 -12.000 -5.700 -10.800 ;
        RECT -3.350 -10.850 -3.180 -9.190 ;
        RECT -3.400 -11.750 -3.100 -10.850 ;
        RECT -2.780 -11.750 -2.610 -8.510 ;
        RECT 0.180 -9.250 0.350 -7.160 ;
        RECT 2.500 -9.250 2.670 -7.160 ;
        RECT 10.080 -7.050 10.250 -4.960 ;
        RECT 11.440 -5.400 11.610 -5.330 ;
        RECT 12.010 -5.400 12.180 -4.960 ;
        RECT 13.080 -4.960 15.180 -4.790 ;
        RECT 13.080 -5.400 13.250 -4.960 ;
        RECT 13.650 -5.400 13.820 -5.330 ;
        RECT 11.440 -6.360 13.820 -5.400 ;
        RECT 11.440 -6.370 13.250 -6.360 ;
        RECT 13.650 -6.370 13.820 -6.360 ;
        RECT 11.600 -7.000 13.250 -6.370 ;
        RECT 15.010 -7.000 15.180 -4.960 ;
        RECT 10.450 -7.050 15.180 -7.000 ;
        RECT 10.080 -7.220 15.180 -7.050 ;
        RECT 30.330 -4.960 32.430 -4.790 ;
        RECT 30.330 -7.050 30.500 -4.960 ;
        RECT 31.690 -5.400 31.860 -5.330 ;
        RECT 32.260 -5.400 32.430 -4.960 ;
        RECT 33.330 -4.960 35.430 -4.790 ;
        RECT 33.330 -5.400 33.500 -4.960 ;
        RECT 33.900 -5.400 34.070 -5.330 ;
        RECT 31.690 -6.360 34.070 -5.400 ;
        RECT 31.690 -6.370 33.500 -6.360 ;
        RECT 33.900 -6.370 34.070 -6.360 ;
        RECT 31.850 -7.000 33.500 -6.370 ;
        RECT 35.260 -7.000 35.430 -4.960 ;
        RECT 30.700 -7.050 35.430 -7.000 ;
        RECT 30.330 -7.220 35.430 -7.050 ;
        RECT 10.450 -8.050 15.150 -7.220 ;
        RECT 30.700 -8.050 35.400 -7.220 ;
        RECT 0.180 -9.420 2.670 -9.250 ;
        RECT 6.450 -8.340 15.150 -8.050 ;
        RECT 26.700 -8.340 35.400 -8.050 ;
        RECT 6.450 -8.510 20.890 -8.340 ;
        RECT 6.450 -8.600 15.150 -8.510 ;
        RECT 1.300 -11.750 1.750 -9.420 ;
        RECT 6.450 -11.750 6.950 -8.600 ;
        RECT 7.250 -10.950 7.420 -9.190 ;
        RECT 9.830 -10.900 10.000 -9.190 ;
        RECT 12.410 -10.900 12.580 -9.190 ;
        RECT 14.990 -10.850 15.160 -9.190 ;
        RECT 17.570 -10.800 17.740 -9.190 ;
        RECT -3.400 -11.850 6.950 -11.750 ;
        RECT 7.150 -11.850 7.450 -10.950 ;
        RECT -3.400 -12.000 7.450 -11.850 ;
        RECT 9.750 -12.000 10.050 -10.900 ;
        RECT 12.350 -12.000 12.650 -10.900 ;
        RECT 14.950 -12.000 15.250 -10.850 ;
        RECT 17.500 -12.000 17.800 -10.800 ;
        RECT 20.150 -10.850 20.320 -9.190 ;
        RECT 20.100 -12.000 20.400 -10.850 ;
        RECT 20.720 -12.000 20.890 -8.510 ;
        RECT 26.700 -8.510 41.140 -8.340 ;
        RECT 26.700 -8.600 35.400 -8.510 ;
        RECT 26.700 -11.850 27.200 -8.600 ;
        RECT 27.500 -10.950 27.670 -9.190 ;
        RECT 30.080 -10.900 30.250 -9.190 ;
        RECT 32.660 -10.900 32.830 -9.190 ;
        RECT 35.240 -10.850 35.410 -9.190 ;
        RECT 37.820 -10.800 37.990 -9.190 ;
        RECT 27.400 -11.850 27.700 -10.950 ;
        RECT 23.750 -12.000 27.700 -11.850 ;
        RECT 30.000 -12.000 30.300 -10.900 ;
        RECT 32.600 -12.000 32.900 -10.900 ;
        RECT 35.200 -12.000 35.500 -10.850 ;
        RECT 37.750 -12.000 38.050 -10.800 ;
        RECT 40.400 -10.850 40.570 -9.190 ;
        RECT 40.350 -12.000 40.650 -10.850 ;
        RECT 40.970 -12.000 41.140 -8.510 ;
        RECT -25.325 -12.250 41.140 -12.000 ;
        RECT 42.850 -12.250 43.400 7.850 ;
        RECT -25.325 -12.700 43.500 -12.250 ;
        RECT -25.325 -13.300 47.700 -12.700 ;
        RECT -25.325 -13.350 43.500 -13.300 ;
        RECT -25.325 -13.475 -18.400 -13.350 ;
        RECT -19.950 -21.400 -18.400 -13.475 ;
        RECT 36.900 -19.450 37.500 -13.350 ;
        RECT 42.850 -13.400 43.400 -13.350 ;
        RECT -19.950 -21.800 18.000 -21.400 ;
        RECT -19.950 -28.000 -18.400 -21.800 ;
        RECT 14.700 -21.900 18.000 -21.800 ;
        RECT 36.900 -21.750 37.400 -19.450 ;
        RECT 38.100 -20.305 39.300 -20.250 ;
        RECT 38.100 -20.475 39.480 -20.305 ;
        RECT 60.000 -20.470 60.170 -19.940 ;
        RECT 60.570 -20.470 60.740 -20.390 ;
        RECT 38.100 -20.650 39.300 -20.475 ;
        RECT 14.700 -22.130 16.000 -21.900 ;
        RECT -18.120 -24.410 -17.950 -22.370 ;
        RECT -15.540 -24.410 -15.370 -22.370 ;
        RECT -12.960 -24.410 -12.790 -22.370 ;
        RECT -10.380 -24.410 -10.210 -22.370 ;
        RECT -7.800 -24.410 -7.630 -22.370 ;
        RECT -5.220 -24.410 -5.050 -22.370 ;
        RECT -2.640 -24.410 -2.470 -22.370 ;
        RECT -0.060 -24.410 0.110 -22.370 ;
        RECT 2.520 -24.410 2.690 -22.370 ;
        RECT 5.100 -24.410 5.270 -22.370 ;
        RECT 7.680 -24.410 7.850 -22.370 ;
        RECT 10.260 -24.410 10.430 -22.370 ;
        RECT 12.840 -24.410 13.010 -22.370 ;
        RECT 14.700 -23.100 16.020 -22.130 ;
        RECT -18.120 -27.500 -17.950 -25.460 ;
        RECT -15.540 -27.500 -15.370 -25.460 ;
        RECT -12.960 -27.500 -12.790 -25.460 ;
        RECT -10.380 -27.500 -10.210 -25.460 ;
        RECT -7.800 -27.500 -7.630 -25.460 ;
        RECT -5.220 -27.500 -5.050 -25.460 ;
        RECT -2.640 -27.500 -2.470 -25.460 ;
        RECT -0.060 -27.500 0.110 -25.460 ;
        RECT 2.520 -27.500 2.690 -25.460 ;
        RECT 5.100 -27.500 5.270 -25.460 ;
        RECT 7.680 -27.500 7.850 -25.460 ;
        RECT 10.260 -27.500 10.430 -25.460 ;
        RECT 12.840 -27.500 13.010 -25.460 ;
        RECT 14.700 -26.900 15.100 -23.100 ;
        RECT 15.280 -23.850 15.450 -23.100 ;
        RECT 15.850 -23.170 16.020 -23.100 ;
        RECT 17.710 -23.850 17.880 -21.900 ;
        RECT 36.900 -22.550 37.500 -21.750 ;
        RECT 38.100 -22.550 38.500 -20.650 ;
        RECT 59.780 -21.000 60.740 -20.470 ;
        RECT 57.700 -21.350 60.740 -21.000 ;
        RECT 57.700 -21.750 60.180 -21.350 ;
        RECT 60.570 -21.430 60.740 -21.350 ;
        RECT 61.580 -21.570 61.750 -19.940 ;
        RECT 62.530 -21.450 62.700 -19.940 ;
        RECT 63.540 -20.450 63.710 -20.390 ;
        RECT 64.110 -20.450 64.280 -19.940 ;
        RECT 63.540 -21.350 64.350 -20.450 ;
        RECT 63.540 -21.430 63.710 -21.350 ;
        RECT 62.450 -21.650 62.750 -21.450 ;
        RECT 64.050 -21.650 64.350 -21.350 ;
        RECT 64.930 -21.450 65.100 -19.940 ;
        RECT 67.250 -21.450 67.420 -19.940 ;
        RECT 67.780 -21.450 67.950 -19.940 ;
        RECT 68.790 -20.450 68.960 -20.390 ;
        RECT 69.360 -20.450 69.530 -19.940 ;
        RECT 68.790 -21.350 69.600 -20.450 ;
        RECT 68.790 -21.430 68.960 -21.350 ;
        RECT 64.850 -21.650 65.150 -21.450 ;
        RECT 67.150 -21.650 67.450 -21.450 ;
        RECT 67.700 -21.650 68.000 -21.450 ;
        RECT 69.300 -21.650 69.600 -21.350 ;
        RECT 70.180 -21.450 70.350 -19.940 ;
        RECT 72.500 -21.450 72.670 -19.940 ;
        RECT 70.100 -21.650 70.400 -21.450 ;
        RECT 72.400 -21.650 72.700 -21.450 ;
        RECT 62.250 -21.750 72.800 -21.650 ;
        RECT 57.700 -22.000 72.800 -21.750 ;
        RECT 59.700 -22.150 72.800 -22.000 ;
        RECT 36.900 -22.950 38.500 -22.550 ;
        RECT 36.900 -23.000 37.500 -22.950 ;
        RECT 15.280 -24.020 17.880 -23.850 ;
        RECT 15.280 -26.160 17.880 -25.990 ;
        RECT 15.280 -26.900 15.450 -26.160 ;
        RECT 15.850 -26.900 16.020 -26.840 ;
        RECT -20.000 -28.100 -18.400 -28.000 ;
        RECT 14.700 -27.800 16.020 -26.900 ;
        RECT 14.700 -28.100 15.100 -27.800 ;
        RECT 15.280 -28.100 15.450 -27.800 ;
        RECT 15.850 -27.880 16.020 -27.800 ;
        RECT 17.710 -28.100 17.880 -26.160 ;
        RECT 18.285 -26.155 20.885 -25.985 ;
        RECT 18.285 -27.000 18.455 -26.155 ;
        RECT 18.855 -27.000 19.025 -26.835 ;
        RECT 18.285 -27.800 19.100 -27.000 ;
        RECT 18.285 -28.100 18.455 -27.800 ;
        RECT 18.855 -27.875 19.025 -27.800 ;
        RECT 20.715 -28.100 20.885 -26.155 ;
        RECT -20.000 -28.500 21.100 -28.100 ;
        RECT 49.120 -28.460 51.220 -28.290 ;
        RECT -20.000 -29.000 21.000 -28.500 ;
        RECT -20.000 -29.200 18.000 -29.000 ;
        RECT -20.000 -35.500 -18.400 -29.200 ;
        RECT 14.700 -29.300 18.000 -29.200 ;
        RECT 14.700 -29.530 16.000 -29.300 ;
        RECT -18.120 -31.810 -17.950 -29.770 ;
        RECT -15.540 -31.810 -15.370 -29.770 ;
        RECT -12.960 -31.810 -12.790 -29.770 ;
        RECT -10.380 -31.810 -10.210 -29.770 ;
        RECT -7.800 -31.810 -7.630 -29.770 ;
        RECT -5.220 -31.810 -5.050 -29.770 ;
        RECT -2.640 -31.810 -2.470 -29.770 ;
        RECT -0.060 -31.810 0.110 -29.770 ;
        RECT 2.520 -31.810 2.690 -29.770 ;
        RECT 5.100 -31.810 5.270 -29.770 ;
        RECT 7.680 -31.810 7.850 -29.770 ;
        RECT 10.260 -31.810 10.430 -29.770 ;
        RECT 12.840 -31.810 13.010 -29.770 ;
        RECT 14.700 -30.500 16.020 -29.530 ;
        RECT -18.120 -34.900 -17.950 -32.860 ;
        RECT -15.540 -34.900 -15.370 -32.860 ;
        RECT -12.960 -34.900 -12.790 -32.860 ;
        RECT -10.380 -34.900 -10.210 -32.860 ;
        RECT -7.800 -34.900 -7.630 -32.860 ;
        RECT -5.220 -34.900 -5.050 -32.860 ;
        RECT -2.640 -34.900 -2.470 -32.860 ;
        RECT -0.060 -34.900 0.110 -32.860 ;
        RECT 2.520 -34.900 2.690 -32.860 ;
        RECT 5.100 -34.900 5.270 -32.860 ;
        RECT 7.680 -34.900 7.850 -32.860 ;
        RECT 10.260 -34.900 10.430 -32.860 ;
        RECT 12.840 -34.900 13.010 -32.860 ;
        RECT 14.700 -34.300 15.100 -30.500 ;
        RECT 15.280 -31.250 15.450 -30.500 ;
        RECT 15.850 -30.570 16.020 -30.500 ;
        RECT 17.710 -31.250 17.880 -29.300 ;
        RECT 49.120 -30.500 49.290 -28.460 ;
        RECT 50.480 -28.900 50.650 -28.830 ;
        RECT 51.050 -28.900 51.220 -28.460 ;
        RECT 52.120 -28.460 54.220 -28.290 ;
        RECT 52.120 -28.900 52.290 -28.460 ;
        RECT 52.690 -28.900 52.860 -28.830 ;
        RECT 50.480 -29.860 52.860 -28.900 ;
        RECT 50.480 -29.870 50.650 -29.860 ;
        RECT 51.050 -29.870 52.860 -29.860 ;
        RECT 51.050 -30.500 52.700 -29.870 ;
        RECT 49.120 -30.550 53.850 -30.500 ;
        RECT 54.050 -30.550 54.220 -28.460 ;
        RECT 49.120 -30.720 54.220 -30.550 ;
        RECT 68.970 -28.460 71.070 -28.290 ;
        RECT 68.970 -30.500 69.140 -28.460 ;
        RECT 70.330 -28.900 70.500 -28.830 ;
        RECT 70.900 -28.900 71.070 -28.460 ;
        RECT 71.970 -28.460 74.070 -28.290 ;
        RECT 71.970 -28.900 72.140 -28.460 ;
        RECT 72.540 -28.900 72.710 -28.830 ;
        RECT 70.330 -29.860 72.710 -28.900 ;
        RECT 70.330 -29.870 70.500 -29.860 ;
        RECT 70.900 -29.870 72.710 -29.860 ;
        RECT 70.900 -30.500 72.550 -29.870 ;
        RECT 68.970 -30.550 73.700 -30.500 ;
        RECT 73.900 -30.550 74.070 -28.460 ;
        RECT 68.970 -30.720 74.070 -30.550 ;
        RECT 15.280 -31.420 17.880 -31.250 ;
        RECT 49.150 -31.550 53.850 -30.720 ;
        RECT 69.000 -31.550 73.700 -30.720 ;
        RECT 49.150 -31.840 57.850 -31.550 ;
        RECT 69.000 -31.840 77.700 -31.550 ;
        RECT 43.410 -32.010 57.850 -31.840 ;
        RECT 22.380 -32.360 37.880 -32.190 ;
        RECT 15.280 -33.560 17.880 -33.390 ;
        RECT 15.280 -34.300 15.450 -33.560 ;
        RECT 15.850 -34.300 16.020 -34.240 ;
        RECT 14.700 -35.200 16.020 -34.300 ;
        RECT 14.700 -35.500 15.100 -35.200 ;
        RECT 15.280 -35.500 15.450 -35.200 ;
        RECT 15.850 -35.280 16.020 -35.200 ;
        RECT 17.710 -35.500 17.880 -33.560 ;
        RECT 18.285 -33.555 20.885 -33.385 ;
        RECT 18.285 -34.400 18.455 -33.555 ;
        RECT 18.855 -34.400 19.025 -34.235 ;
        RECT 18.285 -35.200 19.100 -34.400 ;
        RECT 18.285 -35.500 18.455 -35.200 ;
        RECT 18.855 -35.275 19.025 -35.200 ;
        RECT 20.715 -35.500 20.885 -33.555 ;
        RECT -20.000 -35.600 21.100 -35.500 ;
        RECT 22.380 -35.600 22.550 -32.360 ;
        RECT 22.950 -34.900 23.120 -33.040 ;
        RECT 25.530 -34.800 25.700 -33.040 ;
        RECT 28.110 -34.800 28.280 -33.040 ;
        RECT 30.690 -34.800 30.860 -33.040 ;
        RECT 33.270 -34.700 33.440 -33.040 ;
        RECT 35.850 -34.700 36.020 -33.040 ;
        RECT 22.900 -35.600 23.200 -34.900 ;
        RECT 25.500 -35.600 25.800 -34.800 ;
        RECT 28.000 -35.600 28.300 -34.800 ;
        RECT 30.600 -35.600 30.900 -34.800 ;
        RECT 33.200 -35.600 33.500 -34.700 ;
        RECT 35.800 -35.600 36.100 -34.700 ;
        RECT 37.710 -35.600 37.880 -32.360 ;
        RECT 38.180 -33.560 40.780 -33.390 ;
        RECT 38.180 -34.300 38.350 -33.560 ;
        RECT 38.750 -34.300 38.920 -34.240 ;
        RECT 38.180 -35.280 38.920 -34.300 ;
        RECT 38.180 -35.600 38.900 -35.280 ;
        RECT 40.610 -35.600 40.780 -33.560 ;
        RECT 43.410 -35.400 43.580 -32.010 ;
        RECT 49.150 -32.100 57.850 -32.010 ;
        RECT 43.980 -34.350 44.150 -32.690 ;
        RECT 46.560 -34.300 46.730 -32.690 ;
        RECT 43.200 -35.500 43.700 -35.400 ;
        RECT 43.900 -35.500 44.200 -34.350 ;
        RECT 46.500 -35.500 46.800 -34.300 ;
        RECT 49.140 -34.350 49.310 -32.690 ;
        RECT 49.050 -35.500 49.350 -34.350 ;
        RECT 51.720 -34.400 51.890 -32.690 ;
        RECT 54.300 -34.400 54.470 -32.690 ;
        RECT 51.650 -35.500 51.950 -34.400 ;
        RECT 54.250 -35.500 54.550 -34.400 ;
        RECT 56.880 -34.450 57.050 -32.690 ;
        RECT 56.850 -35.350 57.150 -34.450 ;
        RECT 57.350 -35.350 57.850 -32.100 ;
        RECT 63.260 -32.010 77.700 -31.840 ;
        RECT 63.260 -35.350 63.430 -32.010 ;
        RECT 69.000 -32.100 77.700 -32.010 ;
        RECT 63.830 -34.350 64.000 -32.690 ;
        RECT 66.410 -34.300 66.580 -32.690 ;
        RECT 63.750 -35.350 64.050 -34.350 ;
        RECT 56.850 -35.500 64.050 -35.350 ;
        RECT 66.350 -35.500 66.650 -34.300 ;
        RECT 68.990 -34.350 69.160 -32.690 ;
        RECT 68.900 -35.500 69.200 -34.350 ;
        RECT 71.570 -34.400 71.740 -32.690 ;
        RECT 74.150 -34.400 74.320 -32.690 ;
        RECT 71.500 -35.500 71.800 -34.400 ;
        RECT 74.100 -35.500 74.400 -34.400 ;
        RECT 76.730 -34.450 76.900 -32.690 ;
        RECT 76.700 -35.350 77.000 -34.450 ;
        RECT 77.200 -35.350 77.700 -32.100 ;
        RECT 76.700 -35.500 80.650 -35.350 ;
        RECT 43.200 -35.600 80.650 -35.500 ;
        RECT -20.000 -36.000 80.650 -35.600 ;
        RECT -20.000 -36.200 77.700 -36.000 ;
        RECT -20.000 -36.500 43.200 -36.200 ;
        RECT 43.380 -36.260 45.870 -36.200 ;
        RECT 43.380 -38.350 43.550 -36.260 ;
        RECT 45.700 -38.350 45.870 -36.260 ;
        RECT 43.380 -38.520 45.870 -38.350 ;
        RECT 46.230 -36.260 48.720 -36.200 ;
        RECT 46.230 -38.350 46.400 -36.260 ;
        RECT 48.550 -38.350 48.720 -36.260 ;
        RECT 48.900 -36.550 77.700 -36.200 ;
        RECT 58.000 -37.625 58.750 -36.550 ;
        RECT 46.230 -38.520 48.720 -38.350 ;
      LAYER mcon ;
        RECT 45.920 8.650 46.090 9.530 ;
        RECT 1.925 3.400 2.475 3.950 ;
        RECT -25.325 0.275 -23.775 1.825 ;
        RECT -20.295 1.255 -18.805 2.745 ;
        RECT -12.060 -6.290 -11.890 -5.410 ;
        RECT -9.850 -6.290 -9.680 -5.410 ;
        RECT -16.250 -11.650 -16.080 -9.270 ;
        RECT -13.670 -11.650 -13.500 -9.270 ;
        RECT -11.090 -11.650 -10.920 -9.270 ;
        RECT -8.510 -11.650 -8.340 -9.270 ;
        RECT -5.930 -11.650 -5.760 -9.270 ;
        RECT -3.350 -11.650 -3.180 -9.270 ;
        RECT 11.440 -6.290 11.610 -5.410 ;
        RECT 13.650 -6.290 13.820 -5.410 ;
        RECT 31.690 -6.290 31.860 -5.410 ;
        RECT 33.900 -6.290 34.070 -5.410 ;
        RECT 7.250 -11.650 7.420 -9.270 ;
        RECT 9.830 -11.650 10.000 -9.270 ;
        RECT 12.410 -11.650 12.580 -9.270 ;
        RECT 14.990 -11.650 15.160 -9.270 ;
        RECT 17.570 -11.650 17.740 -9.270 ;
        RECT 20.150 -11.650 20.320 -9.270 ;
        RECT 27.500 -11.650 27.670 -9.270 ;
        RECT 30.080 -11.650 30.250 -9.270 ;
        RECT 32.660 -11.650 32.830 -9.270 ;
        RECT 35.240 -11.650 35.410 -9.270 ;
        RECT 37.820 -11.650 37.990 -9.270 ;
        RECT 40.400 -11.650 40.570 -9.270 ;
        RECT 47.100 -13.300 47.700 -12.700 ;
        RECT -18.100 -21.700 14.600 -21.500 ;
        RECT 38.250 -21.650 38.420 -20.770 ;
        RECT -18.120 -24.330 -17.950 -22.450 ;
        RECT -15.540 -24.330 -15.370 -22.450 ;
        RECT -12.960 -24.330 -12.790 -22.450 ;
        RECT -10.380 -24.330 -10.210 -22.450 ;
        RECT -7.800 -24.330 -7.630 -22.450 ;
        RECT -5.220 -24.330 -5.050 -22.450 ;
        RECT -2.640 -24.330 -2.470 -22.450 ;
        RECT -0.060 -24.330 0.110 -22.450 ;
        RECT 2.520 -24.330 2.690 -22.450 ;
        RECT 5.100 -24.330 5.270 -22.450 ;
        RECT 7.680 -24.330 7.850 -22.450 ;
        RECT 10.260 -24.330 10.430 -22.450 ;
        RECT 12.840 -24.330 13.010 -22.450 ;
        RECT 15.850 -23.090 16.020 -22.210 ;
        RECT -18.120 -27.420 -17.950 -25.540 ;
        RECT -15.540 -27.420 -15.370 -25.540 ;
        RECT -12.960 -27.420 -12.790 -25.540 ;
        RECT -10.380 -27.420 -10.210 -25.540 ;
        RECT -7.800 -27.420 -7.630 -25.540 ;
        RECT -5.220 -27.420 -5.050 -25.540 ;
        RECT -2.640 -27.420 -2.470 -25.540 ;
        RECT -0.060 -27.420 0.110 -25.540 ;
        RECT 2.520 -27.420 2.690 -25.540 ;
        RECT 5.100 -27.420 5.270 -25.540 ;
        RECT 7.680 -27.420 7.850 -25.540 ;
        RECT 10.260 -27.420 10.430 -25.540 ;
        RECT 12.840 -27.420 13.010 -25.540 ;
        RECT 57.830 -21.570 58.370 -21.030 ;
        RECT 60.570 -21.350 60.740 -20.470 ;
        RECT 15.850 -27.800 16.020 -26.920 ;
        RECT 18.855 -27.795 19.025 -26.915 ;
        RECT -18.000 -28.400 14.600 -28.200 ;
        RECT -18.100 -29.100 14.600 -28.900 ;
        RECT -18.120 -31.730 -17.950 -29.850 ;
        RECT -15.540 -31.730 -15.370 -29.850 ;
        RECT -12.960 -31.730 -12.790 -29.850 ;
        RECT -10.380 -31.730 -10.210 -29.850 ;
        RECT -7.800 -31.730 -7.630 -29.850 ;
        RECT -5.220 -31.730 -5.050 -29.850 ;
        RECT -2.640 -31.730 -2.470 -29.850 ;
        RECT -0.060 -31.730 0.110 -29.850 ;
        RECT 2.520 -31.730 2.690 -29.850 ;
        RECT 5.100 -31.730 5.270 -29.850 ;
        RECT 7.680 -31.730 7.850 -29.850 ;
        RECT 10.260 -31.730 10.430 -29.850 ;
        RECT 12.840 -31.730 13.010 -29.850 ;
        RECT 15.850 -30.490 16.020 -29.610 ;
        RECT -18.120 -34.820 -17.950 -32.940 ;
        RECT -15.540 -34.820 -15.370 -32.940 ;
        RECT -12.960 -34.820 -12.790 -32.940 ;
        RECT -10.380 -34.820 -10.210 -32.940 ;
        RECT -7.800 -34.820 -7.630 -32.940 ;
        RECT -5.220 -34.820 -5.050 -32.940 ;
        RECT -2.640 -34.820 -2.470 -32.940 ;
        RECT -0.060 -34.820 0.110 -32.940 ;
        RECT 2.520 -34.820 2.690 -32.940 ;
        RECT 5.100 -34.820 5.270 -32.940 ;
        RECT 7.680 -34.820 7.850 -32.940 ;
        RECT 10.260 -34.820 10.430 -32.940 ;
        RECT 12.840 -34.820 13.010 -32.940 ;
        RECT 50.480 -29.790 50.650 -28.910 ;
        RECT 52.690 -29.790 52.860 -28.910 ;
        RECT 70.330 -29.790 70.500 -28.910 ;
        RECT 72.540 -29.790 72.710 -28.910 ;
        RECT 15.850 -35.200 16.020 -34.320 ;
        RECT 18.855 -35.195 19.025 -34.315 ;
        RECT 22.950 -35.200 23.120 -33.120 ;
        RECT 25.530 -35.200 25.700 -33.120 ;
        RECT 28.110 -35.200 28.280 -33.120 ;
        RECT 30.690 -35.200 30.860 -33.120 ;
        RECT 33.270 -35.200 33.440 -33.120 ;
        RECT 35.850 -35.200 36.020 -33.120 ;
        RECT 38.750 -35.200 38.920 -34.320 ;
        RECT 43.980 -35.150 44.150 -32.770 ;
        RECT 46.560 -35.150 46.730 -32.770 ;
        RECT 49.140 -35.150 49.310 -32.770 ;
        RECT 51.720 -35.150 51.890 -32.770 ;
        RECT 54.300 -35.150 54.470 -32.770 ;
        RECT 56.880 -35.150 57.050 -32.770 ;
        RECT 63.830 -35.150 64.000 -32.770 ;
        RECT 66.410 -35.150 66.580 -32.770 ;
        RECT 68.990 -35.150 69.160 -32.770 ;
        RECT 71.570 -35.150 71.740 -32.770 ;
        RECT 74.150 -35.150 74.320 -32.770 ;
        RECT 76.730 -35.150 76.900 -32.770 ;
        RECT -18.000 -35.800 14.600 -35.600 ;
        RECT 58.030 -37.595 58.720 -36.905 ;
      LAYER met1 ;
        RECT 19.860 8.590 20.090 9.590 ;
        RECT 25.110 8.590 25.340 9.590 ;
        RECT 30.360 8.590 30.590 9.590 ;
        RECT 35.560 8.590 35.790 9.590 ;
        RECT 40.810 8.590 41.040 9.590 ;
        RECT 45.890 8.590 46.120 9.590 ;
        RECT -18.840 4.140 -18.610 5.140 ;
        RECT -13.640 4.140 -13.410 5.140 ;
        RECT -8.440 4.140 -8.210 5.140 ;
        RECT -3.240 4.140 -3.010 5.140 ;
        RECT 1.895 3.340 2.505 4.010 ;
        RECT -51.125 2.625 -47.875 2.655 ;
        RECT -26.500 2.625 -20.700 2.700 ;
        RECT -51.125 2.000 -20.700 2.625 ;
        RECT -20.325 2.000 -18.775 2.805 ;
        RECT -51.125 0.250 -18.750 2.000 ;
        RECT -51.125 -0.600 -20.700 0.250 ;
        RECT -51.125 -0.625 -26.375 -0.600 ;
        RECT -51.125 -0.655 -47.875 -0.625 ;
        RECT -12.090 -6.350 -11.860 -5.350 ;
        RECT -9.880 -6.350 -9.650 -5.350 ;
        RECT 11.410 -6.350 11.640 -5.350 ;
        RECT 13.620 -6.350 13.850 -5.350 ;
        RECT 31.660 -6.350 31.890 -5.350 ;
        RECT 33.870 -6.350 34.100 -5.350 ;
        RECT -16.280 -11.710 -16.050 -9.210 ;
        RECT -13.700 -11.710 -13.470 -9.210 ;
        RECT -11.120 -11.710 -10.890 -9.210 ;
        RECT -8.540 -11.710 -8.310 -9.210 ;
        RECT -5.960 -11.710 -5.730 -9.210 ;
        RECT -3.380 -11.710 -3.150 -9.210 ;
        RECT 7.220 -11.710 7.450 -9.210 ;
        RECT 9.800 -11.710 10.030 -9.210 ;
        RECT 12.380 -11.710 12.610 -9.210 ;
        RECT 14.960 -11.710 15.190 -9.210 ;
        RECT 17.540 -11.710 17.770 -9.210 ;
        RECT 20.120 -11.710 20.350 -9.210 ;
        RECT 27.470 -11.710 27.700 -9.210 ;
        RECT 30.050 -11.710 30.280 -9.210 ;
        RECT 32.630 -11.710 32.860 -9.210 ;
        RECT 35.210 -11.710 35.440 -9.210 ;
        RECT 37.790 -11.710 38.020 -9.210 ;
        RECT 40.370 -11.710 40.600 -9.210 ;
        RECT 47.000 -13.400 47.800 -12.600 ;
        RECT -18.200 -21.800 14.800 -21.400 ;
        RECT 38.220 -21.710 38.450 -20.710 ;
        RECT 57.700 -21.700 58.500 -21.000 ;
        RECT 60.540 -21.410 60.770 -20.410 ;
        RECT 63.510 -21.410 63.740 -20.410 ;
        RECT 68.760 -21.410 68.990 -20.410 ;
        RECT -18.200 -22.600 -17.900 -21.800 ;
        RECT -15.600 -22.600 -15.300 -21.800 ;
        RECT -13.000 -22.600 -12.700 -21.800 ;
        RECT -10.400 -22.390 -10.100 -21.800 ;
        RECT -10.410 -22.600 -10.100 -22.390 ;
        RECT -7.900 -22.600 -7.600 -21.800 ;
        RECT -5.300 -22.600 -5.000 -21.800 ;
        RECT -2.700 -22.600 -2.400 -21.800 ;
        RECT -0.100 -22.600 0.200 -21.800 ;
        RECT 2.400 -22.390 2.700 -21.800 ;
        RECT 2.400 -22.600 2.720 -22.390 ;
        RECT 5.000 -22.600 5.300 -21.800 ;
        RECT 7.600 -22.600 7.900 -21.800 ;
        RECT 10.200 -22.600 10.500 -21.800 ;
        RECT 12.800 -22.600 13.100 -21.800 ;
        RECT -18.150 -24.390 -17.920 -22.600 ;
        RECT -15.570 -24.390 -15.340 -22.600 ;
        RECT -12.990 -24.390 -12.760 -22.600 ;
        RECT -10.410 -24.390 -10.180 -22.600 ;
        RECT -7.830 -24.390 -7.600 -22.600 ;
        RECT -5.250 -24.390 -5.020 -22.600 ;
        RECT -2.670 -24.390 -2.440 -22.600 ;
        RECT -0.090 -24.390 0.140 -22.600 ;
        RECT 2.490 -24.390 2.720 -22.600 ;
        RECT 5.070 -24.390 5.300 -22.600 ;
        RECT 7.650 -24.390 7.880 -22.600 ;
        RECT 10.230 -24.390 10.460 -22.600 ;
        RECT 12.810 -24.390 13.040 -22.600 ;
        RECT 15.820 -23.150 16.050 -22.150 ;
        RECT -18.150 -26.800 -17.920 -25.480 ;
        RECT -18.200 -28.100 -17.900 -26.800 ;
        RECT -15.570 -26.900 -15.340 -25.480 ;
        RECT -12.990 -26.800 -12.760 -25.480 ;
        RECT -15.600 -28.100 -15.300 -26.900 ;
        RECT -13.000 -28.100 -12.700 -26.800 ;
        RECT -10.410 -26.900 -10.180 -25.480 ;
        RECT -7.830 -26.900 -7.600 -25.480 ;
        RECT -5.250 -26.900 -5.020 -25.480 ;
        RECT -2.670 -26.900 -2.440 -25.480 ;
        RECT -0.090 -26.900 0.140 -25.480 ;
        RECT 2.490 -26.900 2.720 -25.480 ;
        RECT 5.070 -26.900 5.300 -25.480 ;
        RECT 7.650 -26.900 7.880 -25.480 ;
        RECT 10.230 -26.900 10.460 -25.480 ;
        RECT 12.810 -26.900 13.040 -25.480 ;
        RECT -10.500 -27.480 -10.180 -26.900 ;
        RECT -10.500 -28.100 -10.200 -27.480 ;
        RECT -7.900 -28.100 -7.600 -26.900 ;
        RECT -5.300 -28.100 -5.000 -26.900 ;
        RECT -2.700 -28.100 -2.400 -26.900 ;
        RECT -0.100 -28.100 0.200 -26.900 ;
        RECT 2.400 -27.480 2.720 -26.900 ;
        RECT 2.400 -28.100 2.700 -27.480 ;
        RECT 5.000 -28.100 5.300 -26.900 ;
        RECT 7.600 -28.100 7.900 -26.900 ;
        RECT 10.200 -28.100 10.500 -26.900 ;
        RECT 12.800 -28.100 13.100 -26.900 ;
        RECT 15.820 -27.860 16.050 -26.860 ;
        RECT 18.825 -27.855 19.055 -26.855 ;
        RECT -18.200 -28.500 14.800 -28.100 ;
        RECT -18.200 -29.200 14.800 -28.800 ;
        RECT -18.200 -30.000 -17.900 -29.200 ;
        RECT -15.600 -30.000 -15.300 -29.200 ;
        RECT -13.000 -30.000 -12.700 -29.200 ;
        RECT -10.400 -29.790 -10.100 -29.200 ;
        RECT -10.410 -30.000 -10.100 -29.790 ;
        RECT -7.900 -30.000 -7.600 -29.200 ;
        RECT -5.300 -30.000 -5.000 -29.200 ;
        RECT -2.700 -30.000 -2.400 -29.200 ;
        RECT -0.100 -30.000 0.200 -29.200 ;
        RECT 2.400 -29.790 2.700 -29.200 ;
        RECT 2.400 -30.000 2.720 -29.790 ;
        RECT 5.000 -30.000 5.300 -29.200 ;
        RECT 7.600 -30.000 7.900 -29.200 ;
        RECT 10.200 -30.000 10.500 -29.200 ;
        RECT 12.800 -30.000 13.100 -29.200 ;
        RECT -18.150 -31.790 -17.920 -30.000 ;
        RECT -15.570 -31.790 -15.340 -30.000 ;
        RECT -12.990 -31.790 -12.760 -30.000 ;
        RECT -10.410 -31.790 -10.180 -30.000 ;
        RECT -7.830 -31.790 -7.600 -30.000 ;
        RECT -5.250 -31.790 -5.020 -30.000 ;
        RECT -2.670 -31.790 -2.440 -30.000 ;
        RECT -0.090 -31.790 0.140 -30.000 ;
        RECT 2.490 -31.790 2.720 -30.000 ;
        RECT 5.070 -31.790 5.300 -30.000 ;
        RECT 7.650 -31.790 7.880 -30.000 ;
        RECT 10.230 -31.790 10.460 -30.000 ;
        RECT 12.810 -31.790 13.040 -30.000 ;
        RECT 15.820 -30.550 16.050 -29.550 ;
        RECT 50.450 -29.850 50.680 -28.850 ;
        RECT 52.660 -29.850 52.890 -28.850 ;
        RECT 70.300 -29.850 70.530 -28.850 ;
        RECT 72.510 -29.850 72.740 -28.850 ;
        RECT -18.150 -34.200 -17.920 -32.880 ;
        RECT -18.200 -35.500 -17.900 -34.200 ;
        RECT -15.570 -34.300 -15.340 -32.880 ;
        RECT -12.990 -34.200 -12.760 -32.880 ;
        RECT -15.600 -35.500 -15.300 -34.300 ;
        RECT -13.000 -35.500 -12.700 -34.200 ;
        RECT -10.410 -34.300 -10.180 -32.880 ;
        RECT -7.830 -34.300 -7.600 -32.880 ;
        RECT -5.250 -34.300 -5.020 -32.880 ;
        RECT -2.670 -34.300 -2.440 -32.880 ;
        RECT -0.090 -34.300 0.140 -32.880 ;
        RECT 2.490 -34.300 2.720 -32.880 ;
        RECT 5.070 -34.300 5.300 -32.880 ;
        RECT 7.650 -34.300 7.880 -32.880 ;
        RECT 10.230 -34.300 10.460 -32.880 ;
        RECT 12.810 -34.300 13.040 -32.880 ;
        RECT -10.500 -34.880 -10.180 -34.300 ;
        RECT -10.500 -35.500 -10.200 -34.880 ;
        RECT -7.900 -35.500 -7.600 -34.300 ;
        RECT -5.300 -35.500 -5.000 -34.300 ;
        RECT -2.700 -35.500 -2.400 -34.300 ;
        RECT -0.100 -35.500 0.200 -34.300 ;
        RECT 2.400 -34.880 2.720 -34.300 ;
        RECT 2.400 -35.500 2.700 -34.880 ;
        RECT 5.000 -35.500 5.300 -34.300 ;
        RECT 7.600 -35.500 7.900 -34.300 ;
        RECT 10.200 -35.500 10.500 -34.300 ;
        RECT 12.800 -35.500 13.100 -34.300 ;
        RECT 15.820 -35.260 16.050 -34.260 ;
        RECT 18.825 -35.255 19.055 -34.255 ;
        RECT 22.920 -35.260 23.150 -33.060 ;
        RECT 25.500 -35.260 25.730 -33.060 ;
        RECT 28.080 -35.260 28.310 -33.060 ;
        RECT 30.660 -35.260 30.890 -33.060 ;
        RECT 33.240 -35.260 33.470 -33.060 ;
        RECT 35.820 -35.260 36.050 -33.060 ;
        RECT 38.720 -35.260 38.950 -34.260 ;
        RECT 43.950 -35.210 44.180 -32.710 ;
        RECT 46.530 -35.210 46.760 -32.710 ;
        RECT 49.110 -35.210 49.340 -32.710 ;
        RECT 51.690 -35.210 51.920 -32.710 ;
        RECT 54.270 -35.210 54.500 -32.710 ;
        RECT 56.850 -35.210 57.080 -32.710 ;
        RECT 63.800 -35.210 64.030 -32.710 ;
        RECT 66.380 -35.210 66.610 -32.710 ;
        RECT 68.960 -35.210 69.190 -32.710 ;
        RECT 71.540 -35.210 71.770 -32.710 ;
        RECT 74.120 -35.210 74.350 -32.710 ;
        RECT 76.700 -35.210 76.930 -32.710 ;
        RECT -18.200 -35.900 14.800 -35.500 ;
        RECT 57.900 -37.700 58.850 -36.800 ;
      LAYER via ;
        RECT 1.895 3.370 2.505 3.980 ;
        RECT 47.070 -13.330 47.730 -12.670 ;
        RECT 57.800 -21.600 58.370 -21.000 ;
        RECT 58.000 -37.625 58.750 -36.875 ;
      LAYER met2 ;
        RECT 1.800 3.300 2.600 4.050 ;
        RECT -62.500 2.500 -59.500 2.545 ;
        RECT -57.500 2.500 -54.500 3.000 ;
        RECT -51.500 2.500 -47.845 2.625 ;
        RECT -63.000 -0.500 -47.845 2.500 ;
        RECT -62.500 -0.545 -59.500 -0.500 ;
        RECT -57.500 -1.000 -54.500 -0.500 ;
        RECT -51.500 -0.625 -47.845 -0.500 ;
        RECT 47.000 -12.700 47.800 -12.600 ;
        RECT 47.000 -13.300 58.400 -12.700 ;
        RECT 47.000 -13.400 47.800 -13.300 ;
        RECT 57.800 -21.000 58.400 -13.300 ;
        RECT 57.700 -21.700 58.500 -21.000 ;
        RECT 57.900 -37.700 58.850 -36.800 ;
      LAYER via2 ;
        RECT 1.895 3.370 2.505 3.980 ;
        RECT -62.500 -0.500 -59.500 2.500 ;
        RECT 58.025 -37.600 58.725 -36.900 ;
      LAYER met3 ;
        RECT -62.550 86.475 -59.440 89.525 ;
        RECT -62.515 2.525 -59.480 86.475 ;
        RECT 1.870 3.345 2.560 4.005 ;
        RECT -62.525 -0.525 -59.475 2.525 ;
        RECT 57.900 -37.700 58.850 -36.800 ;
        RECT 48.950 -52.100 58.445 -43.100 ;
      LAYER via3 ;
        RECT -62.520 86.475 -59.470 89.525 ;
        RECT 1.980 3.345 2.530 4.005 ;
        RECT 58.005 -37.620 58.745 -36.880 ;
        RECT 58.025 -51.960 58.345 -43.240 ;
      LAYER met4 ;
        RECT -65.000 86.000 83.000 90.000 ;
        RECT 1.975 3.950 2.535 4.010 ;
        RECT 3.795 3.950 11.405 9.450 ;
        RECT 1.975 3.400 11.405 3.950 ;
        RECT 1.975 3.340 2.535 3.400 ;
        RECT 3.795 1.840 11.405 3.400 ;
        RECT 57.900 -37.700 58.850 -36.800 ;
        RECT 58.000 -43.160 58.450 -37.700 ;
        RECT 57.945 -43.750 58.450 -43.160 ;
        RECT 57.945 -52.040 58.425 -43.750 ;
    END
  END VSS
  PIN PD1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT -23.670 25.630 -22.630 25.800 ;
        RECT -21.800 25.550 -21.500 26.000 ;
        RECT -21.700 24.750 -21.500 25.550 ;
        RECT -23.670 24.450 -22.630 24.620 ;
        RECT -21.750 24.300 -21.450 24.750 ;
        RECT -23.670 22.430 -22.630 22.600 ;
        RECT -23.670 21.250 -22.630 21.420 ;
      LAYER mcon ;
        RECT -23.590 25.630 -22.710 25.800 ;
        RECT -21.750 25.650 -21.550 25.900 ;
        RECT -23.590 24.450 -22.710 24.620 ;
        RECT -21.700 24.400 -21.500 24.650 ;
        RECT -23.590 22.430 -22.710 22.600 ;
        RECT -23.590 21.250 -22.710 21.420 ;
      LAYER met1 ;
        RECT -22.430 25.900 -22.170 25.935 ;
        RECT -21.800 25.900 -21.500 26.000 ;
        RECT -23.150 25.830 -21.500 25.900 ;
        RECT -23.650 25.650 -21.500 25.830 ;
        RECT -23.650 25.600 -22.650 25.650 ;
        RECT -22.430 25.615 -22.170 25.650 ;
        RECT -21.800 25.550 -21.500 25.650 ;
        RECT -21.750 24.650 -21.450 24.750 ;
        RECT -23.650 24.420 -21.450 24.650 ;
        RECT -23.150 24.400 -21.450 24.420 ;
        RECT -22.325 22.700 -22.075 24.400 ;
        RECT -21.750 24.300 -21.450 24.400 ;
        RECT -23.050 22.630 -20.750 22.700 ;
        RECT -23.650 22.450 -20.750 22.630 ;
        RECT -23.650 22.400 -22.650 22.450 ;
        RECT -23.650 21.400 -22.650 21.450 ;
        RECT -21.000 21.400 -20.750 22.450 ;
        RECT -23.650 21.220 -20.750 21.400 ;
        RECT -23.100 21.150 -20.750 21.220 ;
      LAYER via ;
        RECT -22.430 25.645 -22.170 25.905 ;
      LAYER met2 ;
        RECT -40.000 38.400 -39.400 42.450 ;
        RECT -39.830 35.020 -39.530 38.400 ;
        RECT -39.865 34.740 -39.495 35.020 ;
        RECT -39.830 34.730 -39.530 34.740 ;
        RECT -22.450 25.905 -22.150 26.295 ;
        RECT -22.460 25.645 -22.140 25.905 ;
      LAYER via2 ;
        RECT -39.820 34.740 -39.540 35.020 ;
        RECT -22.450 25.950 -22.150 26.250 ;
      LAYER met3 ;
        RECT -39.845 35.030 -39.515 35.045 ;
        RECT -39.845 34.730 -22.150 35.030 ;
        RECT -39.845 34.715 -39.515 34.730 ;
        RECT -22.450 26.275 -22.150 34.730 ;
        RECT -22.475 25.925 -22.125 26.275 ;
    END
  END PD1
  PIN pd1_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT -24.150 22.385 -23.850 22.450 ;
        RECT -24.150 22.055 -23.840 22.385 ;
        RECT -24.150 21.795 -23.850 22.055 ;
        RECT -24.150 21.465 -23.840 21.795 ;
        RECT -24.150 21.450 -23.850 21.465 ;
      LAYER mcon ;
        RECT -24.100 21.600 -23.900 22.300 ;
      LAYER met1 ;
        RECT -24.150 22.050 -23.850 22.450 ;
        RECT -26.250 21.750 -23.850 22.050 ;
        RECT -26.250 19.450 -25.950 21.750 ;
        RECT -24.150 21.450 -23.850 21.750 ;
        RECT -26.280 19.150 -25.920 19.450 ;
      LAYER via ;
        RECT -26.250 19.150 -25.950 19.450 ;
      LAYER met2 ;
        RECT -26.250 -41.850 -25.950 19.480 ;
        RECT -26.250 -42.150 4.950 -41.850 ;
        RECT 4.650 -64.350 4.950 -42.150 ;
        RECT 4.650 -64.650 20.450 -64.350 ;
        RECT 20.150 -68.350 20.450 -64.650 ;
        RECT 20.000 -72.350 20.600 -68.350 ;
    END
  END pd1_a
  PIN pd1_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT -24.150 25.585 -23.850 25.650 ;
        RECT -24.150 25.255 -23.840 25.585 ;
        RECT -24.150 24.995 -23.850 25.255 ;
        RECT -24.150 24.665 -23.840 24.995 ;
        RECT -24.150 24.650 -23.850 24.665 ;
      LAYER mcon ;
        RECT -24.100 24.800 -23.900 25.500 ;
      LAYER met1 ;
        RECT -26.250 25.250 -25.950 25.280 ;
        RECT -24.150 25.250 -23.850 25.650 ;
        RECT -26.250 24.950 -23.850 25.250 ;
        RECT -26.250 24.920 -25.950 24.950 ;
        RECT -24.150 24.650 -23.850 24.950 ;
      LAYER met2 ;
        RECT -26.280 24.950 -25.920 25.250 ;
        RECT -26.250 23.050 -25.950 24.950 ;
        RECT -26.850 22.750 -25.950 23.050 ;
        RECT -26.850 -42.450 -26.550 22.750 ;
        RECT -26.850 -42.750 4.350 -42.450 ;
        RECT 4.050 -64.850 4.350 -42.750 ;
        RECT 4.050 -65.150 15.450 -64.850 ;
        RECT 15.150 -68.350 15.450 -65.150 ;
        RECT 15.000 -72.350 15.600 -68.350 ;
    END
  END pd1_b
  PIN Ibias
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 206.000000 ;
    ANTENNADIFFAREA 30.160000 ;
    PORT
      LAYER li1 ;
        RECT -17.890 -22.200 -16.890 -22.030 ;
        RECT -16.600 -22.200 -15.600 -22.030 ;
        RECT -15.310 -22.200 -14.310 -22.030 ;
        RECT -14.020 -22.200 -13.020 -22.030 ;
        RECT -12.730 -22.200 -11.730 -22.030 ;
        RECT -11.440 -22.200 -10.440 -22.030 ;
        RECT -10.150 -22.200 -9.150 -22.030 ;
        RECT -8.860 -22.200 -7.860 -22.030 ;
        RECT -7.570 -22.200 -6.570 -22.030 ;
        RECT -6.280 -22.200 -5.280 -22.030 ;
        RECT -4.990 -22.200 -3.990 -22.030 ;
        RECT -3.700 -22.200 -2.700 -22.030 ;
        RECT -2.410 -22.200 -1.410 -22.030 ;
        RECT -1.120 -22.200 -0.120 -22.030 ;
        RECT 0.170 -22.200 1.170 -22.030 ;
        RECT 1.460 -22.200 2.460 -22.030 ;
        RECT 2.750 -22.200 3.750 -22.030 ;
        RECT 4.040 -22.200 5.040 -22.030 ;
        RECT 5.330 -22.200 6.330 -22.030 ;
        RECT 6.620 -22.200 7.620 -22.030 ;
        RECT 7.910 -22.200 8.910 -22.030 ;
        RECT 9.200 -22.200 10.200 -22.030 ;
        RECT 10.490 -22.200 11.490 -22.030 ;
        RECT 11.780 -22.200 12.780 -22.030 ;
        RECT 13.070 -22.200 14.070 -22.030 ;
        RECT -16.830 -24.100 -16.660 -22.370 ;
        RECT -14.250 -24.100 -14.080 -22.370 ;
        RECT -11.670 -24.100 -11.500 -22.370 ;
        RECT -9.090 -24.100 -8.920 -22.370 ;
        RECT -6.510 -24.100 -6.340 -22.370 ;
        RECT -3.930 -24.100 -3.760 -22.370 ;
        RECT -1.350 -24.100 -1.180 -22.370 ;
        RECT 1.230 -24.100 1.400 -22.370 ;
        RECT 3.810 -24.100 3.980 -22.370 ;
        RECT 6.390 -24.100 6.560 -22.370 ;
        RECT 8.970 -24.100 9.140 -22.370 ;
        RECT 11.550 -24.100 11.720 -22.370 ;
        RECT 14.130 -24.100 14.300 -22.370 ;
        RECT 16.080 -23.510 17.080 -23.340 ;
        RECT -17.000 -24.580 -16.600 -24.100 ;
        RECT -14.400 -24.580 -14.000 -24.100 ;
        RECT -11.800 -24.580 -11.400 -24.100 ;
        RECT -9.200 -24.580 -8.800 -24.100 ;
        RECT -6.600 -24.580 -6.200 -24.100 ;
        RECT -4.100 -24.580 -3.700 -24.100 ;
        RECT -1.500 -24.580 -1.100 -24.100 ;
        RECT 1.100 -24.580 1.500 -24.100 ;
        RECT 3.700 -24.580 4.100 -24.100 ;
        RECT 6.300 -24.580 6.700 -24.100 ;
        RECT 8.900 -24.580 9.300 -24.100 ;
        RECT 11.400 -24.580 11.800 -24.100 ;
        RECT 14.000 -24.580 14.400 -24.100 ;
        RECT -17.890 -24.600 -15.600 -24.580 ;
        RECT -15.310 -24.600 -13.020 -24.580 ;
        RECT -12.730 -24.600 -10.440 -24.580 ;
        RECT -10.150 -24.600 -7.860 -24.580 ;
        RECT -7.570 -24.600 -5.280 -24.580 ;
        RECT -4.990 -24.600 -2.700 -24.580 ;
        RECT -2.410 -24.600 -0.120 -24.580 ;
        RECT 0.170 -24.600 2.460 -24.580 ;
        RECT 2.750 -24.600 5.040 -24.580 ;
        RECT 5.330 -24.600 7.620 -24.580 ;
        RECT 7.910 -24.600 10.200 -24.580 ;
        RECT 10.490 -24.600 12.780 -24.580 ;
        RECT 13.070 -24.600 14.400 -24.580 ;
        RECT -17.900 -25.200 14.400 -24.600 ;
        RECT 16.000 -24.800 16.500 -24.700 ;
        RECT 19.300 -24.800 19.700 -24.700 ;
        RECT 16.000 -25.100 19.700 -24.800 ;
        RECT 16.000 -25.200 16.500 -25.100 ;
        RECT 19.300 -25.200 19.700 -25.100 ;
        RECT -17.890 -25.290 -15.600 -25.200 ;
        RECT -15.310 -25.290 -13.020 -25.200 ;
        RECT -12.730 -25.290 -10.440 -25.200 ;
        RECT -10.150 -25.290 -7.860 -25.200 ;
        RECT -7.570 -25.290 -5.280 -25.200 ;
        RECT -4.990 -25.290 -2.700 -25.200 ;
        RECT -2.410 -25.290 -0.120 -25.200 ;
        RECT 0.170 -25.290 2.460 -25.200 ;
        RECT 2.750 -25.290 5.040 -25.200 ;
        RECT 5.330 -25.290 7.620 -25.200 ;
        RECT 7.910 -25.290 10.200 -25.200 ;
        RECT 10.490 -25.290 12.780 -25.200 ;
        RECT 13.070 -25.290 14.400 -25.200 ;
        RECT -17.000 -25.800 -16.600 -25.290 ;
        RECT -14.400 -25.800 -14.000 -25.290 ;
        RECT -11.800 -25.800 -11.400 -25.290 ;
        RECT -9.200 -25.800 -8.800 -25.290 ;
        RECT -6.600 -25.800 -6.200 -25.290 ;
        RECT -4.100 -25.800 -3.700 -25.290 ;
        RECT -1.500 -25.800 -1.100 -25.290 ;
        RECT 1.100 -25.800 1.500 -25.290 ;
        RECT 3.700 -25.800 4.100 -25.290 ;
        RECT 6.300 -25.800 6.700 -25.290 ;
        RECT 8.900 -25.800 9.300 -25.290 ;
        RECT 11.400 -25.800 11.800 -25.290 ;
        RECT 14.000 -25.800 14.400 -25.290 ;
        RECT -16.830 -27.500 -16.660 -25.800 ;
        RECT -14.250 -27.500 -14.080 -25.800 ;
        RECT -11.670 -27.500 -11.500 -25.800 ;
        RECT -9.090 -27.500 -8.920 -25.800 ;
        RECT -6.510 -27.500 -6.340 -25.800 ;
        RECT -3.930 -27.500 -3.760 -25.800 ;
        RECT -1.350 -27.500 -1.180 -25.800 ;
        RECT 1.230 -27.500 1.400 -25.800 ;
        RECT 3.810 -27.500 3.980 -25.800 ;
        RECT 6.390 -27.500 6.560 -25.800 ;
        RECT 8.970 -27.500 9.140 -25.800 ;
        RECT 11.550 -27.500 11.720 -25.800 ;
        RECT 14.130 -27.500 14.300 -25.800 ;
        RECT 16.080 -26.670 17.080 -26.500 ;
        RECT 19.085 -26.665 20.085 -26.495 ;
        RECT -17.890 -27.840 -16.890 -27.670 ;
        RECT -16.600 -27.840 -15.600 -27.670 ;
        RECT -15.310 -27.840 -14.310 -27.670 ;
        RECT -14.020 -27.840 -13.020 -27.670 ;
        RECT -12.730 -27.840 -11.730 -27.670 ;
        RECT -11.440 -27.840 -10.440 -27.670 ;
        RECT -10.150 -27.840 -9.150 -27.670 ;
        RECT -8.860 -27.840 -7.860 -27.670 ;
        RECT -7.570 -27.840 -6.570 -27.670 ;
        RECT -6.280 -27.840 -5.280 -27.670 ;
        RECT -4.990 -27.840 -3.990 -27.670 ;
        RECT -3.700 -27.840 -2.700 -27.670 ;
        RECT -2.410 -27.840 -1.410 -27.670 ;
        RECT -1.120 -27.840 -0.120 -27.670 ;
        RECT 0.170 -27.840 1.170 -27.670 ;
        RECT 1.460 -27.840 2.460 -27.670 ;
        RECT 2.750 -27.840 3.750 -27.670 ;
        RECT 4.040 -27.840 5.040 -27.670 ;
        RECT 5.330 -27.840 6.330 -27.670 ;
        RECT 6.620 -27.840 7.620 -27.670 ;
        RECT 7.910 -27.840 8.910 -27.670 ;
        RECT 9.200 -27.840 10.200 -27.670 ;
        RECT 10.490 -27.840 11.490 -27.670 ;
        RECT 11.780 -27.840 12.780 -27.670 ;
        RECT 13.070 -27.840 14.070 -27.670 ;
        RECT -17.890 -29.600 -16.890 -29.430 ;
        RECT -16.600 -29.600 -15.600 -29.430 ;
        RECT -15.310 -29.600 -14.310 -29.430 ;
        RECT -14.020 -29.600 -13.020 -29.430 ;
        RECT -12.730 -29.600 -11.730 -29.430 ;
        RECT -11.440 -29.600 -10.440 -29.430 ;
        RECT -10.150 -29.600 -9.150 -29.430 ;
        RECT -8.860 -29.600 -7.860 -29.430 ;
        RECT -7.570 -29.600 -6.570 -29.430 ;
        RECT -6.280 -29.600 -5.280 -29.430 ;
        RECT -4.990 -29.600 -3.990 -29.430 ;
        RECT -3.700 -29.600 -2.700 -29.430 ;
        RECT -2.410 -29.600 -1.410 -29.430 ;
        RECT -1.120 -29.600 -0.120 -29.430 ;
        RECT 0.170 -29.600 1.170 -29.430 ;
        RECT 1.460 -29.600 2.460 -29.430 ;
        RECT 2.750 -29.600 3.750 -29.430 ;
        RECT 4.040 -29.600 5.040 -29.430 ;
        RECT 5.330 -29.600 6.330 -29.430 ;
        RECT 6.620 -29.600 7.620 -29.430 ;
        RECT 7.910 -29.600 8.910 -29.430 ;
        RECT 9.200 -29.600 10.200 -29.430 ;
        RECT 10.490 -29.600 11.490 -29.430 ;
        RECT 11.780 -29.600 12.780 -29.430 ;
        RECT 13.070 -29.600 14.070 -29.430 ;
        RECT -16.830 -31.500 -16.660 -29.770 ;
        RECT -14.250 -31.500 -14.080 -29.770 ;
        RECT -11.670 -31.500 -11.500 -29.770 ;
        RECT -9.090 -31.500 -8.920 -29.770 ;
        RECT -6.510 -31.500 -6.340 -29.770 ;
        RECT -3.930 -31.500 -3.760 -29.770 ;
        RECT -1.350 -31.500 -1.180 -29.770 ;
        RECT 1.230 -31.500 1.400 -29.770 ;
        RECT 3.810 -31.500 3.980 -29.770 ;
        RECT 6.390 -31.500 6.560 -29.770 ;
        RECT 8.970 -31.500 9.140 -29.770 ;
        RECT 11.550 -31.500 11.720 -29.770 ;
        RECT 14.130 -31.500 14.300 -29.770 ;
        RECT 16.080 -30.910 17.080 -30.740 ;
        RECT -17.000 -31.980 -16.600 -31.500 ;
        RECT -14.400 -31.980 -14.000 -31.500 ;
        RECT -11.800 -31.980 -11.400 -31.500 ;
        RECT -9.200 -31.980 -8.800 -31.500 ;
        RECT -6.600 -31.980 -6.200 -31.500 ;
        RECT -4.100 -31.980 -3.700 -31.500 ;
        RECT -1.500 -31.980 -1.100 -31.500 ;
        RECT 1.100 -31.980 1.500 -31.500 ;
        RECT 3.700 -31.980 4.100 -31.500 ;
        RECT 6.300 -31.980 6.700 -31.500 ;
        RECT 8.900 -31.980 9.300 -31.500 ;
        RECT 11.400 -31.980 11.800 -31.500 ;
        RECT 14.000 -31.980 14.400 -31.500 ;
        RECT -17.890 -32.000 -15.600 -31.980 ;
        RECT -15.310 -32.000 -13.020 -31.980 ;
        RECT -12.730 -32.000 -10.440 -31.980 ;
        RECT -10.150 -32.000 -7.860 -31.980 ;
        RECT -7.570 -32.000 -5.280 -31.980 ;
        RECT -4.990 -32.000 -2.700 -31.980 ;
        RECT -2.410 -32.000 -0.120 -31.980 ;
        RECT 0.170 -32.000 2.460 -31.980 ;
        RECT 2.750 -32.000 5.040 -31.980 ;
        RECT 5.330 -32.000 7.620 -31.980 ;
        RECT 7.910 -32.000 10.200 -31.980 ;
        RECT 10.490 -32.000 12.780 -31.980 ;
        RECT 13.070 -32.000 14.400 -31.980 ;
        RECT -17.900 -32.600 14.400 -32.000 ;
        RECT 16.000 -32.200 16.500 -32.100 ;
        RECT 19.300 -32.200 19.700 -32.100 ;
        RECT 16.000 -32.500 19.700 -32.200 ;
        RECT 16.000 -32.600 16.500 -32.500 ;
        RECT 19.300 -32.600 19.700 -32.500 ;
        RECT -17.890 -32.690 -15.600 -32.600 ;
        RECT -15.310 -32.690 -13.020 -32.600 ;
        RECT -12.730 -32.690 -10.440 -32.600 ;
        RECT -10.150 -32.690 -7.860 -32.600 ;
        RECT -7.570 -32.690 -5.280 -32.600 ;
        RECT -4.990 -32.690 -2.700 -32.600 ;
        RECT -2.410 -32.690 -0.120 -32.600 ;
        RECT 0.170 -32.690 2.460 -32.600 ;
        RECT 2.750 -32.690 5.040 -32.600 ;
        RECT 5.330 -32.690 7.620 -32.600 ;
        RECT 7.910 -32.690 10.200 -32.600 ;
        RECT 10.490 -32.690 12.780 -32.600 ;
        RECT 13.070 -32.690 14.400 -32.600 ;
        RECT -17.000 -33.200 -16.600 -32.690 ;
        RECT -14.400 -33.200 -14.000 -32.690 ;
        RECT -11.800 -33.200 -11.400 -32.690 ;
        RECT -9.200 -33.200 -8.800 -32.690 ;
        RECT -6.600 -33.200 -6.200 -32.690 ;
        RECT -4.100 -33.200 -3.700 -32.690 ;
        RECT -1.500 -33.200 -1.100 -32.690 ;
        RECT 1.100 -33.200 1.500 -32.690 ;
        RECT 3.700 -33.200 4.100 -32.690 ;
        RECT 6.300 -33.200 6.700 -32.690 ;
        RECT 8.900 -33.200 9.300 -32.690 ;
        RECT 11.400 -33.200 11.800 -32.690 ;
        RECT 14.000 -33.200 14.400 -32.690 ;
        RECT -16.830 -34.900 -16.660 -33.200 ;
        RECT -14.250 -34.900 -14.080 -33.200 ;
        RECT -11.670 -34.900 -11.500 -33.200 ;
        RECT -9.090 -34.900 -8.920 -33.200 ;
        RECT -6.510 -34.900 -6.340 -33.200 ;
        RECT -3.930 -34.900 -3.760 -33.200 ;
        RECT -1.350 -34.900 -1.180 -33.200 ;
        RECT 1.230 -34.900 1.400 -33.200 ;
        RECT 3.810 -34.900 3.980 -33.200 ;
        RECT 6.390 -34.900 6.560 -33.200 ;
        RECT 8.970 -34.900 9.140 -33.200 ;
        RECT 11.550 -34.900 11.720 -33.200 ;
        RECT 14.130 -34.900 14.300 -33.200 ;
        RECT 16.080 -34.070 17.080 -33.900 ;
        RECT 19.085 -34.065 20.085 -33.895 ;
        RECT -17.890 -35.240 -16.890 -35.070 ;
        RECT -16.600 -35.240 -15.600 -35.070 ;
        RECT -15.310 -35.240 -14.310 -35.070 ;
        RECT -14.020 -35.240 -13.020 -35.070 ;
        RECT -12.730 -35.240 -11.730 -35.070 ;
        RECT -11.440 -35.240 -10.440 -35.070 ;
        RECT -10.150 -35.240 -9.150 -35.070 ;
        RECT -8.860 -35.240 -7.860 -35.070 ;
        RECT -7.570 -35.240 -6.570 -35.070 ;
        RECT -6.280 -35.240 -5.280 -35.070 ;
        RECT -4.990 -35.240 -3.990 -35.070 ;
        RECT -3.700 -35.240 -2.700 -35.070 ;
        RECT -2.410 -35.240 -1.410 -35.070 ;
        RECT -1.120 -35.240 -0.120 -35.070 ;
        RECT 0.170 -35.240 1.170 -35.070 ;
        RECT 1.460 -35.240 2.460 -35.070 ;
        RECT 2.750 -35.240 3.750 -35.070 ;
        RECT 4.040 -35.240 5.040 -35.070 ;
        RECT 5.330 -35.240 6.330 -35.070 ;
        RECT 6.620 -35.240 7.620 -35.070 ;
        RECT 7.910 -35.240 8.910 -35.070 ;
        RECT 9.200 -35.240 10.200 -35.070 ;
        RECT 10.490 -35.240 11.490 -35.070 ;
        RECT 11.780 -35.240 12.780 -35.070 ;
        RECT 13.070 -35.240 14.070 -35.070 ;
      LAYER mcon ;
        RECT -16.830 -24.330 -16.660 -22.450 ;
        RECT -14.250 -24.330 -14.080 -22.450 ;
        RECT -11.670 -24.330 -11.500 -22.450 ;
        RECT -9.090 -24.330 -8.920 -22.450 ;
        RECT -6.510 -24.330 -6.340 -22.450 ;
        RECT -3.930 -24.330 -3.760 -22.450 ;
        RECT -1.350 -24.330 -1.180 -22.450 ;
        RECT 1.230 -24.330 1.400 -22.450 ;
        RECT 3.810 -24.330 3.980 -22.450 ;
        RECT 6.390 -24.330 6.560 -22.450 ;
        RECT 8.970 -24.330 9.140 -22.450 ;
        RECT 11.550 -24.330 11.720 -22.450 ;
        RECT 14.130 -24.330 14.300 -22.450 ;
        RECT 16.160 -23.510 17.000 -23.340 ;
        RECT -17.800 -25.100 14.000 -24.700 ;
        RECT 16.100 -25.100 16.400 -24.800 ;
        RECT 19.400 -25.100 19.600 -24.800 ;
        RECT -16.830 -27.420 -16.660 -25.540 ;
        RECT -14.250 -27.420 -14.080 -25.540 ;
        RECT -11.670 -27.420 -11.500 -25.540 ;
        RECT -9.090 -27.420 -8.920 -25.540 ;
        RECT -6.510 -27.420 -6.340 -25.540 ;
        RECT -3.930 -27.420 -3.760 -25.540 ;
        RECT -1.350 -27.420 -1.180 -25.540 ;
        RECT 1.230 -27.420 1.400 -25.540 ;
        RECT 3.810 -27.420 3.980 -25.540 ;
        RECT 6.390 -27.420 6.560 -25.540 ;
        RECT 8.970 -27.420 9.140 -25.540 ;
        RECT 11.550 -27.420 11.720 -25.540 ;
        RECT 14.130 -27.420 14.300 -25.540 ;
        RECT 16.160 -26.670 17.000 -26.500 ;
        RECT 19.205 -26.665 19.965 -26.495 ;
        RECT -16.830 -31.730 -16.660 -29.850 ;
        RECT -14.250 -31.730 -14.080 -29.850 ;
        RECT -11.670 -31.730 -11.500 -29.850 ;
        RECT -9.090 -31.730 -8.920 -29.850 ;
        RECT -6.510 -31.730 -6.340 -29.850 ;
        RECT -3.930 -31.730 -3.760 -29.850 ;
        RECT -1.350 -31.730 -1.180 -29.850 ;
        RECT 1.230 -31.730 1.400 -29.850 ;
        RECT 3.810 -31.730 3.980 -29.850 ;
        RECT 6.390 -31.730 6.560 -29.850 ;
        RECT 8.970 -31.730 9.140 -29.850 ;
        RECT 11.550 -31.730 11.720 -29.850 ;
        RECT 14.130 -31.730 14.300 -29.850 ;
        RECT 16.160 -30.910 17.000 -30.740 ;
        RECT -17.800 -32.500 14.000 -32.100 ;
        RECT 16.100 -32.500 16.400 -32.200 ;
        RECT 19.400 -32.500 19.600 -32.200 ;
        RECT -16.830 -34.820 -16.660 -32.940 ;
        RECT -14.250 -34.820 -14.080 -32.940 ;
        RECT -11.670 -34.820 -11.500 -32.940 ;
        RECT -9.090 -34.820 -8.920 -32.940 ;
        RECT -6.510 -34.820 -6.340 -32.940 ;
        RECT -3.930 -34.820 -3.760 -32.940 ;
        RECT -1.350 -34.820 -1.180 -32.940 ;
        RECT 1.230 -34.820 1.400 -32.940 ;
        RECT 3.810 -34.820 3.980 -32.940 ;
        RECT 6.390 -34.820 6.560 -32.940 ;
        RECT 8.970 -34.820 9.140 -32.940 ;
        RECT 11.550 -34.820 11.720 -32.940 ;
        RECT 14.130 -34.820 14.300 -32.940 ;
        RECT 16.160 -34.070 17.000 -33.900 ;
        RECT 19.205 -34.065 19.965 -33.895 ;
      LAYER met1 ;
        RECT -54.250 -21.000 -49.750 -20.970 ;
        RECT -54.250 -25.500 -30.250 -21.000 ;
        RECT -54.250 -25.530 -49.750 -25.500 ;
        RECT -34.750 -26.750 -30.250 -25.500 ;
        RECT -20.000 -24.600 -18.300 -24.200 ;
        RECT -16.860 -24.390 -16.630 -22.390 ;
        RECT -14.280 -24.390 -14.050 -22.390 ;
        RECT -11.700 -24.390 -11.470 -22.390 ;
        RECT -9.120 -24.390 -8.890 -22.390 ;
        RECT -6.540 -24.390 -6.310 -22.390 ;
        RECT -3.960 -24.390 -3.730 -22.390 ;
        RECT -1.380 -24.390 -1.150 -22.390 ;
        RECT 1.200 -24.390 1.430 -22.390 ;
        RECT 3.780 -24.390 4.010 -22.390 ;
        RECT 6.360 -24.390 6.590 -22.390 ;
        RECT 8.940 -24.390 9.170 -22.390 ;
        RECT 11.520 -24.390 11.750 -22.390 ;
        RECT 14.100 -24.390 14.330 -22.390 ;
        RECT 16.100 -23.310 16.400 -23.300 ;
        RECT 16.100 -23.540 17.060 -23.310 ;
        RECT -20.000 -24.800 14.100 -24.600 ;
        RECT 16.100 -24.700 16.400 -23.540 ;
        RECT 16.000 -24.800 16.500 -24.700 ;
        RECT -20.000 -25.100 16.500 -24.800 ;
        RECT -20.000 -25.200 14.100 -25.100 ;
        RECT 16.000 -25.200 16.500 -25.100 ;
        RECT 19.300 -25.200 19.700 -24.700 ;
        RECT -20.000 -25.500 -18.300 -25.200 ;
        RECT -20.000 -26.750 -18.800 -25.500 ;
        RECT -34.750 -31.500 -18.800 -26.750 ;
        RECT -16.860 -27.480 -16.630 -25.480 ;
        RECT -14.280 -27.480 -14.050 -25.480 ;
        RECT -11.700 -27.480 -11.470 -25.480 ;
        RECT -9.120 -27.480 -8.890 -25.480 ;
        RECT -6.540 -27.480 -6.310 -25.480 ;
        RECT -3.960 -27.480 -3.730 -25.480 ;
        RECT -1.380 -27.480 -1.150 -25.480 ;
        RECT 1.200 -27.480 1.430 -25.480 ;
        RECT 3.780 -27.480 4.010 -25.480 ;
        RECT 6.360 -27.480 6.590 -25.480 ;
        RECT 8.940 -27.480 9.170 -25.480 ;
        RECT 11.520 -27.480 11.750 -25.480 ;
        RECT 14.100 -27.480 14.330 -25.480 ;
        RECT 16.100 -26.470 16.400 -25.200 ;
        RECT 19.400 -26.465 19.600 -25.200 ;
        RECT 16.100 -26.700 17.060 -26.470 ;
        RECT 19.145 -26.695 20.025 -26.465 ;
        RECT 19.400 -26.700 19.600 -26.695 ;
        RECT -34.750 -31.750 -30.250 -31.500 ;
        RECT -20.000 -31.600 -18.800 -31.500 ;
        RECT -20.000 -32.000 -18.300 -31.600 ;
        RECT -16.860 -31.790 -16.630 -29.790 ;
        RECT -14.280 -31.790 -14.050 -29.790 ;
        RECT -11.700 -31.790 -11.470 -29.790 ;
        RECT -9.120 -31.790 -8.890 -29.790 ;
        RECT -6.540 -31.790 -6.310 -29.790 ;
        RECT -3.960 -31.790 -3.730 -29.790 ;
        RECT -1.380 -31.790 -1.150 -29.790 ;
        RECT 1.200 -31.790 1.430 -29.790 ;
        RECT 3.780 -31.790 4.010 -29.790 ;
        RECT 6.360 -31.790 6.590 -29.790 ;
        RECT 8.940 -31.790 9.170 -29.790 ;
        RECT 11.520 -31.790 11.750 -29.790 ;
        RECT 14.100 -31.790 14.330 -29.790 ;
        RECT 16.100 -30.710 16.400 -30.700 ;
        RECT 16.100 -30.940 17.060 -30.710 ;
        RECT -20.000 -32.200 14.100 -32.000 ;
        RECT 16.100 -32.100 16.400 -30.940 ;
        RECT 16.000 -32.200 16.500 -32.100 ;
        RECT -20.000 -32.500 16.500 -32.200 ;
        RECT -20.000 -32.600 14.100 -32.500 ;
        RECT 16.000 -32.600 16.500 -32.500 ;
        RECT 19.300 -32.600 19.700 -32.100 ;
        RECT -20.000 -32.900 -18.300 -32.600 ;
        RECT -20.000 -33.000 -18.800 -32.900 ;
        RECT -16.860 -34.880 -16.630 -32.880 ;
        RECT -14.280 -34.880 -14.050 -32.880 ;
        RECT -11.700 -34.880 -11.470 -32.880 ;
        RECT -9.120 -34.880 -8.890 -32.880 ;
        RECT -6.540 -34.880 -6.310 -32.880 ;
        RECT -3.960 -34.880 -3.730 -32.880 ;
        RECT -1.380 -34.880 -1.150 -32.880 ;
        RECT 1.200 -34.880 1.430 -32.880 ;
        RECT 3.780 -34.880 4.010 -32.880 ;
        RECT 6.360 -34.880 6.590 -32.880 ;
        RECT 8.940 -34.880 9.170 -32.880 ;
        RECT 11.520 -34.880 11.750 -32.880 ;
        RECT 14.100 -34.880 14.330 -32.880 ;
        RECT 16.100 -33.870 16.400 -32.600 ;
        RECT 19.400 -33.865 19.600 -32.600 ;
        RECT 16.100 -34.100 17.060 -33.870 ;
        RECT 19.145 -34.095 20.025 -33.865 ;
        RECT 19.400 -34.100 19.600 -34.095 ;
      LAYER met2 ;
        RECT -57.500 -25.500 -49.720 -21.000 ;
    END
  END Ibias
  PIN Vd1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT -0.850 14.150 -0.350 14.250 ;
        RECT -0.850 13.950 0.500 14.150 ;
        RECT -0.435 13.930 -0.105 13.950 ;
        RECT 0.155 13.930 0.485 13.950 ;
      LAYER mcon ;
        RECT -0.800 14.000 -0.400 14.200 ;
      LAYER met1 ;
        RECT -0.900 13.900 -0.300 14.300 ;
      LAYER via ;
        RECT -0.850 13.950 -0.350 14.250 ;
      LAYER met2 ;
        RECT -0.900 14.250 -0.300 14.300 ;
        RECT -2.150 14.200 -0.300 14.250 ;
        RECT -23.300 13.950 -0.300 14.200 ;
        RECT -23.300 13.900 -1.850 13.950 ;
        RECT -0.900 13.900 -0.300 13.950 ;
        RECT -23.300 -38.800 -23.000 13.900 ;
        RECT -23.300 -39.100 8.200 -38.800 ;
        RECT 7.900 -61.350 8.200 -39.100 ;
        RECT 7.900 -61.650 55.450 -61.350 ;
        RECT 55.150 -68.350 55.450 -61.650 ;
        RECT 55.000 -72.350 55.600 -68.350 ;
    END
  END Vd1
  PIN Vd2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 2.365 12.850 2.695 12.860 ;
        RECT 2.955 12.850 3.285 12.860 ;
        RECT 2.365 12.690 3.600 12.850 ;
        RECT 2.400 12.550 3.600 12.690 ;
      LAYER mcon ;
        RECT 3.000 12.600 3.550 12.800 ;
      LAYER met1 ;
        RECT 2.900 12.350 3.650 12.900 ;
      LAYER via ;
        RECT 3.000 12.400 3.500 12.800 ;
      LAYER met2 ;
        RECT -22.800 12.750 -1.750 12.800 ;
        RECT 2.900 12.750 3.650 12.900 ;
        RECT -22.800 12.500 3.650 12.750 ;
        RECT -22.800 -38.300 -22.500 12.500 ;
        RECT -2.150 12.450 3.650 12.500 ;
        RECT 2.900 12.350 3.650 12.450 ;
        RECT -22.800 -38.600 8.700 -38.300 ;
        RECT 8.400 -60.850 8.700 -38.600 ;
        RECT 8.400 -61.150 60.450 -60.850 ;
        RECT 60.150 -68.350 60.450 -61.150 ;
        RECT 60.000 -72.350 60.600 -68.350 ;
    END
  END Vd2
  PIN sw1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.200000 ;
    PORT
      LAYER li1 ;
        RECT -19.020 7.000 -18.670 7.065 ;
        RECT -8.620 7.000 -8.270 7.065 ;
        RECT -19.100 6.895 -18.670 7.000 ;
        RECT -8.700 6.895 -8.270 7.000 ;
        RECT -19.100 6.800 -18.700 6.895 ;
        RECT -8.700 6.800 -8.300 6.895 ;
        RECT -20.100 6.500 -19.700 6.600 ;
        RECT -19.100 6.500 -18.800 6.800 ;
        RECT -20.100 6.200 -18.800 6.500 ;
        RECT -20.100 6.100 -19.700 6.200 ;
        RECT -19.100 6.000 -18.800 6.200 ;
        RECT -9.700 6.500 -9.200 6.600 ;
        RECT -8.700 6.500 -8.400 6.800 ;
        RECT -9.700 6.200 -8.400 6.500 ;
        RECT -9.700 6.100 -9.200 6.200 ;
        RECT -8.700 6.000 -8.400 6.200 ;
        RECT -19.100 5.800 -16.400 6.000 ;
        RECT -19.100 5.500 -18.800 5.800 ;
        RECT -16.600 5.600 -16.400 5.800 ;
        RECT -8.700 5.800 -6.000 6.000 ;
        RECT -16.600 5.500 -15.700 5.600 ;
        RECT -8.700 5.500 -8.400 5.800 ;
        RECT -6.200 5.600 -6.000 5.800 ;
        RECT -6.200 5.500 -5.300 5.600 ;
        RECT -19.110 5.330 -18.780 5.500 ;
        RECT -16.635 5.400 -15.700 5.500 ;
        RECT -16.635 5.330 -16.305 5.400 ;
        RECT -16.045 5.330 -15.715 5.400 ;
        RECT -8.710 5.330 -8.380 5.500 ;
        RECT -6.235 5.400 -5.300 5.500 ;
        RECT -6.235 5.330 -5.905 5.400 ;
        RECT -5.645 5.330 -5.315 5.400 ;
      LAYER mcon ;
        RECT -20.000 6.200 -19.800 6.500 ;
        RECT -9.600 6.200 -9.300 6.500 ;
      LAYER met1 ;
        RECT -20.100 6.100 -19.600 6.600 ;
        RECT -9.700 6.100 -9.200 6.600 ;
      LAYER via ;
        RECT -20.000 6.200 -19.700 6.500 ;
        RECT -9.600 6.200 -9.300 6.500 ;
      LAYER met2 ;
        RECT -20.100 6.500 -19.600 6.600 ;
        RECT -21.800 6.200 -19.600 6.500 ;
        RECT -21.800 -37.300 -21.500 6.200 ;
        RECT -20.100 6.100 -19.600 6.200 ;
        RECT -9.700 6.100 -9.200 6.600 ;
        RECT -20.000 2.700 -19.700 6.100 ;
        RECT -9.600 2.700 -9.300 6.100 ;
        RECT -20.000 2.400 -9.300 2.700 ;
        RECT -21.800 -37.600 9.700 -37.300 ;
        RECT 9.400 -59.850 9.700 -37.600 ;
        RECT 9.400 -60.150 70.400 -59.850 ;
        RECT 70.100 -68.350 70.400 -60.150 ;
        RECT 70.000 -72.350 70.600 -68.350 ;
    END
  END sw1
  PIN sw2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.200000 ;
    PORT
      LAYER li1 ;
        RECT -13.820 7.000 -13.470 7.065 ;
        RECT -3.420 7.000 -3.070 7.065 ;
        RECT -13.900 6.895 -13.470 7.000 ;
        RECT -3.500 6.895 -3.070 7.000 ;
        RECT -13.900 6.800 -13.500 6.895 ;
        RECT -3.500 6.800 -3.100 6.895 ;
        RECT -15.000 6.500 -14.500 6.600 ;
        RECT -13.900 6.500 -13.600 6.800 ;
        RECT -15.000 6.200 -13.600 6.500 ;
        RECT -15.000 6.100 -14.500 6.200 ;
        RECT -13.900 6.000 -13.600 6.200 ;
        RECT -4.600 6.500 -4.100 6.600 ;
        RECT -3.500 6.500 -3.200 6.800 ;
        RECT -4.600 6.200 -3.200 6.500 ;
        RECT -4.600 6.100 -4.100 6.200 ;
        RECT -3.500 6.000 -3.200 6.200 ;
        RECT -13.900 5.800 -11.200 6.000 ;
        RECT -13.900 5.500 -13.600 5.800 ;
        RECT -11.400 5.600 -11.200 5.800 ;
        RECT -3.500 5.800 -0.800 6.000 ;
        RECT -11.400 5.500 -10.500 5.600 ;
        RECT -3.500 5.500 -3.200 5.800 ;
        RECT -1.000 5.600 -0.800 5.800 ;
        RECT -1.000 5.500 -0.100 5.600 ;
        RECT -13.910 5.330 -13.580 5.500 ;
        RECT -11.435 5.400 -10.500 5.500 ;
        RECT -11.435 5.330 -11.105 5.400 ;
        RECT -10.845 5.330 -10.515 5.400 ;
        RECT -3.510 5.330 -3.180 5.500 ;
        RECT -1.035 5.400 -0.100 5.500 ;
        RECT -1.035 5.330 -0.705 5.400 ;
        RECT -0.445 5.330 -0.115 5.400 ;
      LAYER mcon ;
        RECT -14.900 6.200 -14.600 6.500 ;
        RECT -4.500 6.200 -4.200 6.500 ;
      LAYER met1 ;
        RECT -15.000 6.100 -14.500 6.600 ;
        RECT -4.600 6.100 -4.100 6.600 ;
      LAYER via ;
        RECT -14.900 6.200 -14.600 6.500 ;
        RECT -4.500 6.200 -4.200 6.500 ;
      LAYER met2 ;
        RECT -22.300 10.300 -14.600 10.600 ;
        RECT -22.300 -37.800 -22.000 10.300 ;
        RECT -14.900 9.900 -14.600 10.300 ;
        RECT -14.900 9.600 -4.200 9.900 ;
        RECT -14.900 6.600 -14.600 9.600 ;
        RECT -4.500 6.600 -4.200 9.600 ;
        RECT -15.000 6.100 -14.500 6.600 ;
        RECT -4.600 6.100 -4.100 6.600 ;
        RECT -22.300 -38.100 9.200 -37.800 ;
        RECT 8.900 -60.350 9.200 -38.100 ;
        RECT 8.900 -60.650 65.450 -60.350 ;
        RECT 65.150 -68.350 65.450 -60.650 ;
        RECT 65.000 -72.350 65.600 -68.350 ;
    END
  END sw2
  PIN sh
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 0.965 -8.750 1.295 -8.740 ;
        RECT 1.555 -8.750 1.885 -8.740 ;
        RECT 0.550 -8.950 1.900 -8.750 ;
        RECT 0.550 -9.050 0.950 -8.950 ;
      LAYER mcon ;
        RECT 0.600 -9.000 0.900 -8.800 ;
      LAYER met1 ;
        RECT 0.500 -9.050 1.000 -8.750 ;
        RECT 0.650 -17.800 0.850 -9.050 ;
        RECT 26.670 -17.800 26.930 -17.740 ;
        RECT 0.650 -18.000 26.930 -17.800 ;
        RECT 26.670 -18.060 26.930 -18.000 ;
        RECT 26.640 -37.430 26.960 -37.170 ;
        RECT 26.700 -65.900 26.900 -37.430 ;
        RECT 72.240 -65.900 72.560 -65.870 ;
        RECT 26.700 -66.100 72.560 -65.900 ;
        RECT 72.240 -66.130 72.560 -66.100 ;
      LAYER via ;
        RECT 26.670 -18.030 26.930 -17.770 ;
        RECT 26.670 -37.430 26.930 -37.170 ;
        RECT 72.270 -66.130 72.530 -65.870 ;
      LAYER met2 ;
        RECT 26.640 -18.030 26.960 -17.770 ;
        RECT 26.700 -37.140 26.900 -18.030 ;
        RECT 26.670 -37.460 26.930 -37.140 ;
        RECT 72.270 -65.900 72.530 -65.840 ;
        RECT 72.270 -66.100 85.300 -65.900 ;
        RECT 72.270 -66.160 72.530 -66.100 ;
        RECT 85.100 -68.500 85.300 -66.100 ;
        RECT 85.000 -72.400 85.600 -68.500 ;
    END
  END sh
  PIN sh_cmp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 47.015 -37.850 47.345 -37.840 ;
        RECT 47.605 -37.850 47.935 -37.840 ;
        RECT 47.000 -38.150 48.350 -37.850 ;
      LAYER mcon ;
        RECT 48.050 -38.100 48.250 -37.900 ;
      LAYER met1 ;
        RECT 47.950 -38.150 48.350 -37.850 ;
        RECT 48.000 -52.750 48.300 -38.150 ;
        RECT 48.000 -53.050 80.450 -52.750 ;
        RECT 80.150 -69.430 80.450 -53.050 ;
      LAYER via ;
        RECT 80.150 -69.400 80.450 -69.100 ;
      LAYER met2 ;
        RECT 80.000 -72.350 80.600 -68.350 ;
    END
  END sh_cmp
  PIN sh_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 44.165 -37.900 44.495 -37.840 ;
        RECT 44.755 -37.850 45.085 -37.840 ;
        RECT 44.755 -37.900 45.500 -37.850 ;
        RECT 44.165 -38.010 45.500 -37.900 ;
        RECT 44.200 -38.100 45.500 -38.010 ;
        RECT 45.000 -38.150 45.500 -38.100 ;
      LAYER mcon ;
        RECT 45.100 -38.100 45.400 -37.900 ;
      LAYER met1 ;
        RECT 45.000 -38.150 45.500 -37.850 ;
        RECT 45.100 -53.550 45.400 -38.150 ;
        RECT 45.100 -53.850 75.450 -53.550 ;
        RECT 75.150 -69.430 75.450 -53.850 ;
      LAYER via ;
        RECT 75.150 -69.400 75.450 -69.100 ;
      LAYER met2 ;
        RECT 75.000 -72.350 75.600 -68.350 ;
    END
  END sh_rst
  PIN OTA_out_c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.100000 ;
    PORT
      LAYER li1 ;
        RECT 19.680 11.450 20.030 11.515 ;
        RECT 19.600 11.345 20.030 11.450 ;
        RECT 19.600 11.250 20.000 11.345 ;
        RECT 19.600 10.950 19.900 11.250 ;
        RECT 18.600 10.650 19.900 10.950 ;
        RECT 19.600 10.450 19.900 10.650 ;
        RECT 19.600 10.250 22.300 10.450 ;
        RECT 19.600 9.950 19.900 10.250 ;
        RECT 22.100 10.050 22.300 10.250 ;
        RECT 22.100 9.950 23.000 10.050 ;
        RECT 19.590 9.780 19.920 9.950 ;
        RECT 22.065 9.850 23.000 9.950 ;
        RECT 22.065 9.780 22.395 9.850 ;
        RECT 22.655 9.780 22.985 9.850 ;
      LAYER met1 ;
        RECT 11.700 16.550 12.100 16.950 ;
        RECT 11.750 16.400 12.050 16.550 ;
        RECT 11.750 16.100 18.950 16.400 ;
        RECT 18.540 10.620 18.960 10.980 ;
      LAYER via ;
        RECT 11.750 16.600 12.050 16.900 ;
        RECT 18.600 16.100 18.900 16.400 ;
        RECT 18.570 10.620 18.930 10.980 ;
      LAYER met2 ;
        RECT -25.800 -41.300 -25.500 18.745 ;
        RECT 11.700 16.550 12.100 16.950 ;
        RECT 18.600 11.050 18.900 16.430 ;
        RECT 18.500 10.550 19.000 11.050 ;
        RECT -25.800 -41.600 5.450 -41.300 ;
        RECT 5.150 -63.850 5.450 -41.600 ;
        RECT 5.150 -64.150 30.450 -63.850 ;
        RECT 30.150 -68.350 30.450 -64.150 ;
        RECT 30.000 -72.350 30.600 -68.350 ;
      LAYER via2 ;
        RECT -25.800 18.400 -25.500 18.700 ;
        RECT 11.760 16.610 12.040 16.890 ;
      LAYER met3 ;
        RECT -25.825 18.700 -25.475 18.725 ;
        RECT -25.825 18.400 12.050 18.700 ;
        RECT -25.825 18.375 -25.475 18.400 ;
        RECT 11.750 16.915 12.050 18.400 ;
        RECT 11.735 16.585 12.065 16.915 ;
    END
  END OTA_out_c
  PIN SH_out_c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.100000 ;
    PORT
      LAYER li1 ;
        RECT 24.930 11.450 25.280 11.515 ;
        RECT 24.850 11.345 25.280 11.450 ;
        RECT 24.850 11.250 25.250 11.345 ;
        RECT 24.850 10.950 25.150 11.250 ;
        RECT 23.850 10.650 25.150 10.950 ;
        RECT 24.850 10.450 25.150 10.650 ;
        RECT 24.850 10.250 27.550 10.450 ;
        RECT 24.850 9.950 25.150 10.250 ;
        RECT 27.350 10.050 27.550 10.250 ;
        RECT 27.350 9.950 28.250 10.050 ;
        RECT 24.840 9.780 25.170 9.950 ;
        RECT 27.315 9.850 28.250 9.950 ;
        RECT 27.315 9.780 27.645 9.850 ;
        RECT 27.905 9.780 28.235 9.850 ;
      LAYER met1 ;
        RECT 11.000 15.900 11.400 16.300 ;
        RECT 11.050 15.600 24.180 15.900 ;
        RECT 23.790 10.620 24.210 10.980 ;
      LAYER via ;
        RECT 11.050 15.950 11.350 16.250 ;
        RECT 23.850 15.600 24.150 15.900 ;
        RECT 23.820 10.620 24.180 10.980 ;
      LAYER met2 ;
        RECT -25.300 -40.800 -25.000 18.045 ;
        RECT 11.000 15.900 11.400 16.300 ;
        RECT 23.850 11.050 24.150 15.930 ;
        RECT 23.750 10.550 24.250 11.050 ;
        RECT -25.300 -41.100 6.050 -40.800 ;
        RECT 5.750 -63.350 6.050 -41.100 ;
        RECT 5.750 -63.650 35.450 -63.350 ;
        RECT 35.150 -68.350 35.450 -63.650 ;
        RECT 35.000 -72.350 35.600 -68.350 ;
      LAYER via2 ;
        RECT -25.300 17.700 -25.000 18.000 ;
        RECT 11.060 15.960 11.340 16.240 ;
      LAYER met3 ;
        RECT -25.325 18.000 -24.975 18.025 ;
        RECT -25.325 17.700 11.350 18.000 ;
        RECT -25.325 17.675 -24.975 17.700 ;
        RECT 11.050 16.265 11.350 17.700 ;
        RECT 11.035 15.935 11.365 16.265 ;
    END
  END SH_out_c
  PIN Vref_cmp_c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.100000 ;
    PORT
      LAYER li1 ;
        RECT 30.180 11.450 30.530 11.515 ;
        RECT 30.100 11.345 30.530 11.450 ;
        RECT 30.100 11.250 30.500 11.345 ;
        RECT 30.100 10.950 30.400 11.250 ;
        RECT 29.100 10.650 30.400 10.950 ;
        RECT 30.100 10.450 30.400 10.650 ;
        RECT 30.100 10.250 32.800 10.450 ;
        RECT 30.100 9.950 30.400 10.250 ;
        RECT 32.600 10.050 32.800 10.250 ;
        RECT 32.600 9.950 33.500 10.050 ;
        RECT 30.090 9.780 30.420 9.950 ;
        RECT 32.565 9.850 33.500 9.950 ;
        RECT 32.565 9.780 32.895 9.850 ;
        RECT 33.155 9.780 33.485 9.850 ;
      LAYER mcon ;
        RECT 29.150 10.650 29.450 10.950 ;
      LAYER met1 ;
        RECT 10.300 15.400 10.700 15.700 ;
        RECT 29.100 15.400 29.500 15.450 ;
        RECT 10.300 15.300 29.500 15.400 ;
        RECT 10.350 15.100 29.500 15.300 ;
        RECT 29.100 15.050 29.500 15.100 ;
        RECT 29.090 10.620 29.510 10.980 ;
      LAYER via ;
        RECT 10.350 15.350 10.650 15.650 ;
        RECT 29.150 15.100 29.450 15.400 ;
        RECT 29.120 10.620 29.480 10.980 ;
      LAYER met2 ;
        RECT -24.800 -40.300 -24.500 17.345 ;
        RECT 10.300 15.300 10.700 15.700 ;
        RECT 29.100 15.050 29.500 15.450 ;
        RECT 29.150 11.050 29.450 15.050 ;
        RECT 29.050 10.550 29.550 11.050 ;
        RECT -24.800 -40.600 6.650 -40.300 ;
        RECT 6.350 -62.850 6.650 -40.600 ;
        RECT 6.350 -63.150 40.450 -62.850 ;
        RECT 40.150 -68.350 40.450 -63.150 ;
        RECT 40.000 -72.350 40.600 -68.350 ;
      LAYER via2 ;
        RECT -24.800 17.000 -24.500 17.300 ;
        RECT 10.360 15.360 10.640 15.640 ;
      LAYER met3 ;
        RECT -24.825 17.300 -24.475 17.325 ;
        RECT -24.825 17.000 10.650 17.300 ;
        RECT -24.825 16.975 -24.475 17.000 ;
        RECT 10.350 15.665 10.650 17.000 ;
        RECT 10.335 15.335 10.665 15.665 ;
    END
  END Vref_cmp_c
  PIN OTA_sh_c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.100000 ;
    PORT
      LAYER li1 ;
        RECT 35.380 11.450 35.730 11.515 ;
        RECT 35.300 11.345 35.730 11.450 ;
        RECT 35.300 11.250 35.700 11.345 ;
        RECT 35.300 10.950 35.600 11.250 ;
        RECT 34.300 10.650 35.600 10.950 ;
        RECT 35.300 10.450 35.600 10.650 ;
        RECT 35.300 10.250 38.000 10.450 ;
        RECT 35.300 9.950 35.600 10.250 ;
        RECT 37.800 10.050 38.000 10.250 ;
        RECT 37.800 9.950 38.700 10.050 ;
        RECT 35.290 9.780 35.620 9.950 ;
        RECT 37.765 9.850 38.700 9.950 ;
        RECT 37.765 9.780 38.095 9.850 ;
        RECT 38.355 9.780 38.685 9.850 ;
      LAYER met1 ;
        RECT 9.550 14.900 9.950 15.250 ;
        RECT 34.300 14.900 34.600 14.930 ;
        RECT 9.550 14.850 34.600 14.900 ;
        RECT 9.600 14.600 34.600 14.850 ;
        RECT 34.300 14.570 34.600 14.600 ;
        RECT 34.240 10.620 34.660 10.980 ;
      LAYER via ;
        RECT 9.600 14.900 9.900 15.200 ;
        RECT 34.300 14.600 34.600 14.900 ;
        RECT 34.270 10.620 34.630 10.980 ;
      LAYER met2 ;
        RECT -24.300 -39.800 -24.000 16.695 ;
        RECT 9.550 14.850 9.950 15.250 ;
        RECT 34.270 14.600 34.630 14.900 ;
        RECT 34.300 11.050 34.600 14.600 ;
        RECT 34.200 10.550 34.700 11.050 ;
        RECT -24.300 -40.100 7.150 -39.800 ;
        RECT 6.850 -62.350 7.150 -40.100 ;
        RECT 6.850 -62.650 45.450 -62.350 ;
        RECT 45.150 -68.350 45.450 -62.650 ;
        RECT 45.000 -72.350 45.600 -68.350 ;
      LAYER via2 ;
        RECT -24.300 16.350 -24.000 16.650 ;
        RECT 9.610 14.910 9.890 15.190 ;
      LAYER met3 ;
        RECT -24.325 16.650 -23.975 16.675 ;
        RECT -24.325 16.350 9.900 16.650 ;
        RECT -24.325 16.325 -23.975 16.350 ;
        RECT 9.600 15.250 9.900 16.350 ;
        RECT 9.550 14.850 9.950 15.250 ;
    END
  END OTA_sh_c
  PIN CMP_out_c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.100000 ;
    PORT
      LAYER li1 ;
        RECT 40.630 11.450 40.980 11.515 ;
        RECT 40.550 11.345 40.980 11.450 ;
        RECT 40.550 11.250 40.950 11.345 ;
        RECT 40.550 10.950 40.850 11.250 ;
        RECT 39.550 10.650 40.850 10.950 ;
        RECT 40.550 10.450 40.850 10.650 ;
        RECT 40.550 10.250 43.250 10.450 ;
        RECT 40.550 9.950 40.850 10.250 ;
        RECT 43.050 10.050 43.250 10.250 ;
        RECT 43.050 9.950 43.950 10.050 ;
        RECT 40.540 9.780 40.870 9.950 ;
        RECT 43.015 9.850 43.950 9.950 ;
        RECT 43.015 9.780 43.345 9.850 ;
        RECT 43.605 9.780 43.935 9.850 ;
      LAYER met1 ;
        RECT 39.550 14.450 39.850 14.480 ;
        RECT 8.720 14.400 34.150 14.450 ;
        RECT 34.750 14.400 39.850 14.450 ;
        RECT 8.720 14.150 39.850 14.400 ;
        RECT 39.550 14.120 39.850 14.150 ;
        RECT 39.520 10.980 39.880 11.010 ;
        RECT 39.490 10.620 39.910 10.980 ;
      LAYER via ;
        RECT 8.750 14.150 9.050 14.450 ;
        RECT 39.550 14.150 39.850 14.450 ;
        RECT 39.520 10.680 39.880 10.980 ;
      LAYER met2 ;
        RECT -23.800 -39.300 -23.500 15.995 ;
        RECT 8.750 14.105 9.050 14.495 ;
        RECT 39.520 14.150 39.880 14.450 ;
        RECT 39.550 10.980 39.850 14.150 ;
        RECT 39.490 10.680 39.910 10.980 ;
        RECT -23.800 -39.600 7.700 -39.300 ;
        RECT 7.400 -61.850 7.700 -39.600 ;
        RECT 7.400 -62.150 50.450 -61.850 ;
        RECT 50.150 -68.350 50.450 -62.150 ;
        RECT 50.000 -72.350 50.600 -68.350 ;
      LAYER via2 ;
        RECT -23.800 15.650 -23.500 15.950 ;
        RECT 8.750 14.150 9.050 14.450 ;
      LAYER met3 ;
        RECT -23.825 15.950 -23.475 15.975 ;
        RECT -23.850 15.650 9.050 15.950 ;
        RECT -23.825 15.625 -23.475 15.650 ;
        RECT 8.750 14.475 9.050 15.650 ;
        RECT 8.725 14.125 9.075 14.475 ;
    END
  END CMP_out_c
  PIN PD2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT -17.220 25.630 -16.180 25.800 ;
        RECT -15.350 25.550 -15.050 26.000 ;
        RECT -15.250 24.750 -15.050 25.550 ;
        RECT -17.220 24.450 -16.180 24.620 ;
        RECT -15.300 24.300 -15.000 24.750 ;
        RECT -17.270 22.430 -16.230 22.600 ;
        RECT -17.270 21.250 -16.230 21.420 ;
      LAYER mcon ;
        RECT -17.140 25.630 -16.260 25.800 ;
        RECT -15.300 25.650 -15.100 25.900 ;
        RECT -17.140 24.450 -16.260 24.620 ;
        RECT -15.250 24.400 -15.050 24.650 ;
        RECT -17.190 22.430 -16.310 22.600 ;
        RECT -17.190 21.250 -16.310 21.420 ;
      LAYER met1 ;
        RECT -16.050 26.240 -15.790 26.560 ;
        RECT -16.045 25.900 -15.795 26.240 ;
        RECT -15.350 25.900 -15.050 26.000 ;
        RECT -16.700 25.830 -15.050 25.900 ;
        RECT -17.200 25.650 -15.050 25.830 ;
        RECT -17.200 25.600 -16.200 25.650 ;
        RECT -15.350 25.550 -15.050 25.650 ;
        RECT -15.300 24.650 -15.000 24.750 ;
        RECT -17.200 24.420 -15.000 24.650 ;
        RECT -16.700 24.400 -15.000 24.420 ;
        RECT -16.125 22.700 -15.875 24.400 ;
        RECT -15.300 24.300 -15.000 24.400 ;
        RECT -16.650 22.630 -14.350 22.700 ;
        RECT -17.250 22.450 -14.350 22.630 ;
        RECT -17.250 22.400 -16.250 22.450 ;
        RECT -17.250 21.400 -16.250 21.450 ;
        RECT -14.600 21.400 -14.350 22.450 ;
        RECT -17.250 21.220 -14.350 21.400 ;
        RECT -16.700 21.150 -14.350 21.220 ;
      LAYER via ;
        RECT -16.050 26.270 -15.790 26.530 ;
      LAYER met2 ;
        RECT -32.000 38.400 -31.400 42.450 ;
        RECT -31.830 35.980 -31.530 38.400 ;
        RECT -31.865 35.700 -31.495 35.980 ;
        RECT -31.830 35.690 -31.530 35.700 ;
        RECT -16.160 26.080 -15.680 26.640 ;
      LAYER via2 ;
        RECT -31.820 35.700 -31.540 35.980 ;
        RECT -16.070 26.250 -15.770 26.550 ;
      LAYER met3 ;
        RECT -31.845 35.990 -31.515 36.005 ;
        RECT -31.845 35.690 -15.770 35.990 ;
        RECT -31.845 35.675 -31.515 35.690 ;
        RECT -16.070 26.640 -15.770 35.690 ;
        RECT -16.160 26.080 -15.680 26.640 ;
    END
  END PD2
  PIN pd2_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT -17.750 22.385 -17.450 22.450 ;
        RECT -17.750 22.055 -17.440 22.385 ;
        RECT -17.750 21.795 -17.450 22.055 ;
        RECT -17.750 21.465 -17.440 21.795 ;
        RECT -17.750 21.450 -17.450 21.465 ;
      LAYER mcon ;
        RECT -17.700 21.600 -17.500 22.300 ;
      LAYER met1 ;
        RECT -26.950 26.550 -19.150 26.850 ;
        RECT -26.950 23.850 -26.650 26.550 ;
        RECT -27.380 23.550 -26.650 23.850 ;
        RECT -19.450 21.950 -19.150 26.550 ;
        RECT -17.750 21.950 -17.450 22.450 ;
        RECT -19.450 21.650 -17.450 21.950 ;
        RECT -17.750 21.450 -17.450 21.650 ;
      LAYER via ;
        RECT -27.350 23.550 -27.050 23.850 ;
      LAYER met2 ;
        RECT -27.350 -42.950 -27.050 23.880 ;
        RECT -27.350 -43.250 3.750 -42.950 ;
        RECT 3.450 -65.350 3.750 -43.250 ;
        RECT 3.450 -65.650 10.450 -65.350 ;
        RECT 10.150 -68.300 10.450 -65.650 ;
        RECT 10.000 -68.350 10.450 -68.300 ;
        RECT 10.000 -72.350 10.600 -68.350 ;
    END
  END pd2_a
  PIN pd2_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT -17.700 25.585 -17.400 25.650 ;
        RECT -17.700 25.255 -17.390 25.585 ;
        RECT -17.700 24.995 -17.400 25.255 ;
        RECT -17.700 24.665 -17.390 24.995 ;
        RECT -17.700 24.650 -17.400 24.665 ;
      LAYER mcon ;
        RECT -17.650 24.800 -17.450 25.500 ;
      LAYER met1 ;
        RECT -27.550 27.150 -17.450 27.450 ;
        RECT -27.550 24.350 -27.250 27.150 ;
        RECT -17.750 25.650 -17.450 27.150 ;
        RECT -17.750 24.650 -17.400 25.650 ;
        RECT -27.980 24.050 -27.250 24.350 ;
      LAYER via ;
        RECT -27.950 24.050 -27.650 24.350 ;
      LAYER met2 ;
        RECT -27.950 -43.550 -27.650 24.380 ;
        RECT -27.950 -43.850 3.250 -43.550 ;
        RECT 2.950 -65.850 3.250 -43.850 ;
        RECT 2.950 -66.150 5.450 -65.850 ;
        RECT 5.150 -68.300 5.450 -66.150 ;
        RECT 5.000 -72.350 5.600 -68.300 ;
    END
  END pd2_b
  PIN PD3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT -10.770 25.630 -9.730 25.800 ;
        RECT -8.900 25.550 -8.600 26.000 ;
        RECT -8.800 24.750 -8.600 25.550 ;
        RECT -10.770 24.450 -9.730 24.620 ;
        RECT -8.850 24.300 -8.550 24.750 ;
        RECT -10.770 22.430 -9.730 22.600 ;
        RECT -10.770 21.250 -9.730 21.420 ;
      LAYER mcon ;
        RECT -10.690 25.630 -9.810 25.800 ;
        RECT -8.850 25.650 -8.650 25.900 ;
        RECT -10.690 24.450 -9.810 24.620 ;
        RECT -8.800 24.400 -8.600 24.650 ;
        RECT -10.690 22.430 -9.810 22.600 ;
        RECT -10.690 21.250 -9.810 21.420 ;
      LAYER met1 ;
        RECT -9.650 27.120 -9.390 27.440 ;
        RECT -9.645 25.900 -9.395 27.120 ;
        RECT -8.900 25.900 -8.600 26.000 ;
        RECT -10.250 25.830 -8.600 25.900 ;
        RECT -10.750 25.650 -8.600 25.830 ;
        RECT -10.750 25.600 -9.750 25.650 ;
        RECT -8.900 25.550 -8.600 25.650 ;
        RECT -8.850 24.650 -8.550 24.750 ;
        RECT -10.750 24.420 -8.550 24.650 ;
        RECT -10.250 24.400 -8.550 24.420 ;
        RECT -9.680 22.700 -9.360 24.400 ;
        RECT -8.850 24.300 -8.550 24.400 ;
        RECT -10.150 22.630 -7.850 22.700 ;
        RECT -10.750 22.450 -7.850 22.630 ;
        RECT -10.750 22.400 -9.750 22.450 ;
        RECT -10.750 21.400 -9.750 21.450 ;
        RECT -8.100 21.400 -7.850 22.450 ;
        RECT -10.750 21.220 -7.850 21.400 ;
        RECT -10.200 21.150 -7.850 21.220 ;
      LAYER via ;
        RECT -9.650 27.150 -9.390 27.410 ;
      LAYER met2 ;
        RECT -24.000 38.400 -23.400 42.450 ;
        RECT -23.910 36.860 -23.610 38.400 ;
        RECT -23.945 36.580 -23.575 36.860 ;
        RECT -23.910 36.570 -23.610 36.580 ;
        RECT -9.760 27.120 -9.280 27.520 ;
      LAYER via2 ;
        RECT -23.900 36.580 -23.620 36.860 ;
        RECT -9.670 27.130 -9.370 27.430 ;
      LAYER met3 ;
        RECT -23.925 36.870 -23.595 36.885 ;
        RECT -23.925 36.570 -9.370 36.870 ;
        RECT -23.925 36.555 -23.595 36.570 ;
        RECT -9.670 27.520 -9.370 36.570 ;
        RECT -9.760 27.120 -9.280 27.520 ;
        RECT -9.695 27.105 -9.345 27.120 ;
    END
  END PD3
  PIN pd3_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT -11.250 22.385 -10.950 22.450 ;
        RECT -11.250 22.055 -10.940 22.385 ;
        RECT -11.250 21.795 -10.950 22.055 ;
        RECT -11.250 21.465 -10.940 21.795 ;
        RECT -11.250 21.450 -10.950 21.465 ;
      LAYER mcon ;
        RECT -11.200 21.600 -11.000 22.300 ;
      LAYER met1 ;
        RECT -28.150 27.650 -12.750 27.950 ;
        RECT -28.150 24.850 -27.850 27.650 ;
        RECT -28.480 24.550 -27.850 24.850 ;
        RECT -13.050 22.050 -12.750 27.650 ;
        RECT -11.250 22.050 -10.950 22.450 ;
        RECT -13.050 21.750 -10.950 22.050 ;
        RECT -11.250 21.450 -10.950 21.750 ;
      LAYER via ;
        RECT -28.450 24.550 -28.150 24.850 ;
      LAYER met2 ;
        RECT -28.450 -44.050 -28.150 24.880 ;
        RECT -28.450 -44.350 0.450 -44.050 ;
        RECT 0.150 -68.300 0.450 -44.350 ;
        RECT 0.000 -72.350 0.600 -68.300 ;
    END
  END pd3_a
  PIN pd3_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT -11.250 25.585 -10.950 25.650 ;
        RECT -11.250 25.255 -10.940 25.585 ;
        RECT -11.250 24.995 -10.950 25.255 ;
        RECT -11.250 24.665 -10.940 24.995 ;
        RECT -11.250 24.650 -10.950 24.665 ;
      LAYER mcon ;
        RECT -11.200 24.800 -11.000 25.500 ;
      LAYER met1 ;
        RECT -28.750 28.250 -11.050 28.550 ;
        RECT -28.750 25.450 -28.450 28.250 ;
        RECT -28.980 25.150 -28.450 25.450 ;
        RECT -11.350 25.650 -11.050 28.250 ;
        RECT -11.350 24.750 -10.950 25.650 ;
        RECT -11.250 24.650 -10.950 24.750 ;
      LAYER via ;
        RECT -28.950 25.150 -28.650 25.450 ;
      LAYER met2 ;
        RECT -28.950 -44.650 -28.650 25.480 ;
        RECT -28.950 -44.950 -4.550 -44.650 ;
        RECT -4.850 -68.300 -4.550 -44.950 ;
        RECT -5.000 -72.350 -4.400 -68.300 ;
    END
  END pd3_b
  PIN PD4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT -4.320 25.630 -3.280 25.800 ;
        RECT -2.450 25.550 -2.150 26.000 ;
        RECT -2.350 24.750 -2.150 25.550 ;
        RECT -4.320 24.450 -3.280 24.620 ;
        RECT -2.400 24.300 -2.100 24.750 ;
        RECT -4.370 22.430 -3.330 22.600 ;
        RECT -4.370 21.250 -3.330 21.420 ;
      LAYER mcon ;
        RECT -4.240 25.630 -3.360 25.800 ;
        RECT -2.400 25.650 -2.200 25.900 ;
        RECT -4.240 24.450 -3.360 24.620 ;
        RECT -2.350 24.400 -2.150 24.650 ;
        RECT -4.290 22.430 -3.410 22.600 ;
        RECT -4.290 21.250 -3.410 21.420 ;
      LAYER met1 ;
        RECT -3.250 27.680 -2.990 28.000 ;
        RECT -3.245 25.900 -2.995 27.680 ;
        RECT -2.450 25.900 -2.150 26.000 ;
        RECT -3.800 25.830 -2.150 25.900 ;
        RECT -4.300 25.650 -2.150 25.830 ;
        RECT -4.300 25.600 -3.300 25.650 ;
        RECT -2.450 25.550 -2.150 25.650 ;
        RECT -2.400 24.650 -2.100 24.750 ;
        RECT -4.300 24.420 -2.100 24.650 ;
        RECT -3.800 24.400 -2.100 24.420 ;
        RECT -3.200 22.700 -2.880 24.400 ;
        RECT -2.400 24.300 -2.100 24.400 ;
        RECT -3.750 22.630 -1.450 22.700 ;
        RECT -4.350 22.450 -1.450 22.630 ;
        RECT -4.350 22.400 -3.350 22.450 ;
        RECT -4.350 21.400 -3.350 21.450 ;
        RECT -1.700 21.400 -1.450 22.450 ;
        RECT -4.350 21.220 -1.450 21.400 ;
        RECT -3.800 21.150 -1.450 21.220 ;
      LAYER via ;
        RECT -3.250 27.710 -2.990 27.970 ;
      LAYER met2 ;
        RECT -16.000 38.400 -15.400 42.450 ;
        RECT -15.910 36.870 -15.610 38.400 ;
        RECT -3.260 36.870 -2.980 36.905 ;
        RECT -15.910 36.570 -2.970 36.870 ;
        RECT -3.260 36.535 -2.980 36.570 ;
        RECT -3.360 27.600 -2.880 28.080 ;
      LAYER via2 ;
        RECT -3.260 36.580 -2.980 36.860 ;
        RECT -3.270 27.690 -2.970 28.000 ;
      LAYER met3 ;
        RECT -3.285 36.555 -2.955 36.885 ;
        RECT -3.270 28.080 -2.970 36.555 ;
        RECT -3.360 27.600 -2.880 28.080 ;
    END
  END PD4
  PIN pd4_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT -4.850 22.385 -4.550 22.450 ;
        RECT -4.850 22.055 -4.540 22.385 ;
        RECT -4.850 21.795 -4.550 22.055 ;
        RECT -4.850 21.465 -4.540 21.795 ;
        RECT -4.850 21.450 -4.550 21.465 ;
      LAYER mcon ;
        RECT -4.800 21.600 -4.600 22.300 ;
      LAYER met1 ;
        RECT -29.250 28.850 -6.150 29.150 ;
        RECT -29.250 25.950 -28.950 28.850 ;
        RECT -29.580 25.650 -28.950 25.950 ;
        RECT -6.450 22.050 -6.150 28.850 ;
        RECT -4.850 22.050 -4.550 22.450 ;
        RECT -6.450 21.750 -4.550 22.050 ;
        RECT -4.850 21.450 -4.550 21.750 ;
      LAYER via ;
        RECT -29.550 25.650 -29.250 25.950 ;
      LAYER met2 ;
        RECT -29.550 -45.150 -29.250 25.980 ;
        RECT -29.550 -45.450 -9.550 -45.150 ;
        RECT -9.850 -68.300 -9.550 -45.450 ;
        RECT -10.000 -72.350 -9.400 -68.300 ;
    END
  END pd4_a
  PIN pd4_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT -4.800 25.585 -4.500 25.650 ;
        RECT -4.800 25.255 -4.490 25.585 ;
        RECT -4.800 24.995 -4.500 25.255 ;
        RECT -4.800 24.665 -4.490 24.995 ;
        RECT -4.800 24.650 -4.500 24.665 ;
      LAYER mcon ;
        RECT -4.750 24.800 -4.550 25.500 ;
      LAYER met1 ;
        RECT -29.750 29.450 -4.650 29.750 ;
        RECT -29.750 26.450 -29.450 29.450 ;
        RECT -30.080 26.150 -29.450 26.450 ;
        RECT -4.950 25.650 -4.650 29.450 ;
        RECT -4.950 24.650 -4.500 25.650 ;
      LAYER via ;
        RECT -30.050 26.150 -29.750 26.450 ;
      LAYER met2 ;
        RECT -30.050 -45.650 -29.750 26.480 ;
        RECT -30.050 -45.950 -14.550 -45.650 ;
        RECT -14.850 -68.300 -14.550 -45.950 ;
        RECT -15.000 -72.350 -14.400 -68.300 ;
    END
  END pd4_b
  PIN PD5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 2.130 25.630 3.170 25.800 ;
        RECT 4.000 25.550 4.300 26.000 ;
        RECT 4.100 24.750 4.300 25.550 ;
        RECT 2.130 24.450 3.170 24.620 ;
        RECT 4.050 24.300 4.350 24.750 ;
        RECT 2.130 22.430 3.170 22.600 ;
        RECT 2.130 21.250 3.170 21.420 ;
      LAYER mcon ;
        RECT 2.210 25.630 3.090 25.800 ;
        RECT 4.050 25.650 4.250 25.900 ;
        RECT 2.210 24.450 3.090 24.620 ;
        RECT 4.100 24.400 4.300 24.650 ;
        RECT 2.210 22.430 3.090 22.600 ;
        RECT 2.210 21.250 3.090 21.420 ;
      LAYER met1 ;
        RECT 3.200 26.750 3.520 27.010 ;
        RECT 3.235 25.900 3.485 26.750 ;
        RECT 4.000 25.900 4.300 26.000 ;
        RECT 2.650 25.830 4.300 25.900 ;
        RECT 2.150 25.650 4.300 25.830 ;
        RECT 2.150 25.600 3.150 25.650 ;
        RECT 4.000 25.550 4.300 25.650 ;
        RECT 4.050 24.650 4.350 24.750 ;
        RECT 2.150 24.420 4.350 24.650 ;
        RECT 2.650 24.400 4.350 24.420 ;
        RECT 3.440 22.700 3.760 24.400 ;
        RECT 4.050 24.300 4.350 24.400 ;
        RECT 2.750 22.630 5.050 22.700 ;
        RECT 2.150 22.450 5.050 22.630 ;
        RECT 2.150 22.400 3.150 22.450 ;
        RECT 2.150 21.400 3.150 21.450 ;
        RECT 4.800 21.400 5.050 22.450 ;
        RECT 2.150 21.220 5.050 21.400 ;
        RECT 2.700 21.150 5.050 21.220 ;
      LAYER via ;
        RECT 3.230 26.750 3.490 27.010 ;
      LAYER met2 ;
        RECT -8.000 38.400 -7.400 42.450 ;
        RECT -7.830 37.900 -7.530 38.400 ;
        RECT -7.865 37.620 -7.495 37.900 ;
        RECT -7.830 37.610 -7.530 37.620 ;
        RECT 3.230 27.030 3.490 27.040 ;
        RECT 3.165 26.730 3.555 27.030 ;
        RECT 3.230 26.720 3.490 26.730 ;
      LAYER via2 ;
        RECT -7.820 37.620 -7.540 37.900 ;
        RECT 3.210 26.730 3.510 27.030 ;
      LAYER met3 ;
        RECT -7.845 37.595 -7.515 37.925 ;
        RECT -7.830 27.030 -7.530 37.595 ;
        RECT 3.185 27.030 3.535 27.055 ;
        RECT -7.830 26.730 3.535 27.030 ;
        RECT 3.185 26.705 3.535 26.730 ;
    END
  END PD5
  PIN pd5_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 1.650 22.385 1.950 22.450 ;
        RECT 1.650 22.055 1.960 22.385 ;
        RECT 1.650 21.795 1.950 22.055 ;
        RECT 1.650 21.465 1.960 21.795 ;
        RECT 1.650 21.450 1.950 21.465 ;
      LAYER mcon ;
        RECT 1.700 21.600 1.900 22.300 ;
      LAYER met1 ;
        RECT -30.350 30.050 0.350 30.350 ;
        RECT -30.350 26.950 -30.050 30.050 ;
        RECT -30.680 26.650 -30.050 26.950 ;
        RECT 0.050 22.150 0.350 30.050 ;
        RECT 1.650 22.150 1.950 22.450 ;
        RECT 0.050 21.850 1.950 22.150 ;
        RECT 1.650 21.450 1.950 21.850 ;
      LAYER via ;
        RECT -30.650 26.650 -30.350 26.950 ;
      LAYER met2 ;
        RECT -30.650 -46.150 -30.350 26.980 ;
        RECT -30.650 -46.450 -19.550 -46.150 ;
        RECT -19.850 -68.300 -19.550 -46.450 ;
        RECT -20.000 -68.350 -19.550 -68.300 ;
        RECT -20.000 -72.350 -19.400 -68.350 ;
    END
  END pd5_a
  PIN pd5_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 1.650 25.585 1.950 25.650 ;
        RECT 1.650 25.255 1.960 25.585 ;
        RECT 1.650 24.995 1.950 25.255 ;
        RECT 1.650 24.665 1.960 24.995 ;
        RECT 1.650 24.650 1.950 24.665 ;
      LAYER mcon ;
        RECT 1.700 24.800 1.900 25.500 ;
      LAYER met1 ;
        RECT -30.950 30.550 1.850 30.850 ;
        RECT -30.950 27.580 -30.650 30.550 ;
        RECT -31.250 27.250 -30.650 27.580 ;
        RECT -31.250 27.220 -30.950 27.250 ;
        RECT 1.550 25.650 1.850 30.550 ;
        RECT 1.550 24.650 1.950 25.650 ;
      LAYER met2 ;
        RECT -31.280 27.250 -30.920 27.550 ;
        RECT -31.250 -46.650 -30.950 27.250 ;
        RECT -31.250 -46.950 -24.550 -46.650 ;
        RECT -24.850 -68.300 -24.550 -46.950 ;
        RECT -25.000 -72.350 -24.400 -68.300 ;
    END
  END pd5_b
  PIN PD6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 8.580 25.630 9.620 25.800 ;
        RECT 10.450 25.550 10.750 26.000 ;
        RECT 10.550 24.750 10.750 25.550 ;
        RECT 8.580 24.450 9.620 24.620 ;
        RECT 10.500 24.300 10.800 24.750 ;
        RECT 8.530 22.430 9.570 22.600 ;
        RECT 8.530 21.250 9.570 21.420 ;
      LAYER mcon ;
        RECT 8.660 25.630 9.540 25.800 ;
        RECT 10.500 25.650 10.700 25.900 ;
        RECT 8.660 24.450 9.540 24.620 ;
        RECT 10.550 24.400 10.750 24.650 ;
        RECT 8.610 22.430 9.490 22.600 ;
        RECT 8.610 21.250 9.490 21.420 ;
      LAYER met1 ;
        RECT 9.630 27.520 9.890 27.840 ;
        RECT 9.635 25.900 9.885 27.520 ;
        RECT 10.450 25.900 10.750 26.000 ;
        RECT 9.100 25.830 10.750 25.900 ;
        RECT 8.600 25.650 10.750 25.830 ;
        RECT 8.600 25.600 9.600 25.650 ;
        RECT 10.450 25.550 10.750 25.650 ;
        RECT 10.500 24.650 10.800 24.750 ;
        RECT 8.600 24.420 10.800 24.650 ;
        RECT 9.100 24.400 10.800 24.420 ;
        RECT 9.920 22.700 10.240 24.400 ;
        RECT 10.500 24.300 10.800 24.400 ;
        RECT 9.150 22.630 11.450 22.700 ;
        RECT 8.550 22.450 11.450 22.630 ;
        RECT 8.550 22.400 9.550 22.450 ;
        RECT 8.550 21.400 9.550 21.450 ;
        RECT 11.200 21.400 11.450 22.450 ;
        RECT 8.550 21.220 11.450 21.400 ;
        RECT 9.100 21.150 11.450 21.220 ;
      LAYER via ;
        RECT 9.630 27.550 9.890 27.810 ;
      LAYER met2 ;
        RECT 0.000 38.400 0.600 42.450 ;
        RECT 0.170 38.220 0.470 38.400 ;
        RECT 0.135 37.940 0.505 38.220 ;
        RECT 0.170 37.930 0.470 37.940 ;
        RECT 9.520 27.440 10.000 27.920 ;
      LAYER via2 ;
        RECT 0.180 37.940 0.460 38.220 ;
        RECT 9.610 27.530 9.910 27.830 ;
      LAYER met3 ;
        RECT 0.155 37.915 0.485 38.245 ;
        RECT 0.170 27.830 0.470 37.915 ;
        RECT 9.520 27.830 10.000 27.920 ;
        RECT 0.170 27.530 10.000 27.830 ;
        RECT 9.520 27.440 10.000 27.530 ;
    END
  END PD6
  PIN pd6_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 8.050 22.385 8.350 22.450 ;
        RECT 8.050 22.055 8.360 22.385 ;
        RECT 8.050 21.795 8.350 22.055 ;
        RECT 8.050 21.465 8.360 21.795 ;
        RECT 8.050 21.450 8.350 21.465 ;
      LAYER mcon ;
        RECT 8.100 21.600 8.300 22.300 ;
      LAYER met1 ;
        RECT -31.450 31.050 6.750 31.350 ;
        RECT -31.450 28.250 -31.150 31.050 ;
        RECT -31.780 27.950 -31.150 28.250 ;
        RECT 6.450 22.050 6.750 31.050 ;
        RECT 8.050 22.050 8.350 22.450 ;
        RECT 6.450 21.750 8.350 22.050 ;
        RECT 8.050 21.450 8.350 21.750 ;
      LAYER via ;
        RECT -31.750 27.950 -31.450 28.250 ;
      LAYER met2 ;
        RECT -31.750 -47.250 -31.450 28.280 ;
        RECT -31.750 -47.550 -29.550 -47.250 ;
        RECT -29.850 -68.300 -29.550 -47.550 ;
        RECT -30.000 -72.350 -29.400 -68.300 ;
    END
  END pd6_a
  PIN pd6_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 8.100 25.585 8.400 25.650 ;
        RECT 8.100 25.255 8.410 25.585 ;
        RECT 8.100 24.995 8.400 25.255 ;
        RECT 8.100 24.665 8.410 24.995 ;
        RECT 8.100 24.650 8.400 24.665 ;
      LAYER mcon ;
        RECT 8.150 24.800 8.350 25.500 ;
      LAYER met1 ;
        RECT -32.050 31.650 8.250 31.950 ;
        RECT -32.050 28.750 -31.750 31.650 ;
        RECT -32.380 28.450 -31.750 28.750 ;
        RECT 7.950 25.650 8.250 31.650 ;
        RECT 7.950 24.650 8.400 25.650 ;
      LAYER via ;
        RECT -32.350 28.450 -32.050 28.750 ;
      LAYER met2 ;
        RECT -32.350 -47.250 -32.050 28.780 ;
        RECT -34.850 -47.550 -32.050 -47.250 ;
        RECT -34.850 -68.300 -34.550 -47.550 ;
        RECT -35.000 -72.350 -34.400 -68.300 ;
    END
  END pd6_b
  PIN PD7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 15.030 25.630 16.070 25.800 ;
        RECT 16.900 25.550 17.200 26.000 ;
        RECT 17.000 24.750 17.200 25.550 ;
        RECT 15.030 24.450 16.070 24.620 ;
        RECT 16.950 24.300 17.250 24.750 ;
        RECT 15.030 22.430 16.070 22.600 ;
        RECT 15.030 21.250 16.070 21.420 ;
      LAYER mcon ;
        RECT 15.110 25.630 15.990 25.800 ;
        RECT 16.950 25.650 17.150 25.900 ;
        RECT 15.110 24.450 15.990 24.620 ;
        RECT 17.000 24.400 17.200 24.650 ;
        RECT 15.110 22.430 15.990 22.600 ;
        RECT 15.110 21.250 15.990 21.420 ;
      LAYER met1 ;
        RECT 16.190 28.400 16.450 28.720 ;
        RECT 16.195 25.900 16.445 28.400 ;
        RECT 16.900 25.900 17.200 26.000 ;
        RECT 15.550 25.830 17.200 25.900 ;
        RECT 15.050 25.650 17.200 25.830 ;
        RECT 15.050 25.600 16.050 25.650 ;
        RECT 16.900 25.550 17.200 25.650 ;
        RECT 16.950 24.650 17.250 24.750 ;
        RECT 15.050 24.420 17.250 24.650 ;
        RECT 15.550 24.400 17.250 24.420 ;
        RECT 16.320 22.700 16.640 24.400 ;
        RECT 16.950 24.300 17.250 24.400 ;
        RECT 15.650 22.630 17.950 22.700 ;
        RECT 15.050 22.450 17.950 22.630 ;
        RECT 15.050 22.400 16.050 22.450 ;
        RECT 15.050 21.400 16.050 21.450 ;
        RECT 17.700 21.400 17.950 22.450 ;
        RECT 15.050 21.220 17.950 21.400 ;
        RECT 15.600 21.150 17.950 21.220 ;
      LAYER via ;
        RECT 16.190 28.430 16.450 28.690 ;
      LAYER met2 ;
        RECT 8.000 38.400 8.600 42.450 ;
        RECT 8.170 38.140 8.470 38.400 ;
        RECT 8.135 37.860 8.505 38.140 ;
        RECT 8.170 37.850 8.470 37.860 ;
        RECT 16.080 28.320 16.560 28.800 ;
      LAYER via2 ;
        RECT 8.180 37.860 8.460 38.140 ;
        RECT 16.170 28.410 16.470 28.710 ;
      LAYER met3 ;
        RECT 8.155 37.835 8.485 38.165 ;
        RECT 8.170 28.710 8.470 37.835 ;
        RECT 16.080 28.710 16.560 28.800 ;
        RECT 8.170 28.410 16.560 28.710 ;
        RECT 16.080 28.320 16.560 28.410 ;
    END
  END PD7
  PIN pd7_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 14.550 22.385 14.850 22.450 ;
        RECT 14.550 22.055 14.860 22.385 ;
        RECT 14.550 21.795 14.850 22.055 ;
        RECT 14.550 21.465 14.860 21.795 ;
        RECT 14.550 21.450 14.850 21.465 ;
      LAYER mcon ;
        RECT 14.600 21.600 14.800 22.300 ;
      LAYER met1 ;
        RECT -32.550 32.250 13.150 32.550 ;
        RECT -32.550 29.250 -32.250 32.250 ;
        RECT -32.980 28.950 -32.250 29.250 ;
        RECT 12.850 22.050 13.150 32.250 ;
        RECT 14.550 22.050 14.850 22.450 ;
        RECT 12.850 21.750 14.850 22.050 ;
        RECT 14.550 21.450 14.850 21.750 ;
      LAYER via ;
        RECT -32.950 28.950 -32.650 29.250 ;
      LAYER met2 ;
        RECT -32.950 -46.750 -32.650 29.280 ;
        RECT -37.150 -47.050 -32.650 -46.750 ;
        RECT -37.150 -63.250 -36.850 -47.050 ;
        RECT -39.850 -63.550 -36.850 -63.250 ;
        RECT -39.850 -68.300 -39.550 -63.550 ;
        RECT -40.000 -72.350 -39.400 -68.300 ;
    END
  END pd7_a
  PIN pd7_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 14.550 25.585 14.850 25.650 ;
        RECT 14.550 25.255 14.860 25.585 ;
        RECT 14.550 24.995 14.850 25.255 ;
        RECT 14.550 24.665 14.860 24.995 ;
        RECT 14.550 24.650 14.850 24.665 ;
      LAYER mcon ;
        RECT 14.600 24.800 14.800 25.500 ;
      LAYER met1 ;
        RECT -33.150 32.750 14.650 33.050 ;
        RECT -33.150 29.750 -32.850 32.750 ;
        RECT -33.680 29.450 -32.850 29.750 ;
        RECT 14.350 25.650 14.650 32.750 ;
        RECT 14.350 24.650 14.850 25.650 ;
      LAYER via ;
        RECT -33.650 29.450 -33.350 29.750 ;
      LAYER met2 ;
        RECT -33.650 -46.250 -33.350 29.780 ;
        RECT -37.750 -46.550 -33.350 -46.250 ;
        RECT -37.750 -62.650 -37.450 -46.550 ;
        RECT -44.850 -62.950 -37.450 -62.650 ;
        RECT -44.850 -68.300 -44.550 -62.950 ;
        RECT -45.000 -72.350 -44.400 -68.300 ;
    END
  END pd7_b
  PIN PD8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 21.480 25.630 22.520 25.800 ;
        RECT 23.350 25.550 23.650 26.000 ;
        RECT 23.450 24.750 23.650 25.550 ;
        RECT 21.480 24.450 22.520 24.620 ;
        RECT 23.400 24.300 23.700 24.750 ;
        RECT 21.430 22.430 22.470 22.600 ;
        RECT 21.430 21.250 22.470 21.420 ;
      LAYER mcon ;
        RECT 21.560 25.630 22.440 25.800 ;
        RECT 23.400 25.650 23.600 25.900 ;
        RECT 21.560 24.450 22.440 24.620 ;
        RECT 23.450 24.400 23.650 24.650 ;
        RECT 21.510 22.430 22.390 22.600 ;
        RECT 21.510 21.250 22.390 21.420 ;
      LAYER met1 ;
        RECT 22.670 29.600 22.930 29.920 ;
        RECT 22.675 25.900 22.925 29.600 ;
        RECT 23.350 25.900 23.650 26.000 ;
        RECT 22.000 25.830 23.650 25.900 ;
        RECT 21.500 25.650 23.650 25.830 ;
        RECT 21.500 25.600 22.500 25.650 ;
        RECT 23.350 25.550 23.650 25.650 ;
        RECT 23.400 24.650 23.700 24.750 ;
        RECT 21.500 24.420 23.700 24.650 ;
        RECT 22.000 24.400 23.700 24.420 ;
        RECT 22.880 22.700 23.200 24.400 ;
        RECT 23.400 24.300 23.700 24.400 ;
        RECT 22.050 22.630 24.350 22.700 ;
        RECT 21.450 22.450 24.350 22.630 ;
        RECT 21.450 22.400 22.450 22.450 ;
        RECT 21.450 21.400 22.450 21.450 ;
        RECT 24.100 21.400 24.350 22.450 ;
        RECT 21.450 21.220 24.350 21.400 ;
        RECT 22.000 21.150 24.350 21.220 ;
      LAYER via ;
        RECT 22.670 29.630 22.930 29.890 ;
      LAYER met2 ;
        RECT 16.000 38.400 16.600 42.450 ;
        RECT 16.170 38.140 16.470 38.400 ;
        RECT 16.135 37.860 16.505 38.140 ;
        RECT 16.170 37.850 16.470 37.860 ;
        RECT 22.560 29.520 23.040 30.000 ;
      LAYER via2 ;
        RECT 16.180 37.860 16.460 38.140 ;
        RECT 22.650 29.610 22.950 29.910 ;
      LAYER met3 ;
        RECT 16.155 37.835 16.485 38.165 ;
        RECT 16.170 29.910 16.470 37.835 ;
        RECT 22.560 29.910 23.040 30.000 ;
        RECT 16.170 29.610 23.040 29.910 ;
        RECT 22.560 29.520 23.040 29.610 ;
    END
  END PD8
  PIN pd8_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 20.950 22.385 21.250 22.450 ;
        RECT 20.950 22.055 21.260 22.385 ;
        RECT 20.950 21.795 21.250 22.055 ;
        RECT 20.950 21.465 21.260 21.795 ;
        RECT 20.950 21.450 21.250 21.465 ;
      LAYER mcon ;
        RECT 21.000 21.600 21.200 22.300 ;
      LAYER met1 ;
        RECT -33.750 33.250 19.750 33.550 ;
        RECT -33.750 30.250 -33.450 33.250 ;
        RECT -34.280 29.950 -33.450 30.250 ;
        RECT 19.450 22.050 19.750 33.250 ;
        RECT 20.950 22.050 21.250 22.450 ;
        RECT 19.450 21.750 21.250 22.050 ;
        RECT 20.950 21.450 21.250 21.750 ;
      LAYER via ;
        RECT -34.250 29.950 -33.950 30.250 ;
      LAYER met2 ;
        RECT -34.250 -45.650 -33.950 30.280 ;
        RECT -38.250 -45.950 -33.950 -45.650 ;
        RECT -38.250 -62.150 -37.950 -45.950 ;
        RECT -49.850 -62.450 -37.950 -62.150 ;
        RECT -49.850 -68.300 -49.550 -62.450 ;
        RECT -50.000 -72.350 -49.400 -68.300 ;
    END
  END pd8_a
  PIN pd8_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 21.000 25.585 21.300 25.650 ;
        RECT 21.000 25.255 21.310 25.585 ;
        RECT 21.000 24.995 21.300 25.255 ;
        RECT 21.000 24.665 21.310 24.995 ;
        RECT 21.000 24.650 21.300 24.665 ;
      LAYER mcon ;
        RECT 21.050 24.800 21.250 25.500 ;
      LAYER met1 ;
        RECT 20.850 26.880 21.230 27.200 ;
        RECT 20.880 25.650 21.200 26.880 ;
        RECT 20.880 24.800 21.300 25.650 ;
        RECT 21.000 24.650 21.300 24.800 ;
      LAYER via ;
        RECT 20.880 26.880 21.200 27.200 ;
      LAYER met2 ;
        RECT -25.180 29.600 -24.900 29.625 ;
        RECT -25.200 29.280 21.200 29.600 ;
        RECT -25.180 29.255 -24.900 29.280 ;
        RECT 20.880 26.850 21.200 29.280 ;
        RECT -54.800 -67.600 -51.635 -67.280 ;
        RECT -54.800 -68.400 -54.480 -67.600 ;
        RECT -54.960 -72.400 -54.320 -68.400 ;
      LAYER via2 ;
        RECT -25.180 29.300 -24.900 29.580 ;
        RECT -52.000 -67.600 -51.680 -67.280 ;
      LAYER met3 ;
        RECT -25.205 29.600 -24.875 29.605 ;
        RECT -48.480 29.280 -24.875 29.600 ;
        RECT -52.025 -67.280 -51.655 -67.255 ;
        RECT -48.480 -67.280 -48.160 29.280 ;
        RECT -25.205 29.275 -24.875 29.280 ;
        RECT -52.025 -67.600 -48.160 -67.280 ;
        RECT -52.025 -67.625 -51.655 -67.600 ;
    END
  END pd8_b
  PIN PD9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 27.930 25.630 28.970 25.800 ;
        RECT 29.800 25.550 30.100 26.000 ;
        RECT 29.900 24.750 30.100 25.550 ;
        RECT 27.930 24.450 28.970 24.620 ;
        RECT 29.850 24.300 30.150 24.750 ;
        RECT 27.930 22.430 28.970 22.600 ;
        RECT 27.930 21.250 28.970 21.420 ;
      LAYER mcon ;
        RECT 28.010 25.630 28.890 25.800 ;
        RECT 29.850 25.650 30.050 25.900 ;
        RECT 28.010 24.450 28.890 24.620 ;
        RECT 29.900 24.400 30.100 24.650 ;
        RECT 28.010 22.430 28.890 22.600 ;
        RECT 28.010 21.250 28.890 21.420 ;
      LAYER met1 ;
        RECT 29.070 30.640 29.330 30.960 ;
        RECT 29.075 25.900 29.325 30.640 ;
        RECT 29.800 25.900 30.100 26.000 ;
        RECT 28.450 25.830 30.100 25.900 ;
        RECT 27.950 25.650 30.100 25.830 ;
        RECT 27.950 25.600 28.950 25.650 ;
        RECT 29.800 25.550 30.100 25.650 ;
        RECT 29.850 24.650 30.150 24.750 ;
        RECT 27.950 24.420 30.150 24.650 ;
        RECT 28.450 24.400 30.150 24.420 ;
        RECT 29.280 22.700 29.600 24.400 ;
        RECT 29.850 24.300 30.150 24.400 ;
        RECT 28.550 22.630 30.850 22.700 ;
        RECT 27.950 22.450 30.850 22.630 ;
        RECT 27.950 22.400 28.950 22.450 ;
        RECT 27.950 21.400 28.950 21.450 ;
        RECT 30.600 21.400 30.850 22.450 ;
        RECT 27.950 21.220 30.850 21.400 ;
        RECT 28.500 21.150 30.850 21.220 ;
      LAYER via ;
        RECT 29.070 30.670 29.330 30.930 ;
      LAYER met2 ;
        RECT 24.000 38.400 24.600 42.450 ;
        RECT 24.090 38.060 24.390 38.400 ;
        RECT 24.055 37.780 24.425 38.060 ;
        RECT 24.090 37.770 24.390 37.780 ;
        RECT 28.960 30.560 29.440 31.040 ;
      LAYER via2 ;
        RECT 24.100 37.780 24.380 38.060 ;
        RECT 29.050 30.650 29.350 30.950 ;
      LAYER met3 ;
        RECT 24.075 37.755 24.405 38.085 ;
        RECT 24.090 30.950 24.390 37.755 ;
        RECT 28.960 30.950 29.440 31.040 ;
        RECT 24.090 30.650 29.440 30.950 ;
        RECT 28.960 30.560 29.440 30.650 ;
    END
  END PD9
  PIN pd9_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 27.450 22.385 27.750 22.450 ;
        RECT 27.450 22.055 27.760 22.385 ;
        RECT 27.450 21.795 27.750 22.055 ;
        RECT 27.450 21.465 27.760 21.795 ;
        RECT 27.450 21.450 27.750 21.465 ;
      LAYER mcon ;
        RECT 27.500 21.600 27.700 22.300 ;
      LAYER met1 ;
        RECT -34.350 33.750 26.050 34.050 ;
        RECT -34.350 30.750 -34.050 33.750 ;
        RECT -34.880 30.450 -34.050 30.750 ;
        RECT 25.750 22.050 26.050 33.750 ;
        RECT 27.450 22.050 27.750 22.450 ;
        RECT 25.750 21.750 27.750 22.050 ;
        RECT 27.450 21.450 27.750 21.750 ;
      LAYER via ;
        RECT -34.850 30.450 -34.550 30.750 ;
      LAYER met2 ;
        RECT -34.850 -44.950 -34.550 30.780 ;
        RECT -38.950 -45.250 -34.550 -44.950 ;
        RECT -38.950 -61.650 -38.650 -45.250 ;
        RECT -50.750 -61.950 -38.650 -61.650 ;
        RECT -57.350 -65.150 -53.300 -65.000 ;
        RECT -50.750 -65.150 -50.450 -61.950 ;
        RECT -57.350 -65.450 -50.450 -65.150 ;
        RECT -57.350 -65.600 -53.300 -65.450 ;
    END
  END pd9_a
  PIN pd9_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 27.450 25.585 27.750 25.650 ;
        RECT 27.450 25.255 27.760 25.585 ;
        RECT 27.450 24.995 27.750 25.255 ;
        RECT 27.450 24.665 27.760 24.995 ;
        RECT 27.450 24.650 27.750 24.665 ;
      LAYER mcon ;
        RECT 27.500 24.800 27.700 25.500 ;
      LAYER met1 ;
        RECT -34.950 34.250 27.550 34.550 ;
        RECT -34.950 31.250 -34.650 34.250 ;
        RECT -35.480 30.950 -34.650 31.250 ;
        RECT 27.250 25.650 27.550 34.250 ;
        RECT 27.250 24.750 27.750 25.650 ;
        RECT 27.450 24.650 27.750 24.750 ;
      LAYER via ;
        RECT -35.450 30.950 -35.150 31.250 ;
      LAYER met2 ;
        RECT -35.450 -44.150 -35.150 31.280 ;
        RECT -39.550 -44.450 -35.150 -44.150 ;
        RECT -57.350 -60.150 -53.300 -60.000 ;
        RECT -39.550 -60.150 -39.250 -44.450 ;
        RECT -57.350 -60.450 -39.250 -60.150 ;
        RECT -57.350 -60.600 -53.300 -60.450 ;
    END
  END pd9_b
  PIN PD10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 34.380 25.630 35.420 25.800 ;
        RECT 36.250 25.550 36.550 26.000 ;
        RECT 36.350 24.750 36.550 25.550 ;
        RECT 34.380 24.450 35.420 24.620 ;
        RECT 36.300 24.300 36.600 24.750 ;
        RECT 34.330 22.430 35.370 22.600 ;
        RECT 34.330 21.250 35.370 21.420 ;
      LAYER mcon ;
        RECT 34.460 25.630 35.340 25.800 ;
        RECT 36.300 25.650 36.500 25.900 ;
        RECT 34.460 24.450 35.340 24.620 ;
        RECT 36.350 24.400 36.550 24.650 ;
        RECT 34.410 22.430 35.290 22.600 ;
        RECT 34.410 21.250 35.290 21.420 ;
      LAYER met1 ;
        RECT 35.550 27.040 35.810 27.360 ;
        RECT 35.555 25.900 35.805 27.040 ;
        RECT 36.250 25.900 36.550 26.000 ;
        RECT 34.900 25.830 36.550 25.900 ;
        RECT 34.400 25.650 36.550 25.830 ;
        RECT 34.400 25.600 35.400 25.650 ;
        RECT 36.250 25.550 36.550 25.650 ;
        RECT 36.300 24.650 36.600 24.750 ;
        RECT 34.400 24.420 36.600 24.650 ;
        RECT 34.900 24.400 36.600 24.420 ;
        RECT 35.760 22.700 36.080 24.400 ;
        RECT 36.300 24.300 36.600 24.400 ;
        RECT 34.950 22.630 37.250 22.700 ;
        RECT 34.350 22.450 37.250 22.630 ;
        RECT 34.350 22.400 35.350 22.450 ;
        RECT 34.350 21.400 35.350 21.450 ;
        RECT 37.000 21.400 37.250 22.450 ;
        RECT 34.350 21.220 37.250 21.400 ;
        RECT 34.900 21.150 37.250 21.220 ;
      LAYER via ;
        RECT 35.550 27.070 35.810 27.330 ;
      LAYER met2 ;
        RECT 32.000 38.400 32.600 42.450 ;
        RECT 32.170 38.140 32.470 38.400 ;
        RECT 32.135 37.860 32.505 38.140 ;
        RECT 32.170 37.850 32.470 37.860 ;
        RECT 35.440 26.960 35.920 27.440 ;
      LAYER via2 ;
        RECT 32.180 37.860 32.460 38.140 ;
        RECT 35.530 27.050 35.830 27.350 ;
      LAYER met3 ;
        RECT 32.155 37.835 32.485 38.165 ;
        RECT 32.170 35.350 32.470 37.835 ;
        RECT 32.170 35.050 35.830 35.350 ;
        RECT 35.530 27.440 35.830 35.050 ;
        RECT 35.440 26.960 35.920 27.440 ;
    END
  END PD10
  PIN pd10_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 33.850 22.385 34.150 22.450 ;
        RECT 33.850 22.055 34.160 22.385 ;
        RECT 33.850 21.795 34.150 22.055 ;
        RECT 33.850 21.465 34.160 21.795 ;
        RECT 33.850 21.450 34.150 21.465 ;
      LAYER mcon ;
        RECT 33.900 21.600 34.100 22.300 ;
      LAYER met1 ;
        RECT -35.450 34.750 32.550 35.050 ;
        RECT -35.450 31.750 -35.150 34.750 ;
        RECT -36.180 31.450 -35.150 31.750 ;
        RECT 32.250 22.050 32.550 34.750 ;
        RECT 33.850 22.050 34.150 22.450 ;
        RECT 32.250 21.750 34.150 22.050 ;
        RECT 33.850 21.450 34.150 21.750 ;
      LAYER via ;
        RECT -36.150 31.450 -35.850 31.750 ;
      LAYER met2 ;
        RECT -36.150 -43.550 -35.850 31.780 ;
        RECT -40.250 -43.850 -35.850 -43.550 ;
        RECT -57.350 -55.150 -53.300 -55.000 ;
        RECT -40.250 -55.150 -39.950 -43.850 ;
        RECT -57.350 -55.450 -39.950 -55.150 ;
        RECT -57.350 -55.600 -53.300 -55.450 ;
    END
  END pd10_a
  PIN pd10_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 33.900 25.585 34.200 25.650 ;
        RECT 33.900 25.255 34.210 25.585 ;
        RECT 33.900 24.995 34.200 25.255 ;
        RECT 33.900 24.665 34.210 24.995 ;
        RECT 33.900 24.650 34.200 24.665 ;
      LAYER mcon ;
        RECT 33.950 24.800 34.150 25.500 ;
      LAYER met1 ;
        RECT -36.050 35.250 34.050 35.550 ;
        RECT -36.050 32.250 -35.750 35.250 ;
        RECT -36.780 31.950 -35.750 32.250 ;
        RECT 33.750 25.650 34.050 35.250 ;
        RECT 33.750 24.650 34.200 25.650 ;
      LAYER via ;
        RECT -36.750 31.950 -36.450 32.250 ;
      LAYER met2 ;
        RECT -36.750 -42.950 -36.450 32.280 ;
        RECT -40.850 -43.250 -36.450 -42.950 ;
        RECT -57.350 -50.150 -53.300 -50.000 ;
        RECT -40.850 -50.150 -40.550 -43.250 ;
        RECT -57.350 -50.450 -40.550 -50.150 ;
        RECT -57.350 -50.600 -53.300 -50.450 ;
    END
  END pd10_b
  PIN PD11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 40.830 25.630 41.870 25.800 ;
        RECT 42.700 25.550 43.000 26.000 ;
        RECT 42.800 24.750 43.000 25.550 ;
        RECT 40.830 24.450 41.870 24.620 ;
        RECT 42.750 24.300 43.050 24.750 ;
        RECT 40.830 22.430 41.870 22.600 ;
        RECT 40.830 21.250 41.870 21.420 ;
      LAYER mcon ;
        RECT 40.910 25.630 41.790 25.800 ;
        RECT 42.750 25.650 42.950 25.900 ;
        RECT 40.910 24.450 41.790 24.620 ;
        RECT 42.800 24.400 43.000 24.650 ;
        RECT 40.910 22.430 41.790 22.600 ;
        RECT 40.910 21.250 41.790 21.420 ;
      LAYER met1 ;
        RECT 41.950 27.040 42.210 27.360 ;
        RECT 41.955 25.900 42.205 27.040 ;
        RECT 42.700 25.900 43.000 26.000 ;
        RECT 41.350 25.830 43.000 25.900 ;
        RECT 40.850 25.650 43.000 25.830 ;
        RECT 40.850 25.600 41.850 25.650 ;
        RECT 42.700 25.550 43.000 25.650 ;
        RECT 42.750 24.650 43.050 24.750 ;
        RECT 40.850 24.420 43.050 24.650 ;
        RECT 41.350 24.400 43.050 24.420 ;
        RECT 42.240 22.700 42.560 24.400 ;
        RECT 42.750 24.300 43.050 24.400 ;
        RECT 41.450 22.630 43.750 22.700 ;
        RECT 40.850 22.450 43.750 22.630 ;
        RECT 40.850 22.400 41.850 22.450 ;
        RECT 40.850 21.400 41.850 21.450 ;
        RECT 43.500 21.400 43.750 22.450 ;
        RECT 40.850 21.220 43.750 21.400 ;
        RECT 41.400 21.150 43.750 21.220 ;
      LAYER via ;
        RECT 41.950 27.070 42.210 27.330 ;
      LAYER met2 ;
        RECT 40.000 38.400 40.600 42.450 ;
        RECT 40.090 37.850 40.390 38.400 ;
        RECT 40.100 37.815 40.380 37.850 ;
        RECT 41.840 26.960 42.320 27.440 ;
      LAYER via2 ;
        RECT 40.100 37.860 40.380 38.140 ;
        RECT 41.930 27.050 42.230 27.350 ;
      LAYER met3 ;
        RECT 40.075 38.150 40.405 38.165 ;
        RECT 40.075 37.850 42.230 38.150 ;
        RECT 40.075 37.835 40.405 37.850 ;
        RECT 41.930 27.440 42.230 37.850 ;
        RECT 41.840 26.960 42.320 27.440 ;
    END
  END PD11
  PIN pd11_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -37.350 -42.450 -37.050 -20.000 ;
        RECT -41.350 -42.750 -37.050 -42.450 ;
        RECT -57.350 -45.150 -53.300 -45.000 ;
        RECT -41.350 -45.150 -41.050 -42.750 ;
        RECT -57.350 -45.450 -41.050 -45.150 ;
        RECT -57.350 -45.600 -53.300 -45.450 ;
    END
  END pd11_a
  PIN pd11_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -57.350 -40.150 -53.300 -40.000 ;
        RECT -37.850 -40.150 -37.550 -20.000 ;
        RECT -57.350 -40.450 -37.550 -40.150 ;
        RECT -57.350 -40.600 -53.350 -40.450 ;
    END
  END pd11_b
  PIN PD12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.160000 ;
    PORT
      LAYER li1 ;
        RECT 47.280 25.630 48.320 25.800 ;
        RECT 49.150 25.550 49.450 26.000 ;
        RECT 49.250 24.750 49.450 25.550 ;
        RECT 47.280 24.450 48.320 24.620 ;
        RECT 49.200 24.300 49.500 24.750 ;
        RECT 47.230 22.430 48.270 22.600 ;
        RECT 47.230 21.250 48.270 21.420 ;
      LAYER mcon ;
        RECT 47.360 25.630 48.240 25.800 ;
        RECT 49.200 25.650 49.400 25.900 ;
        RECT 47.360 24.450 48.240 24.620 ;
        RECT 49.250 24.400 49.450 24.650 ;
        RECT 47.310 22.430 48.190 22.600 ;
        RECT 47.310 21.250 48.190 21.420 ;
      LAYER met1 ;
        RECT 48.510 27.040 48.770 27.360 ;
        RECT 48.515 25.900 48.765 27.040 ;
        RECT 49.150 25.900 49.450 26.000 ;
        RECT 47.800 25.830 49.450 25.900 ;
        RECT 47.300 25.650 49.450 25.830 ;
        RECT 47.300 25.600 48.300 25.650 ;
        RECT 49.150 25.550 49.450 25.650 ;
        RECT 49.200 24.650 49.500 24.750 ;
        RECT 47.300 24.420 49.500 24.650 ;
        RECT 47.800 24.400 49.500 24.420 ;
        RECT 48.800 24.300 49.500 24.400 ;
        RECT 48.800 24.160 49.360 24.300 ;
        RECT 48.800 22.700 49.120 24.160 ;
        RECT 47.850 22.630 50.150 22.700 ;
        RECT 47.250 22.450 50.150 22.630 ;
        RECT 47.250 22.400 48.250 22.450 ;
        RECT 47.250 21.400 48.250 21.450 ;
        RECT 49.900 21.400 50.150 22.450 ;
        RECT 47.250 21.220 50.150 21.400 ;
        RECT 47.800 21.150 50.150 21.220 ;
      LAYER via ;
        RECT 48.510 27.070 48.770 27.330 ;
      LAYER met2 ;
        RECT 48.000 38.400 48.600 42.450 ;
        RECT 48.170 38.230 48.470 38.400 ;
        RECT 48.170 37.930 48.790 38.230 ;
        RECT 48.490 37.580 48.790 37.930 ;
        RECT 48.455 37.300 48.825 37.580 ;
        RECT 48.490 37.290 48.790 37.300 ;
        RECT 48.445 27.050 48.835 27.350 ;
      LAYER via2 ;
        RECT 48.500 37.300 48.780 37.580 ;
        RECT 48.490 27.050 48.790 27.350 ;
      LAYER met3 ;
        RECT 48.475 37.275 48.805 37.605 ;
        RECT 48.490 27.375 48.790 37.275 ;
        RECT 48.465 27.025 48.815 27.375 ;
    END
  END PD12
  PIN pd12_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -57.350 -35.150 -53.300 -35.000 ;
        RECT -38.450 -35.150 -38.150 -20.000 ;
        RECT -57.350 -35.450 -38.150 -35.150 ;
        RECT -57.350 -35.600 -53.300 -35.450 ;
    END
  END pd12_a
  PIN pd12_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -57.350 -30.150 -53.300 -30.000 ;
        RECT -39.050 -30.150 -38.750 -20.000 ;
        RECT -57.350 -30.450 -38.750 -30.150 ;
        RECT -57.350 -30.600 -53.300 -30.450 ;
    END
  END pd12_b
  PIN Vref_sel_c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.600000 ;
    PORT
      LAYER li1 ;
        RECT 60.800 -18.655 61.150 -18.485 ;
        RECT 68.580 -18.550 68.930 -18.485 ;
        RECT 68.500 -18.655 68.930 -18.550 ;
        RECT 59.700 -19.230 60.180 -19.110 ;
        RECT 60.860 -19.230 61.060 -18.655 ;
        RECT 68.500 -18.750 68.900 -18.655 ;
        RECT 68.500 -19.050 68.800 -18.750 ;
        RECT 59.700 -19.470 61.060 -19.230 ;
        RECT 67.500 -19.350 68.800 -19.050 ;
        RECT 59.700 -19.590 60.180 -19.470 ;
        RECT 60.780 -20.050 60.980 -19.470 ;
        RECT 68.500 -19.550 68.800 -19.350 ;
        RECT 68.500 -19.750 71.200 -19.550 ;
        RECT 68.500 -20.050 68.800 -19.750 ;
        RECT 71.000 -19.950 71.200 -19.750 ;
        RECT 71.000 -20.050 71.900 -19.950 ;
        RECT 60.710 -20.220 61.040 -20.050 ;
        RECT 68.490 -20.220 68.820 -20.050 ;
        RECT 70.965 -20.150 71.900 -20.050 ;
        RECT 70.965 -20.220 71.295 -20.150 ;
        RECT 71.555 -20.220 71.885 -20.150 ;
      LAYER mcon ;
        RECT 59.780 -19.510 60.100 -19.190 ;
      LAYER met1 ;
        RECT 67.500 -15.600 67.800 -15.570 ;
        RECT 59.600 -15.900 67.800 -15.600 ;
        RECT 59.600 -19.110 59.900 -15.900 ;
        RECT 67.500 -15.930 67.800 -15.900 ;
        RECT 59.600 -19.200 60.180 -19.110 ;
        RECT 25.750 -19.500 60.180 -19.200 ;
        RECT 67.440 -19.380 67.860 -19.020 ;
        RECT 25.750 -23.080 26.050 -19.500 ;
        RECT 59.700 -19.590 60.180 -19.500 ;
        RECT 25.750 -67.380 26.050 -37.120 ;
      LAYER via ;
        RECT 67.500 -15.900 67.800 -15.600 ;
        RECT 67.470 -19.380 67.830 -19.020 ;
        RECT 25.750 -23.050 26.050 -22.750 ;
        RECT 25.750 -37.450 26.050 -37.150 ;
        RECT 25.750 -67.350 26.050 -67.050 ;
      LAYER met2 ;
        RECT 67.470 -15.900 67.830 -15.600 ;
        RECT 67.500 -18.950 67.800 -15.900 ;
        RECT 67.400 -19.450 67.900 -18.950 ;
        RECT 25.720 -23.050 26.080 -22.750 ;
        RECT 25.750 -37.150 26.050 -23.050 ;
        RECT 25.720 -37.450 26.080 -37.150 ;
        RECT 25.150 -67.350 26.080 -67.050 ;
        RECT 25.150 -68.350 25.450 -67.350 ;
        RECT 25.000 -72.350 25.600 -68.350 ;
    END
  END Vref_sel_c
  OBS
      LAYER nwell ;
        RECT 37.500 -22.450 40.460 -19.610 ;
        RECT 33.000 -26.650 35.960 -23.810 ;
        RECT 37.500 -26.650 40.460 -23.810 ;
      LAYER li1 ;
        RECT 40.350 25.585 40.650 25.650 ;
        RECT 46.800 25.585 47.100 25.650 ;
        RECT 40.350 25.255 40.660 25.585 ;
        RECT 46.800 25.255 47.110 25.585 ;
        RECT -23.670 25.040 -22.630 25.210 ;
        RECT -17.220 25.040 -16.180 25.210 ;
        RECT -10.770 25.040 -9.730 25.210 ;
        RECT -4.320 25.040 -3.280 25.210 ;
        RECT 2.130 25.040 3.170 25.210 ;
        RECT 8.580 25.040 9.620 25.210 ;
        RECT 15.030 25.040 16.070 25.210 ;
        RECT 21.480 25.040 22.520 25.210 ;
        RECT 27.930 25.040 28.970 25.210 ;
        RECT 34.380 25.040 35.420 25.210 ;
        RECT 40.350 24.995 40.650 25.255 ;
        RECT 40.830 25.040 41.870 25.210 ;
        RECT 46.800 24.995 47.100 25.255 ;
        RECT 47.280 25.040 48.320 25.210 ;
        RECT 40.350 24.665 40.660 24.995 ;
        RECT 46.800 24.665 47.110 24.995 ;
        RECT 40.350 24.650 40.650 24.665 ;
        RECT 46.800 24.650 47.100 24.665 ;
        RECT 40.350 22.385 40.650 22.450 ;
        RECT 46.750 22.385 47.050 22.450 ;
        RECT 40.350 22.055 40.660 22.385 ;
        RECT 46.750 22.055 47.060 22.385 ;
        RECT -23.670 21.840 -22.630 22.010 ;
        RECT -17.270 21.840 -16.230 22.010 ;
        RECT -10.770 21.840 -9.730 22.010 ;
        RECT -4.370 21.840 -3.330 22.010 ;
        RECT 2.130 21.840 3.170 22.010 ;
        RECT 8.530 21.840 9.570 22.010 ;
        RECT 15.030 21.840 16.070 22.010 ;
        RECT 21.430 21.840 22.470 22.010 ;
        RECT 27.930 21.840 28.970 22.010 ;
        RECT 34.330 21.840 35.370 22.010 ;
        RECT 40.350 21.795 40.650 22.055 ;
        RECT 40.830 21.840 41.870 22.010 ;
        RECT 46.750 21.795 47.050 22.055 ;
        RECT 47.230 21.840 48.270 22.010 ;
        RECT 40.350 21.465 40.660 21.795 ;
        RECT 46.750 21.465 47.060 21.795 ;
        RECT 40.350 21.450 40.650 21.465 ;
        RECT 46.750 21.450 47.050 21.465 ;
        RECT -0.650 12.720 -0.480 13.760 ;
        RECT -0.060 12.720 0.110 13.760 ;
        RECT 0.530 12.720 0.700 13.760 ;
        RECT 2.150 13.030 2.320 14.070 ;
        RECT 2.740 13.030 2.910 14.070 ;
        RECT 3.330 13.030 3.500 14.070 ;
        RECT 19.450 11.730 19.620 12.770 ;
        RECT 22.390 11.730 22.560 12.770 ;
        RECT 24.700 11.730 24.870 12.770 ;
        RECT 27.640 11.730 27.810 12.770 ;
        RECT 29.950 11.730 30.120 12.770 ;
        RECT 32.890 11.730 33.060 12.770 ;
        RECT 35.150 11.730 35.320 12.770 ;
        RECT 38.090 11.730 38.260 12.770 ;
        RECT 40.400 11.730 40.570 12.770 ;
        RECT 43.340 11.730 43.510 12.770 ;
        RECT 46.560 11.730 46.730 12.770 ;
        RECT 21.980 11.450 22.330 11.515 ;
        RECT 22.620 11.450 22.970 11.515 ;
        RECT 27.230 11.450 27.580 11.515 ;
        RECT 27.870 11.450 28.220 11.515 ;
        RECT 32.480 11.450 32.830 11.515 ;
        RECT 33.120 11.450 33.470 11.515 ;
        RECT 37.680 11.450 38.030 11.515 ;
        RECT 38.320 11.450 38.670 11.515 ;
        RECT 42.930 11.450 43.280 11.515 ;
        RECT 43.570 11.450 43.920 11.515 ;
        RECT 21.980 11.345 23.000 11.450 ;
        RECT 27.230 11.345 28.250 11.450 ;
        RECT 32.480 11.345 33.500 11.450 ;
        RECT 37.680 11.345 38.700 11.450 ;
        RECT 42.930 11.345 43.950 11.450 ;
        RECT 46.150 11.345 46.500 11.515 ;
        RECT 22.000 11.250 23.000 11.345 ;
        RECT 27.250 11.250 28.250 11.345 ;
        RECT 32.500 11.250 33.500 11.345 ;
        RECT 37.700 11.250 38.700 11.345 ;
        RECT 42.950 11.250 43.950 11.345 ;
        RECT 20.100 10.950 20.500 11.050 ;
        RECT 22.000 10.950 22.200 11.250 ;
        RECT 20.100 10.750 22.200 10.950 ;
        RECT 25.350 10.950 25.750 11.050 ;
        RECT 27.250 10.950 27.450 11.250 ;
        RECT 25.350 10.750 27.450 10.950 ;
        RECT 30.600 10.950 31.000 11.050 ;
        RECT 32.500 10.950 32.700 11.250 ;
        RECT 30.600 10.750 32.700 10.950 ;
        RECT 35.800 10.950 36.200 11.050 ;
        RECT 37.700 10.950 37.900 11.250 ;
        RECT 35.800 10.750 37.900 10.950 ;
        RECT 41.050 10.950 41.450 11.050 ;
        RECT 42.950 10.950 43.150 11.250 ;
        RECT 41.050 10.750 43.150 10.950 ;
        RECT 45.050 10.770 45.530 10.890 ;
        RECT 46.210 10.770 46.410 11.345 ;
        RECT 20.100 10.650 20.500 10.750 ;
        RECT 25.350 10.650 25.750 10.750 ;
        RECT 30.600 10.650 31.000 10.750 ;
        RECT 35.800 10.650 36.200 10.750 ;
        RECT 41.050 10.650 41.450 10.750 ;
        RECT 45.050 10.530 46.410 10.770 ;
        RECT 45.050 10.410 45.530 10.530 ;
        RECT 46.130 9.950 46.330 10.530 ;
        RECT 46.060 9.780 46.390 9.950 ;
        RECT 19.450 8.570 19.620 9.610 ;
        RECT 21.850 8.570 22.020 9.610 ;
        RECT 23.030 8.570 23.200 9.610 ;
        RECT 24.700 8.570 24.870 9.610 ;
        RECT 27.100 8.570 27.270 9.610 ;
        RECT 28.280 8.570 28.450 9.610 ;
        RECT 29.950 8.570 30.120 9.610 ;
        RECT 32.350 8.570 32.520 9.610 ;
        RECT 33.530 8.570 33.700 9.610 ;
        RECT 35.150 8.570 35.320 9.610 ;
        RECT 37.550 8.570 37.720 9.610 ;
        RECT 38.730 8.570 38.900 9.610 ;
        RECT 40.400 8.570 40.570 9.610 ;
        RECT 42.800 8.570 42.970 9.610 ;
        RECT 43.980 8.570 44.150 9.610 ;
        RECT 46.360 8.570 46.530 9.610 ;
        RECT -19.250 7.280 -19.080 8.320 ;
        RECT -16.950 7.280 -16.780 8.320 ;
        RECT -16.310 7.280 -16.140 8.320 ;
        RECT -15.670 7.280 -15.500 8.320 ;
        RECT -14.050 7.280 -13.880 8.320 ;
        RECT -11.750 7.280 -11.580 8.320 ;
        RECT -11.110 7.280 -10.940 8.320 ;
        RECT -10.470 7.280 -10.300 8.320 ;
        RECT -8.850 7.280 -8.680 8.320 ;
        RECT -6.550 7.280 -6.380 8.320 ;
        RECT -5.910 7.280 -5.740 8.320 ;
        RECT -5.270 7.280 -5.100 8.320 ;
        RECT -3.650 7.280 -3.480 8.320 ;
        RECT -1.350 7.280 -1.180 8.320 ;
        RECT -0.710 7.280 -0.540 8.320 ;
        RECT -0.070 7.280 0.100 8.320 ;
        RECT -16.720 7.000 -16.370 7.065 ;
        RECT -16.080 7.000 -15.730 7.065 ;
        RECT -11.520 7.000 -11.170 7.065 ;
        RECT -10.880 7.000 -10.530 7.065 ;
        RECT -6.320 7.000 -5.970 7.065 ;
        RECT -5.680 7.000 -5.330 7.065 ;
        RECT -1.120 7.000 -0.770 7.065 ;
        RECT -0.480 7.000 -0.130 7.065 ;
        RECT -16.720 6.895 -15.700 7.000 ;
        RECT -11.520 6.895 -10.500 7.000 ;
        RECT -6.320 6.895 -5.300 7.000 ;
        RECT -1.120 6.895 -0.100 7.000 ;
        RECT -16.700 6.800 -15.700 6.895 ;
        RECT -11.500 6.800 -10.500 6.895 ;
        RECT -6.300 6.800 -5.300 6.895 ;
        RECT -1.100 6.800 -0.100 6.895 ;
        RECT -18.600 6.500 -18.200 6.600 ;
        RECT -16.700 6.500 -16.500 6.800 ;
        RECT -18.600 6.300 -16.500 6.500 ;
        RECT -13.400 6.500 -13.000 6.600 ;
        RECT -11.500 6.500 -11.300 6.800 ;
        RECT -13.400 6.300 -11.300 6.500 ;
        RECT -8.200 6.500 -7.800 6.600 ;
        RECT -6.300 6.500 -6.100 6.800 ;
        RECT -8.200 6.300 -6.100 6.500 ;
        RECT -3.000 6.500 -2.600 6.600 ;
        RECT -1.100 6.500 -0.900 6.800 ;
        RECT -3.000 6.300 -0.900 6.500 ;
        RECT -18.600 6.200 -18.200 6.300 ;
        RECT -13.400 6.200 -13.000 6.300 ;
        RECT -8.200 6.200 -7.800 6.300 ;
        RECT -3.000 6.200 -2.600 6.300 ;
        RECT -19.250 4.120 -19.080 5.160 ;
        RECT -16.850 4.120 -16.680 5.160 ;
        RECT -16.260 4.120 -16.090 5.160 ;
        RECT -15.670 4.120 -15.500 5.160 ;
        RECT -14.050 4.120 -13.880 5.160 ;
        RECT -11.650 4.120 -11.480 5.160 ;
        RECT -11.060 4.120 -10.890 5.160 ;
        RECT -10.470 4.120 -10.300 5.160 ;
        RECT -8.850 4.120 -8.680 5.160 ;
        RECT -6.450 4.120 -6.280 5.160 ;
        RECT -5.860 4.120 -5.690 5.160 ;
        RECT -5.270 4.120 -5.100 5.160 ;
        RECT -3.650 4.120 -3.480 5.160 ;
        RECT -1.250 4.120 -1.080 5.160 ;
        RECT -0.660 4.120 -0.490 5.160 ;
        RECT -0.070 4.120 0.100 5.160 ;
        RECT -12.800 -1.040 -12.080 -0.880 ;
        RECT -9.680 -1.040 -8.840 -0.920 ;
        RECT 10.700 -1.040 11.420 -0.880 ;
        RECT 13.820 -1.040 14.660 -0.920 ;
        RECT 30.950 -1.040 31.670 -0.880 ;
        RECT 34.070 -1.040 34.910 -0.920 ;
        RECT -19.040 -1.240 -11.840 -1.040 ;
        RECT -9.800 -1.055 -2.640 -1.040 ;
        RECT -9.820 -1.225 -2.640 -1.055 ;
        RECT -9.800 -1.240 -2.640 -1.225 ;
        RECT 4.460 -1.240 11.660 -1.040 ;
        RECT 13.700 -1.055 20.860 -1.040 ;
        RECT 13.680 -1.225 20.860 -1.055 ;
        RECT 13.700 -1.240 20.860 -1.225 ;
        RECT 24.710 -1.240 31.910 -1.040 ;
        RECT 33.950 -1.055 41.110 -1.040 ;
        RECT 33.930 -1.225 41.110 -1.055 ;
        RECT 33.950 -1.240 41.110 -1.225 ;
        RECT -19.250 -3.880 -19.080 -1.440 ;
        RECT -17.760 -3.880 -17.590 -1.440 ;
        RECT -16.270 -3.880 -16.100 -1.440 ;
        RECT -14.780 -3.880 -14.610 -1.440 ;
        RECT -13.290 -3.880 -13.120 -1.440 ;
        RECT -11.800 -3.880 -11.630 -1.440 ;
        RECT -10.050 -3.880 -9.880 -1.440 ;
        RECT -8.560 -3.880 -8.390 -1.440 ;
        RECT -7.070 -3.880 -6.900 -1.440 ;
        RECT -5.580 -3.880 -5.410 -1.440 ;
        RECT -4.090 -3.880 -3.920 -1.440 ;
        RECT -2.600 -3.880 -2.430 -1.440 ;
        RECT 4.250 -3.880 4.420 -1.440 ;
        RECT 5.740 -3.880 5.910 -1.440 ;
        RECT 7.230 -3.880 7.400 -1.440 ;
        RECT 8.720 -3.880 8.890 -1.440 ;
        RECT 10.210 -3.880 10.380 -1.440 ;
        RECT 11.700 -3.880 11.870 -1.440 ;
        RECT 13.450 -3.880 13.620 -1.440 ;
        RECT 14.940 -3.880 15.110 -1.440 ;
        RECT 16.430 -3.880 16.600 -1.440 ;
        RECT 17.920 -3.880 18.090 -1.440 ;
        RECT 19.410 -3.880 19.580 -1.440 ;
        RECT 20.900 -3.880 21.070 -1.440 ;
        RECT 24.500 -3.880 24.670 -1.440 ;
        RECT 25.990 -3.880 26.160 -1.440 ;
        RECT 27.480 -3.880 27.650 -1.440 ;
        RECT 28.970 -3.880 29.140 -1.440 ;
        RECT 30.460 -3.880 30.630 -1.440 ;
        RECT 31.950 -3.880 32.120 -1.440 ;
        RECT 33.700 -3.880 33.870 -1.440 ;
        RECT 35.190 -3.880 35.360 -1.440 ;
        RECT 36.680 -3.880 36.850 -1.440 ;
        RECT 38.170 -3.880 38.340 -1.440 ;
        RECT 39.660 -3.880 39.830 -1.440 ;
        RECT 41.150 -3.880 41.320 -1.440 ;
        RECT -19.250 -7.320 -19.080 -5.280 ;
        RECT -16.250 -6.320 -16.080 -5.280 ;
        RECT -12.850 -6.370 -12.680 -5.330 ;
        RECT -9.060 -6.370 -8.890 -5.330 ;
        RECT -16.020 -6.705 -15.020 -6.535 ;
        RECT -12.620 -6.710 -12.120 -6.540 ;
        RECT -9.620 -6.710 -9.120 -6.540 ;
        RECT -5.260 -7.020 -5.090 -5.270 ;
        RECT -2.680 -7.020 -2.510 -5.270 ;
        RECT -6.700 -7.400 -2.700 -7.200 ;
        RECT 4.250 -7.320 4.420 -5.280 ;
        RECT 7.250 -6.320 7.420 -5.280 ;
        RECT 10.650 -6.370 10.820 -5.330 ;
        RECT 14.440 -6.370 14.610 -5.330 ;
        RECT 7.480 -6.705 8.480 -6.535 ;
        RECT 10.880 -6.710 11.380 -6.540 ;
        RECT 13.880 -6.710 14.380 -6.540 ;
        RECT 18.240 -7.020 18.410 -5.270 ;
        RECT 20.820 -7.020 20.990 -5.270 ;
        RECT 16.800 -7.400 20.800 -7.200 ;
        RECT 24.500 -7.320 24.670 -5.280 ;
        RECT 27.500 -6.320 27.670 -5.280 ;
        RECT 30.900 -6.370 31.070 -5.330 ;
        RECT 34.690 -6.370 34.860 -5.330 ;
        RECT 27.730 -6.705 28.730 -6.535 ;
        RECT 31.130 -6.710 31.630 -6.540 ;
        RECT 34.130 -6.710 34.630 -6.540 ;
        RECT 38.490 -7.020 38.660 -5.270 ;
        RECT 41.070 -7.020 41.240 -5.270 ;
        RECT 37.050 -7.400 41.050 -7.200 ;
        RECT -6.700 -7.405 -5.320 -7.400 ;
        RECT -5.030 -7.405 -4.030 -7.400 ;
        RECT -3.740 -7.405 -2.740 -7.400 ;
        RECT 16.800 -7.405 18.180 -7.400 ;
        RECT 18.470 -7.405 19.470 -7.400 ;
        RECT 19.760 -7.405 20.760 -7.400 ;
        RECT 37.050 -7.405 38.430 -7.400 ;
        RECT 38.720 -7.405 39.720 -7.400 ;
        RECT 40.010 -7.405 41.010 -7.400 ;
        RECT -6.700 -7.500 -5.800 -7.405 ;
        RECT 16.800 -7.500 17.700 -7.405 ;
        RECT 37.050 -7.500 37.950 -7.405 ;
        RECT -19.020 -7.705 -18.020 -7.535 ;
        RECT 0.750 -8.570 0.920 -7.530 ;
        RECT 1.340 -8.570 1.510 -7.530 ;
        RECT 1.930 -8.570 2.100 -7.530 ;
        RECT 4.480 -7.705 5.480 -7.535 ;
        RECT 24.730 -7.705 25.730 -7.535 ;
        RECT -16.100 -9.000 -3.400 -8.800 ;
        RECT 7.400 -9.000 20.100 -8.800 ;
        RECT 27.650 -9.000 40.350 -8.800 ;
        RECT -16.020 -9.020 -15.020 -9.000 ;
        RECT -14.730 -9.020 -13.730 -9.000 ;
        RECT -13.440 -9.020 -12.440 -9.000 ;
        RECT -12.150 -9.020 -11.150 -9.000 ;
        RECT -10.860 -9.020 -9.860 -9.000 ;
        RECT -9.570 -9.020 -8.570 -9.000 ;
        RECT -8.280 -9.020 -7.280 -9.000 ;
        RECT -6.990 -9.020 -5.990 -9.000 ;
        RECT -5.700 -9.020 -4.700 -9.000 ;
        RECT -4.410 -9.020 -3.410 -9.000 ;
        RECT 7.480 -9.020 8.480 -9.000 ;
        RECT 8.770 -9.020 9.770 -9.000 ;
        RECT 10.060 -9.020 11.060 -9.000 ;
        RECT 11.350 -9.020 12.350 -9.000 ;
        RECT 12.640 -9.020 13.640 -9.000 ;
        RECT 13.930 -9.020 14.930 -9.000 ;
        RECT 15.220 -9.020 16.220 -9.000 ;
        RECT 16.510 -9.020 17.510 -9.000 ;
        RECT 17.800 -9.020 18.800 -9.000 ;
        RECT 19.090 -9.020 20.090 -9.000 ;
        RECT 27.730 -9.020 28.730 -9.000 ;
        RECT 29.020 -9.020 30.020 -9.000 ;
        RECT 30.310 -9.020 31.310 -9.000 ;
        RECT 31.600 -9.020 32.600 -9.000 ;
        RECT 32.890 -9.020 33.890 -9.000 ;
        RECT 34.180 -9.020 35.180 -9.000 ;
        RECT 35.470 -9.020 36.470 -9.000 ;
        RECT 36.760 -9.020 37.760 -9.000 ;
        RECT 38.050 -9.020 39.050 -9.000 ;
        RECT 39.340 -9.020 40.340 -9.000 ;
        RECT -8.100 -9.150 -7.500 -9.020 ;
        RECT 15.400 -9.150 16.000 -9.020 ;
        RECT 35.650 -9.150 36.250 -9.020 ;
        RECT -14.960 -11.730 -14.790 -9.190 ;
        RECT -12.380 -11.730 -12.210 -9.190 ;
        RECT -9.800 -11.730 -9.630 -9.190 ;
        RECT -7.220 -11.730 -7.050 -9.190 ;
        RECT -4.640 -11.730 -4.470 -9.190 ;
        RECT 8.540 -11.730 8.710 -9.190 ;
        RECT 11.120 -11.730 11.290 -9.190 ;
        RECT 13.700 -11.730 13.870 -9.190 ;
        RECT 16.280 -11.730 16.450 -9.190 ;
        RECT 18.860 -11.730 19.030 -9.190 ;
        RECT 28.790 -11.730 28.960 -9.190 ;
        RECT 31.370 -11.730 31.540 -9.190 ;
        RECT 33.950 -11.730 34.120 -9.190 ;
        RECT 36.530 -11.730 36.700 -9.190 ;
        RECT 39.110 -11.730 39.280 -9.190 ;
        RECT 61.210 -18.270 61.380 -17.230 ;
        RECT 63.100 -18.270 63.270 -17.230 ;
        RECT 65.400 -18.270 65.570 -17.230 ;
        RECT 66.040 -18.270 66.210 -17.230 ;
        RECT 66.680 -18.270 66.850 -17.230 ;
        RECT 68.350 -18.270 68.520 -17.230 ;
        RECT 70.650 -18.270 70.820 -17.230 ;
        RECT 71.290 -18.270 71.460 -17.230 ;
        RECT 71.930 -18.270 72.100 -17.230 ;
        RECT 63.330 -18.550 63.680 -18.485 ;
        RECT 63.250 -18.655 63.680 -18.550 ;
        RECT 65.630 -18.550 65.980 -18.485 ;
        RECT 66.270 -18.550 66.620 -18.485 ;
        RECT 70.880 -18.550 71.230 -18.485 ;
        RECT 71.520 -18.550 71.870 -18.485 ;
        RECT 65.630 -18.655 66.650 -18.550 ;
        RECT 70.880 -18.655 71.900 -18.550 ;
        RECT 63.250 -18.750 63.650 -18.655 ;
        RECT 65.650 -18.750 66.650 -18.655 ;
        RECT 70.900 -18.750 71.900 -18.655 ;
        RECT 62.000 -19.050 62.400 -19.000 ;
        RECT 63.250 -19.050 63.550 -18.750 ;
        RECT 62.000 -19.350 63.550 -19.050 ;
        RECT 63.750 -19.050 64.150 -18.950 ;
        RECT 65.650 -19.050 65.850 -18.750 ;
        RECT 63.750 -19.250 65.850 -19.050 ;
        RECT 69.000 -19.050 69.400 -18.950 ;
        RECT 70.900 -19.050 71.100 -18.750 ;
        RECT 69.000 -19.250 71.100 -19.050 ;
        RECT 63.750 -19.350 64.150 -19.250 ;
        RECT 69.000 -19.350 69.400 -19.250 ;
        RECT 62.000 -19.600 62.400 -19.350 ;
        RECT 63.250 -19.550 63.550 -19.350 ;
        RECT 37.600 -20.050 40.300 -19.650 ;
        RECT 63.250 -19.750 65.950 -19.550 ;
        RECT 63.250 -20.050 63.550 -19.750 ;
        RECT 65.750 -19.950 65.950 -19.750 ;
        RECT 65.750 -20.050 66.650 -19.950 ;
        RECT 33.700 -20.305 34.800 -20.250 ;
        RECT 33.700 -20.475 34.980 -20.305 ;
        RECT 17.140 -23.170 17.310 -22.130 ;
        RECT 33.180 -24.550 33.350 -24.395 ;
        RECT 33.700 -24.550 34.000 -20.475 ;
        RECT 37.600 -21.550 37.900 -20.050 ;
        RECT 39.540 -20.850 39.710 -20.690 ;
        RECT 39.900 -20.850 40.300 -20.050 ;
        RECT 63.240 -20.220 63.570 -20.050 ;
        RECT 65.715 -20.150 66.650 -20.050 ;
        RECT 65.715 -20.220 66.045 -20.150 ;
        RECT 66.305 -20.220 66.635 -20.150 ;
        RECT 37.680 -21.865 37.850 -21.550 ;
        RECT 39.500 -21.650 40.300 -20.850 ;
        RECT 61.010 -21.430 61.180 -20.390 ;
        RECT 63.100 -21.430 63.270 -20.390 ;
        RECT 65.500 -21.430 65.670 -20.390 ;
        RECT 66.090 -21.430 66.260 -20.390 ;
        RECT 66.680 -21.430 66.850 -20.390 ;
        RECT 68.350 -21.430 68.520 -20.390 ;
        RECT 70.750 -21.430 70.920 -20.390 ;
        RECT 71.340 -21.430 71.510 -20.390 ;
        RECT 71.930 -21.430 72.100 -20.390 ;
        RECT 39.500 -22.950 39.800 -21.650 ;
        RECT 40.110 -21.865 40.280 -21.650 ;
        RECT 39.500 -23.200 50.250 -22.950 ;
        RECT 39.500 -23.450 40.100 -23.200 ;
        RECT 33.180 -25.550 34.000 -24.550 ;
        RECT 35.000 -24.050 37.900 -23.750 ;
        RECT 33.180 -26.065 33.500 -25.550 ;
        RECT 33.750 -25.570 33.920 -25.550 ;
        RECT 35.000 -25.750 35.300 -24.050 ;
        RECT 36.590 -24.150 37.100 -24.050 ;
        RECT 35.610 -24.450 35.780 -24.395 ;
        RECT 34.000 -25.785 35.300 -25.750 ;
        RECT 33.980 -25.950 35.300 -25.785 ;
        RECT 33.980 -25.955 34.980 -25.950 ;
        RECT 33.200 -26.150 33.500 -26.065 ;
        RECT 35.500 -26.150 35.800 -24.450 ;
        RECT 36.600 -24.650 37.100 -24.150 ;
        RECT 37.600 -24.550 37.900 -24.050 ;
        RECT 38.250 -24.550 38.420 -24.530 ;
        RECT 36.600 -24.700 37.050 -24.650 ;
        RECT 33.200 -26.550 35.800 -26.150 ;
        RECT 37.600 -25.450 38.420 -24.550 ;
        RECT 37.600 -26.250 37.900 -25.450 ;
        RECT 38.250 -25.570 38.420 -25.450 ;
        RECT 39.500 -25.750 39.800 -23.450 ;
        RECT 49.800 -23.600 50.300 -23.200 ;
        RECT 40.110 -24.450 40.280 -24.395 ;
        RECT 38.500 -25.785 39.800 -25.750 ;
        RECT 38.480 -25.950 39.800 -25.785 ;
        RECT 38.480 -25.955 39.480 -25.950 ;
        RECT 40.000 -26.250 40.300 -24.450 ;
        RECT 49.640 -24.540 50.480 -24.420 ;
        RECT 52.880 -24.540 53.600 -24.380 ;
        RECT 69.490 -24.540 70.330 -24.420 ;
        RECT 72.730 -24.540 73.450 -24.380 ;
        RECT 43.440 -24.555 50.600 -24.540 ;
        RECT 43.440 -24.725 50.620 -24.555 ;
        RECT 43.440 -24.740 50.600 -24.725 ;
        RECT 52.640 -24.740 59.840 -24.540 ;
        RECT 63.290 -24.555 70.450 -24.540 ;
        RECT 63.290 -24.725 70.470 -24.555 ;
        RECT 63.290 -24.740 70.450 -24.725 ;
        RECT 72.490 -24.740 79.690 -24.540 ;
        RECT 37.600 -26.650 40.300 -26.250 ;
        RECT 40.000 -26.750 40.300 -26.650 ;
        RECT 17.140 -27.880 17.310 -26.840 ;
        RECT 20.145 -27.875 20.315 -26.835 ;
        RECT 43.230 -27.380 43.400 -24.940 ;
        RECT 44.720 -27.380 44.890 -24.940 ;
        RECT 46.210 -27.380 46.380 -24.940 ;
        RECT 47.700 -27.380 47.870 -24.940 ;
        RECT 49.190 -27.380 49.360 -24.940 ;
        RECT 50.680 -27.380 50.850 -24.940 ;
        RECT 52.430 -27.380 52.600 -24.940 ;
        RECT 53.920 -27.380 54.090 -24.940 ;
        RECT 55.410 -27.380 55.580 -24.940 ;
        RECT 56.900 -27.380 57.070 -24.940 ;
        RECT 58.390 -27.380 58.560 -24.940 ;
        RECT 59.880 -27.380 60.050 -24.940 ;
        RECT 63.080 -27.380 63.250 -24.940 ;
        RECT 64.570 -27.380 64.740 -24.940 ;
        RECT 66.060 -27.380 66.230 -24.940 ;
        RECT 67.550 -27.380 67.720 -24.940 ;
        RECT 69.040 -27.380 69.210 -24.940 ;
        RECT 70.530 -27.380 70.700 -24.940 ;
        RECT 72.280 -27.380 72.450 -24.940 ;
        RECT 73.770 -27.380 73.940 -24.940 ;
        RECT 75.260 -27.380 75.430 -24.940 ;
        RECT 76.750 -27.380 76.920 -24.940 ;
        RECT 78.240 -27.380 78.410 -24.940 ;
        RECT 79.730 -27.380 79.900 -24.940 ;
        RECT 17.140 -30.570 17.310 -29.530 ;
        RECT 22.950 -30.920 23.120 -28.680 ;
        RECT 25.530 -30.920 25.700 -28.680 ;
        RECT 28.110 -30.920 28.280 -28.680 ;
        RECT 30.690 -30.920 30.860 -28.680 ;
        RECT 33.270 -30.920 33.440 -28.680 ;
        RECT 35.850 -30.920 36.020 -28.680 ;
        RECT 40.040 -30.920 40.210 -29.880 ;
        RECT 43.310 -30.520 43.480 -28.770 ;
        RECT 45.890 -30.520 46.060 -28.770 ;
        RECT 49.690 -29.870 49.860 -28.830 ;
        RECT 53.480 -29.870 53.650 -28.830 ;
        RECT 56.880 -29.820 57.050 -28.780 ;
        RECT 49.920 -30.210 50.420 -30.040 ;
        RECT 52.920 -30.210 53.420 -30.040 ;
        RECT 55.820 -30.205 56.820 -30.035 ;
        RECT 43.500 -30.900 47.500 -30.700 ;
        RECT 59.880 -30.820 60.050 -28.780 ;
        RECT 63.160 -30.520 63.330 -28.770 ;
        RECT 65.740 -30.520 65.910 -28.770 ;
        RECT 69.540 -29.870 69.710 -28.830 ;
        RECT 73.330 -29.870 73.500 -28.830 ;
        RECT 76.730 -29.820 76.900 -28.780 ;
        RECT 69.770 -30.210 70.270 -30.040 ;
        RECT 72.770 -30.210 73.270 -30.040 ;
        RECT 75.670 -30.205 76.670 -30.035 ;
        RECT 63.350 -30.900 67.350 -30.700 ;
        RECT 79.730 -30.820 79.900 -28.780 ;
        RECT 43.540 -30.905 44.540 -30.900 ;
        RECT 44.830 -30.905 45.830 -30.900 ;
        RECT 46.120 -30.905 47.500 -30.900 ;
        RECT 63.390 -30.905 64.390 -30.900 ;
        RECT 64.680 -30.905 65.680 -30.900 ;
        RECT 65.970 -30.905 67.350 -30.900 ;
        RECT 46.600 -31.000 47.500 -30.905 ;
        RECT 66.450 -31.000 67.350 -30.905 ;
        RECT 23.180 -31.305 24.180 -31.135 ;
        RECT 24.470 -31.305 25.470 -31.135 ;
        RECT 25.760 -31.305 26.760 -31.135 ;
        RECT 27.050 -31.305 28.050 -31.135 ;
        RECT 28.340 -31.305 29.340 -31.135 ;
        RECT 29.630 -31.305 30.630 -31.135 ;
        RECT 30.920 -31.305 31.920 -31.135 ;
        RECT 32.210 -31.305 33.210 -31.135 ;
        RECT 33.500 -31.305 34.500 -31.135 ;
        RECT 34.790 -31.305 35.790 -31.135 ;
        RECT 36.080 -31.305 37.080 -31.135 ;
        RECT 38.980 -31.305 39.980 -31.135 ;
        RECT 58.820 -31.205 59.820 -31.035 ;
        RECT 78.670 -31.205 79.670 -31.035 ;
        RECT 44.200 -32.500 56.900 -32.300 ;
        RECT 64.050 -32.500 76.750 -32.300 ;
        RECT 44.210 -32.520 45.210 -32.500 ;
        RECT 45.500 -32.520 46.500 -32.500 ;
        RECT 46.790 -32.520 47.790 -32.500 ;
        RECT 48.080 -32.520 49.080 -32.500 ;
        RECT 49.370 -32.520 50.370 -32.500 ;
        RECT 50.660 -32.520 51.660 -32.500 ;
        RECT 51.950 -32.520 52.950 -32.500 ;
        RECT 53.240 -32.520 54.240 -32.500 ;
        RECT 54.530 -32.520 55.530 -32.500 ;
        RECT 55.820 -32.520 56.820 -32.500 ;
        RECT 64.060 -32.520 65.060 -32.500 ;
        RECT 65.350 -32.520 66.350 -32.500 ;
        RECT 66.640 -32.520 67.640 -32.500 ;
        RECT 67.930 -32.520 68.930 -32.500 ;
        RECT 69.220 -32.520 70.220 -32.500 ;
        RECT 70.510 -32.520 71.510 -32.500 ;
        RECT 71.800 -32.520 72.800 -32.500 ;
        RECT 73.090 -32.520 74.090 -32.500 ;
        RECT 74.380 -32.520 75.380 -32.500 ;
        RECT 75.670 -32.520 76.670 -32.500 ;
        RECT 48.300 -32.650 48.900 -32.520 ;
        RECT 68.150 -32.650 68.750 -32.520 ;
        RECT 23.180 -32.870 24.180 -32.700 ;
        RECT 24.470 -32.870 25.470 -32.700 ;
        RECT 25.760 -32.870 26.760 -32.700 ;
        RECT 27.050 -32.870 28.050 -32.700 ;
        RECT 28.340 -32.870 29.340 -32.700 ;
        RECT 29.630 -32.870 30.630 -32.700 ;
        RECT 30.920 -32.870 31.920 -32.700 ;
        RECT 32.210 -32.870 33.210 -32.700 ;
        RECT 33.500 -32.870 34.500 -32.700 ;
        RECT 34.790 -32.870 35.790 -32.700 ;
        RECT 36.080 -32.870 37.080 -32.700 ;
        RECT 17.140 -35.280 17.310 -34.240 ;
        RECT 20.145 -35.275 20.315 -34.235 ;
        RECT 24.240 -35.280 24.410 -33.040 ;
        RECT 26.820 -35.280 26.990 -33.040 ;
        RECT 29.400 -35.280 29.570 -33.040 ;
        RECT 31.980 -35.280 32.150 -33.040 ;
        RECT 34.560 -35.280 34.730 -33.040 ;
        RECT 37.140 -35.280 37.310 -33.040 ;
        RECT 38.980 -34.070 39.980 -33.900 ;
        RECT 40.040 -35.280 40.210 -34.240 ;
        RECT 45.270 -35.230 45.440 -32.690 ;
        RECT 47.850 -35.230 48.020 -32.690 ;
        RECT 50.430 -35.230 50.600 -32.690 ;
        RECT 53.010 -35.230 53.180 -32.690 ;
        RECT 55.590 -35.230 55.760 -32.690 ;
        RECT 65.120 -35.230 65.290 -32.690 ;
        RECT 67.700 -35.230 67.870 -32.690 ;
        RECT 70.280 -35.230 70.450 -32.690 ;
        RECT 72.860 -35.230 73.030 -32.690 ;
        RECT 75.440 -35.230 75.610 -32.690 ;
        RECT 43.950 -37.670 44.120 -36.630 ;
        RECT 44.540 -37.670 44.710 -36.630 ;
        RECT 45.130 -37.670 45.300 -36.630 ;
        RECT 46.800 -37.670 46.970 -36.630 ;
        RECT 47.390 -37.670 47.560 -36.630 ;
        RECT 47.980 -37.670 48.150 -36.630 ;
      LAYER mcon ;
        RECT -23.590 25.040 -22.710 25.210 ;
        RECT -17.140 25.040 -16.260 25.210 ;
        RECT -10.690 25.040 -9.810 25.210 ;
        RECT -4.240 25.040 -3.360 25.210 ;
        RECT 2.210 25.040 3.090 25.210 ;
        RECT 8.660 25.040 9.540 25.210 ;
        RECT 15.110 25.040 15.990 25.210 ;
        RECT 21.560 25.040 22.440 25.210 ;
        RECT 28.010 25.040 28.890 25.210 ;
        RECT 34.460 25.040 35.340 25.210 ;
        RECT 40.400 24.800 40.600 25.500 ;
        RECT 40.910 25.040 41.790 25.210 ;
        RECT 46.850 24.800 47.050 25.500 ;
        RECT 47.360 25.040 48.240 25.210 ;
        RECT -23.590 21.840 -22.710 22.010 ;
        RECT -17.190 21.840 -16.310 22.010 ;
        RECT -10.690 21.840 -9.810 22.010 ;
        RECT -4.290 21.840 -3.410 22.010 ;
        RECT 2.210 21.840 3.090 22.010 ;
        RECT 8.610 21.840 9.490 22.010 ;
        RECT 15.110 21.840 15.990 22.010 ;
        RECT 21.510 21.840 22.390 22.010 ;
        RECT 28.010 21.840 28.890 22.010 ;
        RECT 34.410 21.840 35.290 22.010 ;
        RECT 40.400 21.600 40.600 22.300 ;
        RECT 40.910 21.840 41.790 22.010 ;
        RECT 46.800 21.600 47.000 22.300 ;
        RECT 47.310 21.840 48.190 22.010 ;
        RECT -0.650 12.800 -0.480 13.680 ;
        RECT -0.060 12.800 0.110 13.680 ;
        RECT 0.530 12.800 0.700 13.680 ;
        RECT 2.150 13.110 2.320 13.990 ;
        RECT 2.740 13.110 2.910 13.990 ;
        RECT 3.330 13.110 3.500 13.990 ;
        RECT 19.450 11.810 19.620 12.690 ;
        RECT 22.390 11.810 22.560 12.690 ;
        RECT 24.700 11.810 24.870 12.690 ;
        RECT 27.640 11.810 27.810 12.690 ;
        RECT 29.950 11.810 30.120 12.690 ;
        RECT 32.890 11.810 33.060 12.690 ;
        RECT 35.150 11.810 35.320 12.690 ;
        RECT 38.090 11.810 38.260 12.690 ;
        RECT 40.400 11.810 40.570 12.690 ;
        RECT 43.340 11.810 43.510 12.690 ;
        RECT 46.560 11.810 46.730 12.690 ;
        RECT 20.200 10.750 20.400 10.950 ;
        RECT 25.450 10.750 25.650 10.950 ;
        RECT 30.700 10.750 30.900 10.950 ;
        RECT 35.900 10.750 36.100 10.950 ;
        RECT 41.150 10.750 41.350 10.950 ;
        RECT 45.130 10.490 45.450 10.810 ;
        RECT 19.450 8.650 19.620 9.530 ;
        RECT 21.850 8.650 22.020 9.530 ;
        RECT 23.030 8.650 23.200 9.530 ;
        RECT 24.700 8.650 24.870 9.530 ;
        RECT 27.100 8.650 27.270 9.530 ;
        RECT 28.280 8.650 28.450 9.530 ;
        RECT 29.950 8.650 30.120 9.530 ;
        RECT 32.350 8.650 32.520 9.530 ;
        RECT 33.530 8.650 33.700 9.530 ;
        RECT 35.150 8.650 35.320 9.530 ;
        RECT 37.550 8.650 37.720 9.530 ;
        RECT 38.730 8.650 38.900 9.530 ;
        RECT 40.400 8.650 40.570 9.530 ;
        RECT 42.800 8.650 42.970 9.530 ;
        RECT 43.980 8.650 44.150 9.530 ;
        RECT 46.360 8.650 46.530 9.530 ;
        RECT -19.250 7.360 -19.080 8.240 ;
        RECT -16.950 7.360 -16.780 8.240 ;
        RECT -16.310 7.360 -16.140 8.240 ;
        RECT -15.670 7.360 -15.500 8.240 ;
        RECT -14.050 7.360 -13.880 8.240 ;
        RECT -11.750 7.360 -11.580 8.240 ;
        RECT -11.110 7.360 -10.940 8.240 ;
        RECT -10.470 7.360 -10.300 8.240 ;
        RECT -8.850 7.360 -8.680 8.240 ;
        RECT -6.550 7.360 -6.380 8.240 ;
        RECT -5.910 7.360 -5.740 8.240 ;
        RECT -5.270 7.360 -5.100 8.240 ;
        RECT -3.650 7.360 -3.480 8.240 ;
        RECT -1.350 7.360 -1.180 8.240 ;
        RECT -0.710 7.360 -0.540 8.240 ;
        RECT -0.070 7.360 0.100 8.240 ;
        RECT -18.500 6.300 -18.300 6.500 ;
        RECT -13.300 6.300 -13.100 6.500 ;
        RECT -8.100 6.300 -7.900 6.500 ;
        RECT -2.900 6.300 -2.700 6.500 ;
        RECT -19.250 4.200 -19.080 5.080 ;
        RECT -16.850 4.200 -16.680 5.080 ;
        RECT -16.260 4.200 -16.090 5.080 ;
        RECT -15.670 4.200 -15.500 5.080 ;
        RECT -14.050 4.200 -13.880 5.080 ;
        RECT -11.650 4.200 -11.480 5.080 ;
        RECT -11.060 4.200 -10.890 5.080 ;
        RECT -10.470 4.200 -10.300 5.080 ;
        RECT -8.850 4.200 -8.680 5.080 ;
        RECT -6.450 4.200 -6.280 5.080 ;
        RECT -5.860 4.200 -5.690 5.080 ;
        RECT -5.270 4.200 -5.100 5.080 ;
        RECT -3.650 4.200 -3.480 5.080 ;
        RECT -1.250 4.200 -1.080 5.080 ;
        RECT -0.660 4.200 -0.490 5.080 ;
        RECT -0.070 4.200 0.100 5.080 ;
        RECT -12.720 -1.200 -12.160 -0.960 ;
        RECT -9.600 -1.200 -8.920 -1.000 ;
        RECT 10.780 -1.200 11.340 -0.960 ;
        RECT 13.900 -1.200 14.580 -1.000 ;
        RECT 31.030 -1.200 31.590 -0.960 ;
        RECT 34.150 -1.200 34.830 -1.000 ;
        RECT -19.250 -3.800 -19.080 -1.520 ;
        RECT -17.760 -3.800 -17.590 -1.520 ;
        RECT -16.270 -3.800 -16.100 -1.520 ;
        RECT -14.780 -3.800 -14.610 -1.520 ;
        RECT -13.290 -3.800 -13.120 -1.520 ;
        RECT -11.800 -3.800 -11.630 -1.520 ;
        RECT -10.050 -3.800 -9.880 -1.520 ;
        RECT -8.560 -3.800 -8.390 -1.520 ;
        RECT -7.070 -3.800 -6.900 -1.520 ;
        RECT -5.580 -3.800 -5.410 -1.520 ;
        RECT -4.090 -3.800 -3.920 -1.520 ;
        RECT -2.600 -3.800 -2.430 -1.520 ;
        RECT 4.250 -3.800 4.420 -1.520 ;
        RECT 5.740 -3.800 5.910 -1.520 ;
        RECT 7.230 -3.800 7.400 -1.520 ;
        RECT 8.720 -3.800 8.890 -1.520 ;
        RECT 10.210 -3.800 10.380 -1.520 ;
        RECT 11.700 -3.800 11.870 -1.520 ;
        RECT 13.450 -3.800 13.620 -1.520 ;
        RECT 14.940 -3.800 15.110 -1.520 ;
        RECT 16.430 -3.800 16.600 -1.520 ;
        RECT 17.920 -3.800 18.090 -1.520 ;
        RECT 19.410 -3.800 19.580 -1.520 ;
        RECT 20.900 -3.800 21.070 -1.520 ;
        RECT 24.500 -3.800 24.670 -1.520 ;
        RECT 25.990 -3.800 26.160 -1.520 ;
        RECT 27.480 -3.800 27.650 -1.520 ;
        RECT 28.970 -3.800 29.140 -1.520 ;
        RECT 30.460 -3.800 30.630 -1.520 ;
        RECT 31.950 -3.800 32.120 -1.520 ;
        RECT 33.700 -3.800 33.870 -1.520 ;
        RECT 35.190 -3.800 35.360 -1.520 ;
        RECT 36.680 -3.800 36.850 -1.520 ;
        RECT 38.170 -3.800 38.340 -1.520 ;
        RECT 39.660 -3.800 39.830 -1.520 ;
        RECT 41.150 -3.800 41.320 -1.520 ;
        RECT -19.250 -7.240 -19.080 -5.360 ;
        RECT -16.250 -6.240 -16.080 -5.360 ;
        RECT -12.850 -6.290 -12.680 -5.410 ;
        RECT -9.060 -6.290 -8.890 -5.410 ;
        RECT -15.940 -6.705 -15.100 -6.535 ;
        RECT -12.540 -6.710 -12.200 -6.540 ;
        RECT -9.540 -6.710 -9.200 -6.540 ;
        RECT -5.260 -6.940 -5.090 -5.350 ;
        RECT -2.680 -6.940 -2.510 -5.350 ;
        RECT -6.600 -7.450 -5.950 -7.250 ;
        RECT 4.250 -7.240 4.420 -5.360 ;
        RECT 7.250 -6.240 7.420 -5.360 ;
        RECT 10.650 -6.290 10.820 -5.410 ;
        RECT 14.440 -6.290 14.610 -5.410 ;
        RECT 7.560 -6.705 8.400 -6.535 ;
        RECT 10.960 -6.710 11.300 -6.540 ;
        RECT 13.960 -6.710 14.300 -6.540 ;
        RECT 18.240 -6.940 18.410 -5.350 ;
        RECT 20.820 -6.940 20.990 -5.350 ;
        RECT 16.900 -7.450 17.550 -7.250 ;
        RECT 24.500 -7.240 24.670 -5.360 ;
        RECT 27.500 -6.240 27.670 -5.360 ;
        RECT 30.900 -6.290 31.070 -5.410 ;
        RECT 34.690 -6.290 34.860 -5.410 ;
        RECT 27.810 -6.705 28.650 -6.535 ;
        RECT 31.210 -6.710 31.550 -6.540 ;
        RECT 34.210 -6.710 34.550 -6.540 ;
        RECT 38.490 -6.940 38.660 -5.350 ;
        RECT 41.070 -6.940 41.240 -5.350 ;
        RECT 37.150 -7.450 37.800 -7.250 ;
        RECT -18.940 -7.705 -18.100 -7.535 ;
        RECT 0.750 -8.490 0.920 -7.610 ;
        RECT 1.340 -8.490 1.510 -7.610 ;
        RECT 1.930 -8.490 2.100 -7.610 ;
        RECT 4.560 -7.705 5.400 -7.535 ;
        RECT 24.810 -7.705 25.650 -7.535 ;
        RECT -8.000 -9.100 -7.600 -8.900 ;
        RECT 15.500 -9.100 15.900 -8.900 ;
        RECT 35.750 -9.100 36.150 -8.900 ;
        RECT -14.960 -11.650 -14.790 -9.270 ;
        RECT -12.380 -11.650 -12.210 -9.270 ;
        RECT -9.800 -11.650 -9.630 -9.270 ;
        RECT -7.220 -11.650 -7.050 -9.270 ;
        RECT -4.640 -11.650 -4.470 -9.270 ;
        RECT 8.540 -11.650 8.710 -9.270 ;
        RECT 11.120 -11.650 11.290 -9.270 ;
        RECT 13.700 -11.650 13.870 -9.270 ;
        RECT 16.280 -11.650 16.450 -9.270 ;
        RECT 18.860 -11.650 19.030 -9.270 ;
        RECT 28.790 -11.650 28.960 -9.270 ;
        RECT 31.370 -11.650 31.540 -9.270 ;
        RECT 33.950 -11.650 34.120 -9.270 ;
        RECT 36.530 -11.650 36.700 -9.270 ;
        RECT 39.110 -11.650 39.280 -9.270 ;
        RECT 61.210 -18.190 61.380 -17.310 ;
        RECT 63.100 -18.190 63.270 -17.310 ;
        RECT 65.400 -18.190 65.570 -17.310 ;
        RECT 66.040 -18.190 66.210 -17.310 ;
        RECT 66.680 -18.190 66.850 -17.310 ;
        RECT 68.350 -18.190 68.520 -17.310 ;
        RECT 70.650 -18.190 70.820 -17.310 ;
        RECT 71.290 -18.190 71.460 -17.310 ;
        RECT 71.930 -18.190 72.100 -17.310 ;
        RECT 62.100 -19.500 62.300 -19.100 ;
        RECT 63.850 -19.250 64.050 -19.050 ;
        RECT 69.100 -19.250 69.300 -19.050 ;
        RECT 33.750 -21.650 33.920 -20.770 ;
        RECT 17.140 -23.090 17.310 -22.210 ;
        RECT 39.540 -21.650 39.710 -20.770 ;
        RECT 61.010 -21.350 61.180 -20.470 ;
        RECT 63.100 -21.350 63.270 -20.470 ;
        RECT 65.500 -21.350 65.670 -20.470 ;
        RECT 66.090 -21.350 66.260 -20.470 ;
        RECT 66.680 -21.350 66.850 -20.470 ;
        RECT 68.350 -21.350 68.520 -20.470 ;
        RECT 70.750 -21.350 70.920 -20.470 ;
        RECT 71.340 -21.350 71.510 -20.470 ;
        RECT 71.930 -21.350 72.100 -20.470 ;
        RECT 33.750 -25.490 33.920 -24.610 ;
        RECT 35.040 -25.490 35.210 -24.610 ;
        RECT 38.250 -25.490 38.420 -24.610 ;
        RECT 49.900 -23.500 50.200 -23.300 ;
        RECT 39.540 -25.490 39.710 -24.610 ;
        RECT 49.720 -24.700 50.400 -24.500 ;
        RECT 52.960 -24.700 53.520 -24.460 ;
        RECT 69.570 -24.700 70.250 -24.500 ;
        RECT 72.810 -24.700 73.370 -24.460 ;
        RECT 17.140 -27.800 17.310 -26.920 ;
        RECT 20.145 -27.795 20.315 -26.915 ;
        RECT 43.230 -27.300 43.400 -25.020 ;
        RECT 44.720 -27.300 44.890 -25.020 ;
        RECT 46.210 -27.300 46.380 -25.020 ;
        RECT 47.700 -27.300 47.870 -25.020 ;
        RECT 49.190 -27.300 49.360 -25.020 ;
        RECT 50.680 -27.300 50.850 -25.020 ;
        RECT 52.430 -27.300 52.600 -25.020 ;
        RECT 53.920 -27.300 54.090 -25.020 ;
        RECT 55.410 -27.300 55.580 -25.020 ;
        RECT 56.900 -27.300 57.070 -25.020 ;
        RECT 58.390 -27.300 58.560 -25.020 ;
        RECT 59.880 -27.300 60.050 -25.020 ;
        RECT 63.080 -27.300 63.250 -25.020 ;
        RECT 64.570 -27.300 64.740 -25.020 ;
        RECT 66.060 -27.300 66.230 -25.020 ;
        RECT 67.550 -27.300 67.720 -25.020 ;
        RECT 69.040 -27.300 69.210 -25.020 ;
        RECT 70.530 -27.300 70.700 -25.020 ;
        RECT 72.280 -27.300 72.450 -25.020 ;
        RECT 73.770 -27.300 73.940 -25.020 ;
        RECT 75.260 -27.300 75.430 -25.020 ;
        RECT 76.750 -27.300 76.920 -25.020 ;
        RECT 78.240 -27.300 78.410 -25.020 ;
        RECT 79.730 -27.300 79.900 -25.020 ;
        RECT 17.140 -30.490 17.310 -29.610 ;
        RECT 22.950 -30.840 23.120 -28.760 ;
        RECT 25.530 -30.840 25.700 -28.760 ;
        RECT 28.110 -30.840 28.280 -28.760 ;
        RECT 30.690 -30.840 30.860 -28.760 ;
        RECT 33.270 -30.840 33.440 -28.760 ;
        RECT 35.850 -30.840 36.020 -28.760 ;
        RECT 40.040 -30.840 40.210 -29.960 ;
        RECT 43.310 -30.440 43.480 -28.850 ;
        RECT 45.890 -30.440 46.060 -28.850 ;
        RECT 49.690 -29.790 49.860 -28.910 ;
        RECT 53.480 -29.790 53.650 -28.910 ;
        RECT 56.880 -29.740 57.050 -28.860 ;
        RECT 50.000 -30.210 50.340 -30.040 ;
        RECT 53.000 -30.210 53.340 -30.040 ;
        RECT 55.900 -30.205 56.740 -30.035 ;
        RECT 46.750 -30.950 47.400 -30.750 ;
        RECT 59.880 -30.740 60.050 -28.860 ;
        RECT 63.160 -30.440 63.330 -28.850 ;
        RECT 65.740 -30.440 65.910 -28.850 ;
        RECT 69.540 -29.790 69.710 -28.910 ;
        RECT 73.330 -29.790 73.500 -28.910 ;
        RECT 76.730 -29.740 76.900 -28.860 ;
        RECT 69.850 -30.210 70.190 -30.040 ;
        RECT 72.850 -30.210 73.190 -30.040 ;
        RECT 75.750 -30.205 76.590 -30.035 ;
        RECT 66.600 -30.950 67.250 -30.750 ;
        RECT 79.730 -30.740 79.900 -28.860 ;
        RECT 23.260 -31.305 24.100 -31.135 ;
        RECT 24.550 -31.305 25.390 -31.135 ;
        RECT 25.840 -31.305 26.680 -31.135 ;
        RECT 27.130 -31.305 27.970 -31.135 ;
        RECT 28.420 -31.305 29.260 -31.135 ;
        RECT 29.710 -31.305 30.550 -31.135 ;
        RECT 31.000 -31.305 31.840 -31.135 ;
        RECT 32.290 -31.305 33.130 -31.135 ;
        RECT 33.580 -31.305 34.420 -31.135 ;
        RECT 34.870 -31.305 35.710 -31.135 ;
        RECT 36.160 -31.305 37.000 -31.135 ;
        RECT 39.060 -31.305 39.900 -31.135 ;
        RECT 58.900 -31.205 59.740 -31.035 ;
        RECT 78.750 -31.205 79.590 -31.035 ;
        RECT 48.400 -32.600 48.800 -32.400 ;
        RECT 68.250 -32.600 68.650 -32.400 ;
        RECT 23.260 -32.870 24.100 -32.700 ;
        RECT 24.550 -32.870 25.390 -32.700 ;
        RECT 25.840 -32.870 26.680 -32.700 ;
        RECT 27.130 -32.870 27.970 -32.700 ;
        RECT 28.420 -32.870 29.260 -32.700 ;
        RECT 29.710 -32.870 30.550 -32.700 ;
        RECT 31.000 -32.870 31.840 -32.700 ;
        RECT 32.290 -32.870 33.130 -32.700 ;
        RECT 33.580 -32.870 34.420 -32.700 ;
        RECT 34.870 -32.870 35.710 -32.700 ;
        RECT 36.160 -32.870 37.000 -32.700 ;
        RECT 17.140 -35.200 17.310 -34.320 ;
        RECT 20.145 -35.195 20.315 -34.315 ;
        RECT 24.240 -35.200 24.410 -33.120 ;
        RECT 26.820 -35.200 26.990 -33.120 ;
        RECT 29.400 -35.200 29.570 -33.120 ;
        RECT 31.980 -35.200 32.150 -33.120 ;
        RECT 34.560 -35.200 34.730 -33.120 ;
        RECT 37.140 -35.200 37.310 -33.120 ;
        RECT 39.060 -34.070 39.900 -33.900 ;
        RECT 40.040 -35.200 40.210 -34.320 ;
        RECT 45.270 -35.150 45.440 -32.770 ;
        RECT 47.850 -35.150 48.020 -32.770 ;
        RECT 50.430 -35.150 50.600 -32.770 ;
        RECT 53.010 -35.150 53.180 -32.770 ;
        RECT 55.590 -35.150 55.760 -32.770 ;
        RECT 65.120 -35.150 65.290 -32.770 ;
        RECT 67.700 -35.150 67.870 -32.770 ;
        RECT 70.280 -35.150 70.450 -32.770 ;
        RECT 72.860 -35.150 73.030 -32.770 ;
        RECT 75.440 -35.150 75.610 -32.770 ;
        RECT 43.950 -37.590 44.120 -36.710 ;
        RECT 44.540 -37.590 44.710 -36.710 ;
        RECT 45.130 -37.590 45.300 -36.710 ;
        RECT 46.800 -37.590 46.970 -36.710 ;
        RECT 47.390 -37.590 47.560 -36.710 ;
        RECT 47.980 -37.590 48.150 -36.710 ;
      LAYER met1 ;
        RECT -38.450 37.250 46.950 37.550 ;
        RECT -39.050 34.450 -38.750 34.480 ;
        RECT -38.450 34.450 -38.150 37.250 ;
        RECT -39.050 34.150 -38.150 34.450 ;
        RECT -37.850 36.750 45.550 37.050 ;
        RECT -39.050 34.120 -38.750 34.150 ;
        RECT -38.450 33.850 -38.150 33.880 ;
        RECT -37.850 33.850 -37.550 36.750 ;
        RECT -38.450 33.550 -37.550 33.850 ;
        RECT -37.350 36.250 40.450 36.550 ;
        RECT -38.450 33.520 -38.150 33.550 ;
        RECT -37.350 33.250 -37.050 36.250 ;
        RECT -37.880 32.950 -37.050 33.250 ;
        RECT -36.650 35.750 38.850 36.050 ;
        RECT -36.650 32.750 -36.350 35.750 ;
        RECT -37.380 32.450 -36.350 32.750 ;
        RECT -23.150 25.240 -20.100 25.250 ;
        RECT -16.700 25.240 -13.650 25.250 ;
        RECT -10.250 25.240 -7.200 25.250 ;
        RECT -3.800 25.240 -0.750 25.250 ;
        RECT 2.650 25.240 5.700 25.250 ;
        RECT 9.100 25.240 12.150 25.250 ;
        RECT 15.550 25.240 18.600 25.250 ;
        RECT 22.000 25.240 25.050 25.250 ;
        RECT 28.450 25.240 31.500 25.250 ;
        RECT 34.900 25.240 37.950 25.250 ;
        RECT -23.650 25.010 -20.100 25.240 ;
        RECT -17.200 25.010 -13.650 25.240 ;
        RECT -10.750 25.010 -7.200 25.240 ;
        RECT -4.300 25.010 -0.750 25.240 ;
        RECT 2.150 25.010 5.700 25.240 ;
        RECT 8.600 25.010 12.150 25.240 ;
        RECT 15.050 25.010 18.600 25.240 ;
        RECT 21.500 25.010 25.050 25.240 ;
        RECT 27.950 25.010 31.500 25.240 ;
        RECT 34.400 25.010 37.950 25.240 ;
        RECT -23.150 25.000 -20.100 25.010 ;
        RECT -16.700 25.000 -13.650 25.010 ;
        RECT -10.250 25.000 -7.200 25.010 ;
        RECT -3.800 25.000 -0.750 25.010 ;
        RECT 2.650 25.000 5.700 25.010 ;
        RECT 9.100 25.000 12.150 25.010 ;
        RECT 15.550 25.000 18.600 25.010 ;
        RECT 22.000 25.000 25.050 25.010 ;
        RECT 28.450 25.000 31.500 25.010 ;
        RECT 34.900 25.000 37.950 25.010 ;
        RECT -21.550 22.050 -21.200 22.100 ;
        RECT -23.100 22.040 -21.200 22.050 ;
        RECT -23.650 21.810 -21.200 22.040 ;
        RECT -23.100 21.800 -21.200 21.810 ;
        RECT -21.550 21.750 -21.200 21.800 ;
        RECT -20.350 20.500 -20.100 25.000 ;
        RECT -15.150 22.050 -14.800 22.100 ;
        RECT -16.700 22.040 -14.800 22.050 ;
        RECT -17.250 21.810 -14.800 22.040 ;
        RECT -16.700 21.800 -14.800 21.810 ;
        RECT -15.150 21.750 -14.800 21.800 ;
        RECT -13.900 20.500 -13.650 25.000 ;
        RECT -8.650 22.050 -8.300 22.100 ;
        RECT -10.200 22.040 -8.300 22.050 ;
        RECT -10.750 21.810 -8.300 22.040 ;
        RECT -10.200 21.800 -8.300 21.810 ;
        RECT -8.650 21.750 -8.300 21.800 ;
        RECT -7.450 20.500 -7.200 25.000 ;
        RECT -2.250 22.050 -1.900 22.100 ;
        RECT -3.800 22.040 -1.900 22.050 ;
        RECT -4.350 21.810 -1.900 22.040 ;
        RECT -3.800 21.800 -1.900 21.810 ;
        RECT -2.250 21.750 -1.900 21.800 ;
        RECT -1.000 20.500 -0.750 25.000 ;
        RECT 4.250 22.050 4.600 22.100 ;
        RECT 2.700 22.040 4.600 22.050 ;
        RECT 2.150 21.810 4.600 22.040 ;
        RECT 2.700 21.800 4.600 21.810 ;
        RECT 4.250 21.750 4.600 21.800 ;
        RECT 5.450 20.500 5.700 25.000 ;
        RECT 10.650 22.050 11.000 22.100 ;
        RECT 9.100 22.040 11.000 22.050 ;
        RECT 8.550 21.810 11.000 22.040 ;
        RECT 9.100 21.800 11.000 21.810 ;
        RECT 10.650 21.750 11.000 21.800 ;
        RECT 11.900 20.500 12.150 25.000 ;
        RECT 17.150 22.050 17.500 22.100 ;
        RECT 15.600 22.040 17.500 22.050 ;
        RECT 15.050 21.810 17.500 22.040 ;
        RECT 15.600 21.800 17.500 21.810 ;
        RECT 17.150 21.750 17.500 21.800 ;
        RECT 18.350 20.500 18.600 25.000 ;
        RECT 23.550 22.050 23.900 22.100 ;
        RECT 22.000 22.040 23.900 22.050 ;
        RECT 21.450 21.810 23.900 22.040 ;
        RECT 22.000 21.800 23.900 21.810 ;
        RECT 23.550 21.750 23.900 21.800 ;
        RECT 24.800 20.500 25.050 25.000 ;
        RECT 30.050 22.050 30.400 22.100 ;
        RECT 28.500 22.040 30.400 22.050 ;
        RECT 27.950 21.810 30.400 22.040 ;
        RECT 28.500 21.800 30.400 21.810 ;
        RECT 30.050 21.750 30.400 21.800 ;
        RECT 31.250 20.500 31.500 25.000 ;
        RECT 36.450 22.050 36.800 22.100 ;
        RECT 34.900 22.040 36.800 22.050 ;
        RECT 34.350 21.810 36.800 22.040 ;
        RECT 34.900 21.800 36.800 21.810 ;
        RECT 36.450 21.750 36.800 21.800 ;
        RECT 37.700 20.500 37.950 25.000 ;
        RECT 38.550 22.050 38.850 35.750 ;
        RECT 40.150 25.650 40.450 36.250 ;
        RECT 40.150 24.650 40.650 25.650 ;
        RECT 41.350 25.240 44.400 25.250 ;
        RECT 40.850 25.010 44.400 25.240 ;
        RECT 41.350 25.000 44.400 25.010 ;
        RECT 40.350 22.050 40.650 22.450 ;
        RECT 42.950 22.050 43.300 22.100 ;
        RECT 38.550 21.750 40.650 22.050 ;
        RECT 41.400 22.040 43.300 22.050 ;
        RECT 40.850 21.810 43.300 22.040 ;
        RECT 41.400 21.800 43.300 21.810 ;
        RECT 42.950 21.750 43.300 21.800 ;
        RECT 40.350 21.450 40.650 21.750 ;
        RECT 44.150 20.500 44.400 25.000 ;
        RECT 45.250 21.950 45.550 36.750 ;
        RECT 46.650 25.650 46.950 37.250 ;
        RECT 46.650 24.650 47.100 25.650 ;
        RECT 47.800 25.240 50.850 25.250 ;
        RECT 47.300 25.010 50.850 25.240 ;
        RECT 47.800 25.000 50.850 25.010 ;
        RECT 46.750 21.950 47.050 22.450 ;
        RECT 49.350 22.050 49.700 22.100 ;
        RECT 47.800 22.040 49.700 22.050 ;
        RECT 45.250 21.650 47.050 21.950 ;
        RECT 47.250 21.810 49.700 22.040 ;
        RECT 47.800 21.800 49.700 21.810 ;
        RECT 49.350 21.750 49.700 21.800 ;
        RECT 46.750 21.450 47.050 21.650 ;
        RECT 50.600 20.500 50.850 25.000 ;
        RECT -23.650 20.000 50.950 20.500 ;
        RECT -23.650 19.150 49.800 19.650 ;
        RECT -0.680 13.700 -0.450 13.740 ;
        RECT -1.200 12.800 -0.450 13.700 ;
        RECT -0.100 13.500 0.200 19.150 ;
        RECT 2.120 14.000 2.350 14.050 ;
        RECT -1.200 11.900 -0.900 12.800 ;
        RECT -0.680 12.740 -0.450 12.800 ;
        RECT -0.090 12.740 0.140 13.500 ;
        RECT 0.500 11.900 0.800 13.800 ;
        RECT 2.000 13.050 2.350 14.000 ;
        RECT 2.700 13.500 3.000 17.630 ;
        RECT 3.300 14.000 3.530 14.050 ;
        RECT 2.710 13.050 2.940 13.500 ;
        RECT 3.300 13.100 4.100 14.000 ;
        RECT 3.300 13.050 3.530 13.100 ;
        RECT 2.000 11.900 2.300 13.050 ;
        RECT 3.800 11.900 4.100 13.100 ;
        RECT 19.420 12.150 19.650 12.750 ;
        RECT -1.200 11.600 4.100 11.900 ;
        RECT 19.400 11.750 19.650 12.150 ;
        RECT 22.360 11.950 22.590 12.750 ;
        RECT 24.670 12.150 24.900 12.750 ;
        RECT 22.360 11.750 22.600 11.950 ;
        RECT 1.150 11.400 1.650 11.600 ;
        RECT 19.400 10.950 19.600 11.750 ;
        RECT 22.400 11.050 22.600 11.750 ;
        RECT 24.650 11.750 24.900 12.150 ;
        RECT 27.610 11.950 27.840 12.750 ;
        RECT 29.920 12.150 30.150 12.750 ;
        RECT 27.610 11.750 27.850 11.950 ;
        RECT 20.100 10.950 20.500 11.050 ;
        RECT 19.400 10.750 20.500 10.950 ;
        RECT 22.400 10.850 23.300 11.050 ;
        RECT -17.930 9.600 -17.470 10.000 ;
        RECT -17.900 8.900 -17.500 9.600 ;
        RECT -12.700 8.900 -12.300 10.730 ;
        RECT -1.900 10.050 -0.900 10.200 ;
        RECT -2.350 10.000 -0.900 10.050 ;
        RECT -7.500 9.600 -0.900 10.000 ;
        RECT -7.500 8.900 -7.100 9.600 ;
        RECT -2.350 9.350 -0.900 9.600 ;
        RECT -2.300 9.200 -0.900 9.350 ;
        RECT 19.400 9.590 19.600 10.750 ;
        RECT 20.100 10.650 20.500 10.750 ;
        RECT -2.300 8.900 -1.900 9.200 ;
        RECT 19.400 9.150 19.650 9.590 ;
        RECT 21.820 9.550 22.050 9.590 ;
        RECT -17.900 8.600 -15.400 8.900 ;
        RECT -12.700 8.600 -10.200 8.900 ;
        RECT -7.500 8.600 -5.000 8.900 ;
        RECT -2.300 8.600 0.200 8.900 ;
        RECT -17.100 8.300 -16.800 8.600 ;
        RECT -19.280 7.700 -19.050 8.300 ;
        RECT -19.300 7.300 -19.050 7.700 ;
        RECT -17.100 7.300 -16.750 8.300 ;
        RECT -16.340 7.500 -16.110 8.300 ;
        RECT -16.340 7.300 -16.100 7.500 ;
        RECT -15.700 7.300 -15.400 8.600 ;
        RECT -11.900 8.300 -11.600 8.600 ;
        RECT -14.080 7.700 -13.850 8.300 ;
        RECT -14.100 7.300 -13.850 7.700 ;
        RECT -11.900 7.300 -11.550 8.300 ;
        RECT -11.140 7.500 -10.910 8.300 ;
        RECT -11.140 7.300 -10.900 7.500 ;
        RECT -10.500 7.300 -10.200 8.600 ;
        RECT -6.700 8.300 -6.400 8.600 ;
        RECT -8.880 7.700 -8.650 8.300 ;
        RECT -8.900 7.300 -8.650 7.700 ;
        RECT -6.700 7.300 -6.350 8.300 ;
        RECT -5.940 7.500 -5.710 8.300 ;
        RECT -5.940 7.300 -5.700 7.500 ;
        RECT -5.300 7.300 -5.000 8.600 ;
        RECT -1.500 8.300 -1.200 8.600 ;
        RECT -3.680 7.700 -3.450 8.300 ;
        RECT -3.700 7.300 -3.450 7.700 ;
        RECT -1.500 7.300 -1.150 8.300 ;
        RECT -0.740 7.500 -0.510 8.300 ;
        RECT -0.740 7.300 -0.500 7.500 ;
        RECT -0.100 7.300 0.200 8.600 ;
        RECT 19.420 8.590 19.650 9.150 ;
        RECT 21.700 8.590 22.050 9.550 ;
        RECT 21.700 8.350 22.000 8.590 ;
        RECT 23.000 8.350 23.300 10.850 ;
        RECT 24.650 10.950 24.850 11.750 ;
        RECT 27.650 11.050 27.850 11.750 ;
        RECT 29.900 11.750 30.150 12.150 ;
        RECT 32.860 11.950 33.090 12.750 ;
        RECT 35.120 12.150 35.350 12.750 ;
        RECT 32.860 11.750 33.100 11.950 ;
        RECT 25.350 10.950 25.750 11.050 ;
        RECT 24.650 10.750 25.750 10.950 ;
        RECT 27.650 10.850 28.550 11.050 ;
        RECT 24.650 9.590 24.850 10.750 ;
        RECT 25.350 10.650 25.750 10.750 ;
        RECT 24.650 9.150 24.900 9.590 ;
        RECT 27.070 9.550 27.300 9.590 ;
        RECT 24.670 8.590 24.900 9.150 ;
        RECT 26.950 8.590 27.300 9.550 ;
        RECT 26.950 8.350 27.250 8.590 ;
        RECT 28.250 8.350 28.550 10.850 ;
        RECT 29.900 10.950 30.100 11.750 ;
        RECT 32.900 11.050 33.100 11.750 ;
        RECT 35.100 11.750 35.350 12.150 ;
        RECT 38.060 11.950 38.290 12.750 ;
        RECT 40.370 12.150 40.600 12.750 ;
        RECT 38.060 11.750 38.300 11.950 ;
        RECT 30.600 10.950 31.000 11.050 ;
        RECT 29.900 10.750 31.000 10.950 ;
        RECT 32.900 10.850 33.800 11.050 ;
        RECT 29.900 9.590 30.100 10.750 ;
        RECT 30.600 10.650 31.000 10.750 ;
        RECT 29.900 9.150 30.150 9.590 ;
        RECT 32.320 9.550 32.550 9.590 ;
        RECT 29.920 8.590 30.150 9.150 ;
        RECT 32.200 8.590 32.550 9.550 ;
        RECT 32.200 8.350 32.500 8.590 ;
        RECT 33.500 8.350 33.800 10.850 ;
        RECT 35.100 10.950 35.300 11.750 ;
        RECT 38.100 11.050 38.300 11.750 ;
        RECT 40.350 11.750 40.600 12.150 ;
        RECT 43.310 11.950 43.540 12.750 ;
        RECT 46.530 12.730 46.760 12.750 ;
        RECT 43.310 11.750 43.550 11.950 ;
        RECT 46.530 11.750 46.810 12.730 ;
        RECT 35.800 10.950 36.200 11.050 ;
        RECT 35.100 10.750 36.200 10.950 ;
        RECT 38.100 10.850 39.000 11.050 ;
        RECT 35.100 9.590 35.300 10.750 ;
        RECT 35.800 10.650 36.200 10.750 ;
        RECT 35.100 9.150 35.350 9.590 ;
        RECT 37.520 9.550 37.750 9.590 ;
        RECT 35.120 8.590 35.350 9.150 ;
        RECT 37.400 8.590 37.750 9.550 ;
        RECT 37.400 8.350 37.700 8.590 ;
        RECT 38.700 8.350 39.000 10.850 ;
        RECT 40.350 10.950 40.550 11.750 ;
        RECT 43.350 11.050 43.550 11.750 ;
        RECT 41.050 10.950 41.450 11.050 ;
        RECT 40.350 10.750 41.450 10.950 ;
        RECT 43.350 10.850 44.250 11.050 ;
        RECT 40.350 9.590 40.550 10.750 ;
        RECT 41.050 10.650 41.450 10.750 ;
        RECT 40.350 9.150 40.600 9.590 ;
        RECT 42.770 9.550 43.000 9.590 ;
        RECT 40.370 8.590 40.600 9.150 ;
        RECT 42.650 8.590 43.000 9.550 ;
        RECT 42.650 8.350 42.950 8.590 ;
        RECT 43.950 8.350 44.250 10.850 ;
        RECT 20.750 8.050 23.300 8.350 ;
        RECT 26.050 8.050 28.550 8.350 ;
        RECT 31.300 8.050 33.800 8.350 ;
        RECT 36.350 8.050 39.000 8.350 ;
        RECT 41.750 8.200 44.250 8.350 ;
        RECT 44.800 10.890 45.300 10.900 ;
        RECT 44.800 10.410 45.530 10.890 ;
        RECT 46.570 10.850 46.810 11.750 ;
        RECT 47.075 10.890 48.055 10.925 ;
        RECT 46.450 10.810 46.810 10.850 ;
        RECT 47.050 10.810 48.055 10.890 ;
        RECT 46.450 10.530 48.055 10.810 ;
        RECT 46.450 10.450 46.810 10.530 ;
        RECT 47.050 10.475 48.055 10.530 ;
        RECT 44.800 8.200 45.300 10.410 ;
        RECT 46.450 9.590 46.690 10.450 ;
        RECT 47.050 10.410 47.530 10.475 ;
        RECT 46.330 8.590 46.690 9.590 ;
        RECT 46.450 8.570 46.690 8.590 ;
        RECT 20.750 7.850 21.250 8.050 ;
        RECT -19.300 6.500 -19.100 7.300 ;
        RECT -18.600 6.500 -18.200 6.600 ;
        RECT -19.300 6.300 -18.200 6.500 ;
        RECT -19.300 5.140 -19.100 6.300 ;
        RECT -18.600 6.200 -18.200 6.300 ;
        RECT -17.100 6.200 -16.800 7.300 ;
        RECT -16.300 6.600 -16.100 7.300 ;
        RECT -16.300 6.400 -15.400 6.600 ;
        RECT -17.100 6.000 -16.100 6.200 ;
        RECT -16.300 5.140 -16.100 6.000 ;
        RECT -19.300 4.700 -19.050 5.140 ;
        RECT -16.880 5.100 -16.650 5.140 ;
        RECT -19.280 4.140 -19.050 4.700 ;
        RECT -17.000 4.140 -16.650 5.100 ;
        RECT -16.300 4.900 -16.060 5.140 ;
        RECT -16.290 4.140 -16.060 4.900 ;
        RECT -17.000 3.900 -16.700 4.140 ;
        RECT -15.700 3.900 -15.400 6.400 ;
        RECT -14.100 6.500 -13.900 7.300 ;
        RECT -13.400 6.500 -13.000 6.600 ;
        RECT -14.100 6.300 -13.000 6.500 ;
        RECT -14.100 5.140 -13.900 6.300 ;
        RECT -13.400 6.200 -13.000 6.300 ;
        RECT -11.900 6.200 -11.600 7.300 ;
        RECT -11.100 6.600 -10.900 7.300 ;
        RECT -11.100 6.400 -10.200 6.600 ;
        RECT -11.900 6.000 -10.900 6.200 ;
        RECT -11.100 5.140 -10.900 6.000 ;
        RECT -14.100 4.700 -13.850 5.140 ;
        RECT -11.680 5.100 -11.450 5.140 ;
        RECT -14.080 4.140 -13.850 4.700 ;
        RECT -11.800 4.140 -11.450 5.100 ;
        RECT -11.100 4.900 -10.860 5.140 ;
        RECT -11.090 4.140 -10.860 4.900 ;
        RECT -11.800 3.900 -11.500 4.140 ;
        RECT -10.500 3.900 -10.200 6.400 ;
        RECT -8.900 6.500 -8.700 7.300 ;
        RECT -8.200 6.500 -7.800 6.600 ;
        RECT -8.900 6.300 -7.800 6.500 ;
        RECT -8.900 5.140 -8.700 6.300 ;
        RECT -8.200 6.200 -7.800 6.300 ;
        RECT -6.700 6.200 -6.400 7.300 ;
        RECT -5.900 6.600 -5.700 7.300 ;
        RECT -5.900 6.400 -5.000 6.600 ;
        RECT -6.700 6.000 -5.700 6.200 ;
        RECT -5.900 5.140 -5.700 6.000 ;
        RECT -8.900 4.700 -8.650 5.140 ;
        RECT -6.480 5.100 -6.250 5.140 ;
        RECT -8.880 4.140 -8.650 4.700 ;
        RECT -6.600 4.140 -6.250 5.100 ;
        RECT -5.900 4.900 -5.660 5.140 ;
        RECT -5.890 4.140 -5.660 4.900 ;
        RECT -6.600 3.900 -6.300 4.140 ;
        RECT -5.300 3.900 -5.000 6.400 ;
        RECT -3.700 6.500 -3.500 7.300 ;
        RECT -3.000 6.500 -2.600 6.600 ;
        RECT -3.700 6.300 -2.600 6.500 ;
        RECT -3.700 5.140 -3.500 6.300 ;
        RECT -3.000 6.200 -2.600 6.300 ;
        RECT -1.500 6.200 -1.200 7.300 ;
        RECT -0.700 6.600 -0.500 7.300 ;
        RECT 20.770 7.230 21.225 7.850 ;
        RECT 26.050 7.250 26.450 8.050 ;
        RECT 31.300 7.750 31.700 8.050 ;
        RECT 36.350 7.825 36.900 8.050 ;
        RECT 20.740 6.775 21.255 7.230 ;
        RECT 25.950 6.650 26.550 7.250 ;
        RECT -0.700 6.400 0.200 6.600 ;
        RECT -1.500 6.000 -0.500 6.200 ;
        RECT -0.700 5.140 -0.500 6.000 ;
        RECT -3.700 4.700 -3.450 5.140 ;
        RECT -1.280 5.100 -1.050 5.140 ;
        RECT -3.680 4.140 -3.450 4.700 ;
        RECT -1.400 4.140 -1.050 5.100 ;
        RECT -0.700 4.900 -0.460 5.140 ;
        RECT -0.690 4.140 -0.460 4.900 ;
        RECT -1.400 3.900 -1.100 4.140 ;
        RECT -0.100 3.900 0.200 6.400 ;
        RECT -17.900 3.600 -15.400 3.900 ;
        RECT -12.700 3.600 -10.200 3.900 ;
        RECT -7.500 3.600 -5.000 3.900 ;
        RECT -2.300 3.600 0.200 3.900 ;
        RECT -17.900 3.400 -17.500 3.600 ;
        RECT -12.700 3.400 -12.300 3.600 ;
        RECT -17.900 3.100 -12.200 3.400 ;
        RECT -12.600 0.900 -12.200 3.100 ;
        RECT -7.500 1.900 -7.100 3.600 ;
        RECT -6.600 1.900 -6.200 1.930 ;
        RECT -8.300 1.200 -7.900 1.730 ;
        RECT -7.500 1.500 -6.200 1.900 ;
        RECT -6.600 1.470 -6.200 1.500 ;
        RECT -2.300 1.200 -1.900 3.600 ;
        RECT 31.325 1.675 31.675 7.750 ;
        RECT 36.325 7.400 36.900 7.825 ;
        RECT 41.750 7.750 45.300 8.200 ;
        RECT 36.325 1.825 36.775 7.400 ;
        RECT 31.325 1.325 34.650 1.675 ;
        RECT 36.295 1.375 36.805 1.825 ;
        RECT -12.600 0.400 -10.920 0.900 ;
        RECT -8.300 0.800 -1.900 1.200 ;
        RECT -12.600 -0.100 -12.200 0.400 ;
        RECT -19.520 -1.000 -13.080 -0.480 ;
        RECT -12.600 -0.880 -12.250 -0.100 ;
        RECT -9.500 -0.300 0.080 0.100 ;
        RECT -19.520 -1.460 -19.080 -1.000 ;
        RECT -16.320 -1.460 -16.080 -1.000 ;
        RECT -19.520 -3.860 -19.050 -1.460 ;
        RECT -17.790 -3.240 -17.560 -1.460 ;
        RECT -16.320 -1.640 -16.070 -1.460 ;
        RECT -19.520 -4.600 -19.080 -3.860 ;
        RECT -17.800 -4.040 -17.560 -3.240 ;
        RECT -16.300 -3.860 -16.070 -1.640 ;
        RECT -14.810 -3.240 -14.580 -1.460 ;
        RECT -13.320 -1.640 -13.080 -1.000 ;
        RECT -12.800 -1.240 -12.080 -0.880 ;
        RECT -9.450 -0.920 -9.100 -0.300 ;
        RECT -0.850 -0.400 0.080 -0.300 ;
        RECT 2.500 0.000 11.250 0.250 ;
        RECT 12.545 0.125 14.400 0.475 ;
        RECT 2.500 -0.275 3.750 0.000 ;
        RECT -9.680 -1.240 -8.840 -0.920 ;
        RECT -8.640 -0.960 -8.000 -0.480 ;
        RECT -7.920 -0.960 -2.400 -0.480 ;
        RECT -8.640 -1.000 -2.400 -0.960 ;
        RECT -14.810 -3.860 -14.560 -3.240 ;
        RECT -13.320 -3.860 -13.090 -1.640 ;
        RECT -11.830 -3.240 -11.600 -1.460 ;
        RECT -14.800 -4.040 -14.560 -3.860 ;
        RECT -11.840 -4.040 -11.600 -3.240 ;
        RECT -10.080 -3.280 -9.850 -1.460 ;
        RECT -8.600 -1.560 -8.360 -1.000 ;
        RECT -5.600 -1.460 -5.360 -1.000 ;
        RECT -17.800 -4.240 -11.600 -4.040 ;
        RECT -10.120 -3.860 -9.850 -3.280 ;
        RECT -8.590 -3.860 -8.360 -1.560 ;
        RECT -7.100 -3.360 -6.870 -1.460 ;
        RECT -7.120 -3.860 -6.870 -3.360 ;
        RECT -5.610 -1.560 -5.360 -1.460 ;
        RECT -5.610 -3.860 -5.380 -1.560 ;
        RECT -4.120 -3.320 -3.890 -1.460 ;
        RECT -2.640 -1.520 -2.400 -1.000 ;
        RECT -10.120 -4.040 -9.880 -3.860 ;
        RECT -7.120 -4.040 -6.880 -3.860 ;
        RECT -4.120 -4.040 -3.880 -3.320 ;
        RECT -2.630 -3.860 -2.400 -1.520 ;
        RECT -10.120 -4.240 -3.880 -4.040 ;
        RECT -19.520 -5.120 -16.440 -4.600 ;
        RECT -19.280 -5.720 -19.050 -5.300 ;
        RECT -20.000 -6.960 -19.050 -5.720 ;
        RECT -16.960 -5.320 -16.440 -5.120 ;
        RECT -16.280 -5.320 -16.050 -5.300 ;
        RECT -16.960 -6.160 -16.050 -5.320 ;
        RECT -16.280 -6.300 -16.050 -6.160 ;
        RECT -12.880 -6.480 -12.640 -4.240 ;
        RECT -9.080 -5.350 -8.800 -4.240 ;
        RECT -9.090 -5.550 -8.800 -5.350 ;
        RECT -9.090 -6.000 -7.600 -5.550 ;
        RECT -9.090 -6.350 -8.860 -6.000 ;
        RECT -19.900 -8.550 -19.500 -6.960 ;
        RECT -19.280 -7.300 -19.050 -6.960 ;
        RECT -17.400 -6.500 -15.040 -6.480 ;
        RECT -17.400 -6.680 -13.900 -6.500 ;
        RECT -19.240 -7.480 -19.080 -7.300 ;
        RECT -17.400 -7.480 -17.160 -6.680 ;
        RECT -16.000 -6.735 -13.900 -6.680 ;
        RECT -12.880 -6.510 -12.440 -6.480 ;
        RECT -12.880 -6.520 -12.140 -6.510 ;
        RECT -9.600 -6.520 -9.140 -6.510 ;
        RECT -12.880 -6.720 -9.120 -6.520 ;
        RECT -15.500 -6.750 -13.900 -6.735 ;
        RECT -12.600 -6.740 -12.140 -6.720 ;
        RECT -9.600 -6.740 -9.140 -6.720 ;
        RECT -14.100 -7.200 -13.900 -6.750 ;
        RECT -5.290 -6.800 -5.060 -5.290 ;
        RECT -2.710 -5.300 -2.480 -5.290 ;
        RECT -14.100 -7.400 -5.800 -7.200 ;
        RECT -19.240 -7.760 -17.160 -7.480 ;
        RECT -6.700 -7.500 -5.800 -7.400 ;
        RECT -5.400 -7.600 -5.000 -6.800 ;
        RECT -2.710 -7.000 -2.400 -5.300 ;
        RECT -2.700 -7.600 -2.400 -7.000 ;
        RECT -5.400 -7.650 -2.400 -7.600 ;
        RECT 0.600 -7.300 2.300 -7.000 ;
        RECT 0.600 -7.550 0.900 -7.300 ;
        RECT 2.000 -7.550 2.300 -7.300 ;
        RECT -5.400 -7.900 -1.750 -7.650 ;
        RECT 0.600 -7.900 0.950 -7.550 ;
        RECT -4.800 -8.200 -4.400 -7.900 ;
        RECT -15.000 -8.500 -4.400 -8.200 ;
        RECT -2.850 -8.400 -1.750 -7.900 ;
        RECT -1.530 -8.300 0.950 -7.900 ;
        RECT 1.310 -8.100 1.540 -7.550 ;
        RECT -19.900 -8.950 -18.270 -8.550 ;
        RECT -15.000 -9.400 -14.750 -8.500 ;
        RECT -12.450 -9.210 -12.200 -8.500 ;
        RECT -14.990 -11.710 -14.760 -9.400 ;
        RECT -12.450 -9.450 -12.180 -9.210 ;
        RECT -9.850 -9.450 -9.600 -8.500 ;
        RECT -8.100 -9.150 -7.500 -8.650 ;
        RECT -12.410 -11.710 -12.180 -9.450 ;
        RECT -9.830 -11.710 -9.600 -9.450 ;
        RECT -7.250 -9.450 -7.000 -8.500 ;
        RECT -4.650 -9.210 -4.400 -8.500 ;
        RECT 0.720 -8.550 0.950 -8.300 ;
        RECT -7.250 -11.710 -7.020 -9.450 ;
        RECT -4.670 -9.500 -4.400 -9.210 ;
        RECT 1.300 -9.100 1.600 -8.100 ;
        RECT 1.900 -8.300 2.300 -7.550 ;
        RECT 1.900 -8.550 2.130 -8.300 ;
        RECT 2.500 -9.100 2.750 -0.275 ;
        RECT 3.200 -0.300 3.750 -0.275 ;
        RECT 3.980 -1.000 10.420 -0.480 ;
        RECT 10.900 -0.880 11.250 0.000 ;
        RECT 3.980 -1.460 4.420 -1.000 ;
        RECT 7.180 -1.460 7.420 -1.000 ;
        RECT 3.980 -3.860 4.450 -1.460 ;
        RECT 5.710 -3.240 5.940 -1.460 ;
        RECT 7.180 -1.640 7.430 -1.460 ;
        RECT 3.980 -4.600 4.420 -3.860 ;
        RECT 5.700 -4.040 5.940 -3.240 ;
        RECT 7.200 -3.860 7.430 -1.640 ;
        RECT 8.690 -3.240 8.920 -1.460 ;
        RECT 10.180 -1.640 10.420 -1.000 ;
        RECT 10.700 -1.240 11.420 -0.880 ;
        RECT 14.050 -0.920 14.400 0.125 ;
        RECT 22.075 0.075 31.475 0.425 ;
        RECT 13.820 -1.240 14.660 -0.920 ;
        RECT 14.860 -0.960 15.500 -0.480 ;
        RECT 15.580 -0.960 21.100 -0.480 ;
        RECT 14.860 -1.000 21.100 -0.960 ;
        RECT 8.690 -3.860 8.940 -3.240 ;
        RECT 10.180 -3.860 10.410 -1.640 ;
        RECT 11.670 -3.240 11.900 -1.460 ;
        RECT 8.700 -4.040 8.940 -3.860 ;
        RECT 11.660 -4.040 11.900 -3.240 ;
        RECT 13.420 -3.280 13.650 -1.460 ;
        RECT 14.900 -1.560 15.140 -1.000 ;
        RECT 17.900 -1.460 18.140 -1.000 ;
        RECT 5.700 -4.240 11.900 -4.040 ;
        RECT 13.380 -3.860 13.650 -3.280 ;
        RECT 14.910 -3.860 15.140 -1.560 ;
        RECT 16.400 -3.360 16.630 -1.460 ;
        RECT 16.380 -3.860 16.630 -3.360 ;
        RECT 17.890 -1.560 18.140 -1.460 ;
        RECT 17.890 -3.860 18.120 -1.560 ;
        RECT 19.380 -3.320 19.610 -1.460 ;
        RECT 20.860 -1.520 21.100 -1.000 ;
        RECT 13.380 -4.040 13.620 -3.860 ;
        RECT 16.380 -4.040 16.620 -3.860 ;
        RECT 19.380 -4.040 19.620 -3.320 ;
        RECT 20.870 -3.860 21.100 -1.520 ;
        RECT 13.380 -4.240 19.620 -4.040 ;
        RECT 3.980 -5.120 7.060 -4.600 ;
        RECT 4.220 -5.720 4.450 -5.300 ;
        RECT 3.500 -6.960 4.450 -5.720 ;
        RECT 6.540 -5.320 7.060 -5.120 ;
        RECT 7.220 -5.320 7.450 -5.300 ;
        RECT 6.540 -6.160 7.450 -5.320 ;
        RECT 7.220 -6.300 7.450 -6.160 ;
        RECT 10.620 -6.480 10.860 -4.240 ;
        RECT 14.420 -5.350 14.700 -4.240 ;
        RECT 14.410 -5.550 14.700 -5.350 ;
        RECT 14.410 -6.000 15.900 -5.550 ;
        RECT 14.410 -6.350 14.640 -6.000 ;
        RECT 3.500 -8.650 3.900 -6.960 ;
        RECT 4.220 -7.300 4.450 -6.960 ;
        RECT 6.100 -6.500 8.460 -6.480 ;
        RECT 6.100 -6.680 9.600 -6.500 ;
        RECT 4.260 -7.480 4.420 -7.300 ;
        RECT 6.100 -7.480 6.340 -6.680 ;
        RECT 7.500 -6.735 9.600 -6.680 ;
        RECT 10.620 -6.510 11.060 -6.480 ;
        RECT 10.620 -6.520 11.360 -6.510 ;
        RECT 13.900 -6.520 14.360 -6.510 ;
        RECT 10.620 -6.720 14.380 -6.520 ;
        RECT 8.000 -6.750 9.600 -6.735 ;
        RECT 10.900 -6.740 11.360 -6.720 ;
        RECT 13.900 -6.740 14.360 -6.720 ;
        RECT 9.400 -7.200 9.600 -6.750 ;
        RECT 18.210 -6.800 18.440 -5.290 ;
        RECT 20.790 -5.300 21.020 -5.290 ;
        RECT 9.400 -7.400 17.700 -7.200 ;
        RECT 4.260 -7.760 6.340 -7.480 ;
        RECT 16.800 -7.500 17.700 -7.400 ;
        RECT 18.100 -7.600 18.500 -6.800 ;
        RECT 20.790 -7.000 21.100 -5.300 ;
        RECT 20.800 -7.600 21.100 -7.000 ;
        RECT 18.100 -7.650 21.100 -7.600 ;
        RECT 18.100 -7.900 21.750 -7.650 ;
        RECT 22.075 -7.900 22.425 0.075 ;
        RECT 31.125 0.050 31.475 0.075 ;
        RECT 34.300 0.350 34.650 1.325 ;
        RECT 34.300 0.325 37.100 0.350 ;
        RECT 31.125 -0.275 31.500 0.050 ;
        RECT 24.230 -1.000 30.670 -0.480 ;
        RECT 31.150 -0.880 31.500 -0.275 ;
        RECT 34.300 -0.025 43.875 0.325 ;
        RECT 34.300 -0.050 37.100 -0.025 ;
        RECT 24.230 -1.460 24.670 -1.000 ;
        RECT 27.430 -1.460 27.670 -1.000 ;
        RECT 24.230 -3.860 24.700 -1.460 ;
        RECT 25.960 -3.240 26.190 -1.460 ;
        RECT 27.430 -1.640 27.680 -1.460 ;
        RECT 24.230 -4.600 24.670 -3.860 ;
        RECT 25.950 -4.040 26.190 -3.240 ;
        RECT 27.450 -3.860 27.680 -1.640 ;
        RECT 28.940 -3.240 29.170 -1.460 ;
        RECT 30.430 -1.640 30.670 -1.000 ;
        RECT 30.950 -1.240 31.670 -0.880 ;
        RECT 34.300 -0.920 34.650 -0.050 ;
        RECT 34.070 -1.240 34.910 -0.920 ;
        RECT 35.110 -0.960 35.750 -0.480 ;
        RECT 35.830 -0.960 41.350 -0.480 ;
        RECT 35.110 -1.000 41.350 -0.960 ;
        RECT 28.940 -3.860 29.190 -3.240 ;
        RECT 30.430 -3.860 30.660 -1.640 ;
        RECT 31.920 -3.240 32.150 -1.460 ;
        RECT 28.950 -4.040 29.190 -3.860 ;
        RECT 31.910 -4.040 32.150 -3.240 ;
        RECT 33.670 -3.280 33.900 -1.460 ;
        RECT 35.150 -1.560 35.390 -1.000 ;
        RECT 38.150 -1.460 38.390 -1.000 ;
        RECT 25.950 -4.240 32.150 -4.040 ;
        RECT 33.630 -3.860 33.900 -3.280 ;
        RECT 35.160 -3.860 35.390 -1.560 ;
        RECT 36.650 -3.360 36.880 -1.460 ;
        RECT 36.630 -3.860 36.880 -3.360 ;
        RECT 38.140 -1.560 38.390 -1.460 ;
        RECT 38.140 -3.860 38.370 -1.560 ;
        RECT 39.630 -3.320 39.860 -1.460 ;
        RECT 41.110 -1.520 41.350 -1.000 ;
        RECT 33.630 -4.040 33.870 -3.860 ;
        RECT 36.630 -4.040 36.870 -3.860 ;
        RECT 39.630 -4.040 39.870 -3.320 ;
        RECT 41.120 -3.860 41.350 -1.520 ;
        RECT 33.630 -4.240 39.870 -4.040 ;
        RECT 24.230 -5.120 27.310 -4.600 ;
        RECT 24.470 -5.720 24.700 -5.300 ;
        RECT 23.750 -6.200 24.700 -5.720 ;
        RECT 26.790 -5.320 27.310 -5.120 ;
        RECT 27.470 -5.320 27.700 -5.300 ;
        RECT 26.790 -6.160 27.700 -5.320 ;
        RECT 23.270 -6.600 24.700 -6.200 ;
        RECT 27.470 -6.300 27.700 -6.160 ;
        RECT 30.870 -6.480 31.110 -4.240 ;
        RECT 34.670 -5.350 34.950 -4.240 ;
        RECT 34.660 -5.550 34.950 -5.350 ;
        RECT 34.660 -6.000 36.150 -5.550 ;
        RECT 34.660 -6.350 34.890 -6.000 ;
        RECT 23.750 -6.960 24.700 -6.600 ;
        RECT 24.470 -7.300 24.700 -6.960 ;
        RECT 26.350 -6.500 28.710 -6.480 ;
        RECT 26.350 -6.680 29.850 -6.500 ;
        RECT 24.510 -7.480 24.670 -7.300 ;
        RECT 26.350 -7.480 26.590 -6.680 ;
        RECT 27.750 -6.735 29.850 -6.680 ;
        RECT 30.870 -6.510 31.310 -6.480 ;
        RECT 30.870 -6.520 31.610 -6.510 ;
        RECT 34.150 -6.520 34.610 -6.510 ;
        RECT 30.870 -6.720 34.630 -6.520 ;
        RECT 28.250 -6.750 29.850 -6.735 ;
        RECT 31.150 -6.740 31.610 -6.720 ;
        RECT 34.150 -6.740 34.610 -6.720 ;
        RECT 29.650 -7.200 29.850 -6.750 ;
        RECT 38.460 -6.800 38.690 -5.290 ;
        RECT 41.040 -5.300 41.270 -5.290 ;
        RECT 29.650 -7.400 37.950 -7.200 ;
        RECT 24.510 -7.760 26.590 -7.480 ;
        RECT 37.050 -7.500 37.950 -7.400 ;
        RECT 38.350 -7.600 38.750 -6.800 ;
        RECT 41.040 -7.000 41.350 -5.300 ;
        RECT 41.050 -7.600 41.350 -7.000 ;
        RECT 38.350 -7.650 41.350 -7.600 ;
        RECT 38.350 -7.900 42.000 -7.650 ;
        RECT 18.700 -8.200 19.100 -7.900 ;
        RECT 8.500 -8.500 19.100 -8.200 ;
        RECT 20.650 -8.250 22.425 -7.900 ;
        RECT 38.950 -8.200 39.350 -7.900 ;
        RECT 20.650 -8.400 21.750 -8.250 ;
        RECT 3.500 -9.050 6.380 -8.650 ;
        RECT 1.300 -9.250 2.750 -9.100 ;
        RECT 1.300 -9.400 2.500 -9.250 ;
        RECT 8.500 -9.400 8.750 -8.500 ;
        RECT 11.050 -9.210 11.300 -8.500 ;
        RECT -4.670 -11.710 -4.440 -9.500 ;
        RECT 8.510 -11.710 8.740 -9.400 ;
        RECT 11.050 -9.450 11.320 -9.210 ;
        RECT 13.650 -9.450 13.900 -8.500 ;
        RECT 15.400 -9.150 16.000 -8.650 ;
        RECT 11.090 -11.710 11.320 -9.450 ;
        RECT 13.670 -11.710 13.900 -9.450 ;
        RECT 16.250 -9.450 16.500 -8.500 ;
        RECT 18.850 -9.210 19.100 -8.500 ;
        RECT 16.250 -11.710 16.480 -9.450 ;
        RECT 18.830 -9.500 19.100 -9.210 ;
        RECT 28.750 -8.500 39.350 -8.200 ;
        RECT 40.900 -8.400 42.000 -7.900 ;
        RECT 28.750 -9.400 29.000 -8.500 ;
        RECT 31.300 -9.210 31.550 -8.500 ;
        RECT 18.830 -11.710 19.060 -9.500 ;
        RECT 28.760 -11.710 28.990 -9.400 ;
        RECT 31.300 -9.450 31.570 -9.210 ;
        RECT 33.900 -9.450 34.150 -8.500 ;
        RECT 35.650 -9.150 36.250 -8.650 ;
        RECT 31.340 -11.710 31.570 -9.450 ;
        RECT 33.920 -11.710 34.150 -9.450 ;
        RECT 36.500 -9.450 36.750 -8.500 ;
        RECT 39.100 -9.210 39.350 -8.500 ;
        RECT 36.500 -11.710 36.730 -9.450 ;
        RECT 39.080 -9.500 39.350 -9.210 ;
        RECT 39.080 -11.710 39.310 -9.500 ;
        RECT 43.525 -14.675 43.875 -0.025 ;
        RECT -44.000 -20.000 -37.000 -15.000 ;
        RECT 43.525 -15.025 68.800 -14.675 ;
        RECT 68.450 -16.150 68.800 -15.025 ;
        RECT 64.450 -16.450 70.100 -16.150 ;
        RECT 64.450 -16.650 64.850 -16.450 ;
        RECT 69.700 -16.650 70.100 -16.450 ;
        RECT 64.450 -16.950 66.950 -16.650 ;
        RECT 69.700 -16.950 72.200 -16.650 ;
        RECT 65.250 -17.250 65.550 -16.950 ;
        RECT 61.180 -17.270 61.410 -17.250 ;
        RECT 61.180 -18.250 61.460 -17.270 ;
        RECT 63.070 -17.850 63.300 -17.250 ;
        RECT 22.200 -19.150 22.700 -19.120 ;
        RECT 61.220 -19.150 61.460 -18.250 ;
        RECT 63.050 -18.250 63.300 -17.850 ;
        RECT 65.250 -18.250 65.600 -17.250 ;
        RECT 66.010 -18.050 66.240 -17.250 ;
        RECT 66.010 -18.250 66.250 -18.050 ;
        RECT 66.650 -18.250 66.950 -16.950 ;
        RECT 70.500 -17.250 70.800 -16.950 ;
        RECT 68.320 -17.850 68.550 -17.250 ;
        RECT 68.300 -18.250 68.550 -17.850 ;
        RECT 70.500 -18.250 70.850 -17.250 ;
        RECT 71.260 -18.050 71.490 -17.250 ;
        RECT 71.260 -18.250 71.500 -18.050 ;
        RECT 71.900 -18.250 72.200 -16.950 ;
        RECT 62.000 -19.110 62.400 -19.000 ;
        RECT -0.480 -19.650 22.700 -19.150 ;
        RECT 22.200 -19.680 22.700 -19.650 ;
        RECT 61.100 -19.190 61.460 -19.150 ;
        RECT 61.700 -19.190 62.400 -19.110 ;
        RECT 61.100 -19.470 62.400 -19.190 ;
        RECT 61.100 -19.550 61.460 -19.470 ;
        RECT 5.920 -20.450 19.780 -20.050 ;
        RECT 61.100 -20.410 61.340 -19.550 ;
        RECT 61.700 -19.590 62.400 -19.470 ;
        RECT 62.000 -19.600 62.400 -19.590 ;
        RECT 63.050 -19.050 63.250 -18.250 ;
        RECT 63.750 -19.050 64.150 -18.950 ;
        RECT 63.050 -19.250 64.150 -19.050 ;
        RECT -18.700 -20.650 -18.300 -20.620 ;
        RECT -18.700 -21.050 18.850 -20.650 ;
        RECT -18.700 -21.080 -18.300 -21.050 ;
        RECT 18.450 -21.600 18.850 -21.050 ;
        RECT 18.300 -22.000 21.100 -21.600 ;
        RECT 33.720 -21.710 33.950 -20.710 ;
        RECT 39.510 -21.710 39.740 -20.710 ;
        RECT 60.980 -21.410 61.340 -20.410 ;
        RECT 63.050 -20.410 63.250 -19.250 ;
        RECT 63.750 -19.350 64.150 -19.250 ;
        RECT 65.250 -19.350 65.550 -18.250 ;
        RECT 66.050 -18.950 66.250 -18.250 ;
        RECT 66.050 -19.150 66.950 -18.950 ;
        RECT 65.250 -19.550 66.250 -19.350 ;
        RECT 66.050 -20.410 66.250 -19.550 ;
        RECT 63.050 -20.850 63.300 -20.410 ;
        RECT 65.470 -20.450 65.700 -20.410 ;
        RECT 63.070 -21.410 63.300 -20.850 ;
        RECT 65.350 -21.410 65.700 -20.450 ;
        RECT 66.050 -20.650 66.290 -20.410 ;
        RECT 66.060 -21.410 66.290 -20.650 ;
        RECT 61.100 -21.430 61.340 -21.410 ;
        RECT 65.350 -21.650 65.650 -21.410 ;
        RECT 66.650 -21.650 66.950 -19.150 ;
        RECT 68.300 -19.050 68.500 -18.250 ;
        RECT 69.000 -19.050 69.400 -18.950 ;
        RECT 68.300 -19.250 69.400 -19.050 ;
        RECT 68.300 -20.410 68.500 -19.250 ;
        RECT 69.000 -19.350 69.400 -19.250 ;
        RECT 70.500 -19.350 70.800 -18.250 ;
        RECT 71.300 -18.950 71.500 -18.250 ;
        RECT 71.300 -19.150 72.200 -18.950 ;
        RECT 70.500 -19.550 71.500 -19.350 ;
        RECT 71.300 -20.410 71.500 -19.550 ;
        RECT 68.300 -20.850 68.550 -20.410 ;
        RECT 70.720 -20.450 70.950 -20.410 ;
        RECT 68.320 -21.410 68.550 -20.850 ;
        RECT 70.600 -21.410 70.950 -20.450 ;
        RECT 71.300 -20.650 71.540 -20.410 ;
        RECT 71.310 -21.410 71.540 -20.650 ;
        RECT 70.600 -21.650 70.900 -21.410 ;
        RECT 71.900 -21.650 72.200 -19.150 ;
        RECT 64.450 -21.950 66.950 -21.650 ;
        RECT 69.700 -21.950 72.200 -21.650 ;
        RECT 64.450 -22.000 64.850 -21.950 ;
        RECT 17.110 -22.500 17.340 -22.150 ;
        RECT 18.300 -22.500 18.700 -22.000 ;
        RECT 17.110 -22.900 18.700 -22.500 ;
        RECT 40.500 -22.500 64.850 -22.000 ;
        RECT 17.110 -23.150 17.340 -22.900 ;
        RECT 19.350 -23.100 19.750 -23.070 ;
        RECT 18.400 -23.500 21.100 -23.100 ;
        RECT 40.500 -23.450 41.000 -22.500 ;
        RECT 18.400 -24.100 18.800 -23.500 ;
        RECT 19.350 -23.530 19.750 -23.500 ;
        RECT 22.170 -23.950 41.000 -23.450 ;
        RECT 41.450 -22.950 53.400 -22.700 ;
        RECT 69.700 -22.850 70.100 -21.950 ;
        RECT 17.200 -24.500 18.800 -24.100 ;
        RECT 36.600 -24.120 37.100 -23.950 ;
        RECT 23.300 -24.300 23.700 -24.270 ;
        RECT 17.200 -26.860 17.600 -24.500 ;
        RECT 20.200 -24.700 23.700 -24.300 ;
        RECT 20.200 -26.855 20.600 -24.700 ;
        RECT 23.300 -24.730 23.700 -24.700 ;
        RECT 33.720 -25.550 33.950 -24.550 ;
        RECT 35.010 -25.550 35.240 -24.550 ;
        RECT 36.540 -24.680 37.160 -24.120 ;
        RECT 38.220 -25.550 38.450 -24.550 ;
        RECT 39.510 -25.550 39.740 -24.550 ;
        RECT 17.110 -27.860 17.600 -26.860 ;
        RECT 20.115 -27.855 20.600 -26.855 ;
        RECT 17.200 -27.900 17.600 -27.860 ;
        RECT 20.200 -27.900 20.600 -27.855 ;
        RECT 18.300 -29.400 21.250 -29.000 ;
        RECT 17.110 -29.900 17.340 -29.550 ;
        RECT 18.300 -29.900 18.700 -29.400 ;
        RECT 20.500 -29.500 21.250 -29.400 ;
        RECT 17.110 -30.300 18.700 -29.900 ;
        RECT 17.110 -30.550 17.340 -30.300 ;
        RECT 18.400 -30.900 21.100 -30.500 ;
        RECT 22.920 -30.600 23.150 -28.700 ;
        RECT 25.500 -30.600 25.730 -28.700 ;
        RECT 28.080 -30.600 28.310 -28.700 ;
        RECT 30.660 -30.600 30.890 -28.700 ;
        RECT 33.240 -30.600 33.470 -28.700 ;
        RECT 35.820 -30.600 36.050 -28.700 ;
        RECT 18.400 -31.500 18.800 -30.900 ;
        RECT 19.250 -31.000 20.000 -30.900 ;
        RECT 22.800 -31.000 23.200 -30.600 ;
        RECT 17.200 -31.900 18.800 -31.500 ;
        RECT 21.600 -31.100 23.200 -31.000 ;
        RECT 25.500 -31.100 25.800 -30.600 ;
        RECT 28.000 -30.900 28.310 -30.600 ;
        RECT 28.000 -31.100 28.300 -30.900 ;
        RECT 30.600 -31.100 30.900 -30.600 ;
        RECT 33.200 -31.100 33.500 -30.600 ;
        RECT 35.800 -31.100 36.100 -30.600 ;
        RECT 40.010 -30.900 40.400 -29.900 ;
        RECT 21.600 -31.105 39.800 -31.100 ;
        RECT 21.600 -31.335 39.960 -31.105 ;
        RECT 21.600 -31.400 39.800 -31.335 ;
        RECT 21.600 -31.700 22.000 -31.400 ;
        RECT 17.200 -34.260 17.600 -31.900 ;
        RECT 20.200 -32.100 22.000 -31.700 ;
        RECT 20.200 -34.255 20.600 -32.100 ;
        RECT 40.100 -32.300 40.400 -30.900 ;
        RECT 37.100 -32.600 40.400 -32.300 ;
        RECT 23.200 -32.900 37.400 -32.600 ;
        RECT 24.200 -33.700 24.500 -32.900 ;
        RECT 26.700 -33.060 27.000 -32.900 ;
        RECT 26.700 -33.700 27.020 -33.060 ;
        RECT 29.300 -33.700 29.600 -32.900 ;
        RECT 31.900 -33.700 32.200 -32.900 ;
        RECT 34.500 -33.700 34.800 -32.900 ;
        RECT 37.100 -33.700 37.400 -32.900 ;
        RECT 17.110 -35.260 17.600 -34.260 ;
        RECT 20.115 -35.255 20.600 -34.255 ;
        RECT 17.200 -35.300 17.600 -35.260 ;
        RECT 20.200 -35.300 20.600 -35.255 ;
        RECT 24.210 -35.260 24.440 -33.700 ;
        RECT 26.790 -35.260 27.020 -33.700 ;
        RECT 29.370 -35.260 29.600 -33.700 ;
        RECT 31.950 -35.260 32.180 -33.700 ;
        RECT 34.530 -35.260 34.760 -33.700 ;
        RECT 37.110 -35.260 37.340 -33.700 ;
        RECT 39.000 -33.870 39.300 -32.600 ;
        RECT 39.000 -34.100 39.960 -33.870 ;
        RECT 40.010 -34.500 40.240 -34.260 ;
        RECT 41.450 -34.500 41.750 -22.950 ;
        RECT 49.800 -23.600 50.300 -23.200 ;
        RECT 43.200 -24.460 48.720 -23.980 ;
        RECT 48.800 -24.460 49.440 -23.980 ;
        RECT 49.900 -24.420 50.250 -23.600 ;
        RECT 53.050 -24.380 53.400 -22.950 ;
        RECT 69.600 -23.450 70.200 -22.850 ;
        RECT 69.700 -23.850 70.100 -23.450 ;
        RECT 71.345 -23.600 73.250 -23.250 ;
        RECT 43.200 -24.500 49.440 -24.460 ;
        RECT 43.200 -25.020 43.440 -24.500 ;
        RECT 46.160 -24.960 46.400 -24.500 ;
        RECT 43.200 -27.360 43.430 -25.020 ;
        RECT 44.690 -26.820 44.920 -24.960 ;
        RECT 46.160 -25.060 46.410 -24.960 ;
        RECT 44.680 -27.540 44.920 -26.820 ;
        RECT 46.180 -27.360 46.410 -25.060 ;
        RECT 47.670 -26.860 47.900 -24.960 ;
        RECT 49.160 -25.060 49.400 -24.500 ;
        RECT 49.640 -24.740 50.480 -24.420 ;
        RECT 52.880 -24.740 53.600 -24.380 ;
        RECT 53.880 -24.500 60.320 -23.980 ;
        RECT 47.670 -27.360 47.920 -26.860 ;
        RECT 49.160 -27.360 49.390 -25.060 ;
        RECT 50.650 -26.780 50.880 -24.960 ;
        RECT 52.400 -26.740 52.630 -24.960 ;
        RECT 53.880 -25.140 54.120 -24.500 ;
        RECT 56.880 -24.960 57.120 -24.500 ;
        RECT 59.880 -24.960 60.320 -24.500 ;
        RECT 50.650 -27.360 50.920 -26.780 ;
        RECT 47.680 -27.540 47.920 -27.360 ;
        RECT 50.680 -27.540 50.920 -27.360 ;
        RECT 44.680 -27.740 50.920 -27.540 ;
        RECT 52.400 -27.540 52.640 -26.740 ;
        RECT 53.890 -27.360 54.120 -25.140 ;
        RECT 55.380 -26.740 55.610 -24.960 ;
        RECT 55.360 -27.360 55.610 -26.740 ;
        RECT 56.870 -25.140 57.120 -24.960 ;
        RECT 56.870 -27.360 57.100 -25.140 ;
        RECT 58.360 -26.740 58.590 -24.960 ;
        RECT 55.360 -27.540 55.600 -27.360 ;
        RECT 58.360 -27.540 58.600 -26.740 ;
        RECT 59.850 -27.360 60.320 -24.960 ;
        RECT 63.050 -24.460 68.570 -23.980 ;
        RECT 68.650 -24.460 69.290 -23.980 ;
        RECT 69.750 -24.420 70.100 -23.850 ;
        RECT 72.900 -24.380 73.250 -23.600 ;
        RECT 63.050 -24.500 69.290 -24.460 ;
        RECT 63.050 -25.020 63.290 -24.500 ;
        RECT 66.010 -24.960 66.250 -24.500 ;
        RECT 63.050 -27.360 63.280 -25.020 ;
        RECT 64.540 -26.820 64.770 -24.960 ;
        RECT 66.010 -25.060 66.260 -24.960 ;
        RECT 52.400 -27.740 58.600 -27.540 ;
        RECT 43.280 -28.800 43.510 -28.790 ;
        RECT 43.200 -30.500 43.510 -28.800 ;
        RECT 45.860 -30.300 46.090 -28.790 ;
        RECT 49.600 -28.850 49.880 -27.740 ;
        RECT 49.600 -29.050 49.890 -28.850 ;
        RECT 48.400 -29.500 49.890 -29.050 ;
        RECT 49.660 -29.850 49.890 -29.500 ;
        RECT 53.440 -29.980 53.680 -27.740 ;
        RECT 59.880 -28.100 60.320 -27.360 ;
        RECT 64.530 -27.540 64.770 -26.820 ;
        RECT 66.030 -27.360 66.260 -25.060 ;
        RECT 67.520 -26.860 67.750 -24.960 ;
        RECT 69.010 -25.060 69.250 -24.500 ;
        RECT 69.490 -24.740 70.330 -24.420 ;
        RECT 72.730 -24.740 73.450 -24.380 ;
        RECT 73.730 -24.500 80.170 -23.980 ;
        RECT 67.520 -27.360 67.770 -26.860 ;
        RECT 69.010 -27.360 69.240 -25.060 ;
        RECT 70.500 -26.780 70.730 -24.960 ;
        RECT 72.250 -26.740 72.480 -24.960 ;
        RECT 73.730 -25.140 73.970 -24.500 ;
        RECT 76.730 -24.960 76.970 -24.500 ;
        RECT 79.730 -24.960 80.170 -24.500 ;
        RECT 70.500 -27.360 70.770 -26.780 ;
        RECT 67.530 -27.540 67.770 -27.360 ;
        RECT 70.530 -27.540 70.770 -27.360 ;
        RECT 64.530 -27.740 70.770 -27.540 ;
        RECT 72.250 -27.540 72.490 -26.740 ;
        RECT 73.740 -27.360 73.970 -25.140 ;
        RECT 75.230 -26.740 75.460 -24.960 ;
        RECT 75.210 -27.360 75.460 -26.740 ;
        RECT 76.720 -25.140 76.970 -24.960 ;
        RECT 76.720 -27.360 76.950 -25.140 ;
        RECT 78.210 -26.740 78.440 -24.960 ;
        RECT 75.210 -27.540 75.450 -27.360 ;
        RECT 78.210 -27.540 78.450 -26.740 ;
        RECT 79.700 -27.360 80.170 -24.960 ;
        RECT 72.250 -27.740 78.450 -27.540 ;
        RECT 57.240 -28.620 60.320 -28.100 ;
        RECT 56.850 -28.820 57.080 -28.800 ;
        RECT 57.240 -28.820 57.760 -28.620 ;
        RECT 63.130 -28.800 63.360 -28.790 ;
        RECT 56.850 -29.660 57.760 -28.820 ;
        RECT 59.850 -29.220 60.080 -28.800 ;
        RECT 56.850 -29.800 57.080 -29.660 ;
        RECT 53.240 -30.010 53.680 -29.980 ;
        RECT 55.840 -30.000 58.200 -29.980 ;
        RECT 49.940 -30.020 50.400 -30.010 ;
        RECT 52.940 -30.020 53.680 -30.010 ;
        RECT 49.920 -30.220 53.680 -30.020 ;
        RECT 54.700 -30.180 58.200 -30.000 ;
        RECT 49.940 -30.240 50.400 -30.220 ;
        RECT 52.940 -30.240 53.400 -30.220 ;
        RECT 54.700 -30.235 56.800 -30.180 ;
        RECT 54.700 -30.250 56.300 -30.235 ;
        RECT 43.200 -31.100 43.500 -30.500 ;
        RECT 45.800 -31.100 46.200 -30.300 ;
        RECT 54.700 -30.700 54.900 -30.250 ;
        RECT 46.600 -30.900 54.900 -30.700 ;
        RECT 46.600 -31.000 47.500 -30.900 ;
        RECT 57.960 -30.980 58.200 -30.180 ;
        RECT 59.850 -30.460 60.800 -29.220 ;
        RECT 59.850 -30.800 60.080 -30.460 ;
        RECT 59.880 -30.980 60.040 -30.800 ;
        RECT 43.200 -31.150 46.200 -31.100 ;
        RECT 42.550 -31.400 46.200 -31.150 ;
        RECT 57.960 -31.260 60.040 -30.980 ;
        RECT 42.550 -31.900 43.650 -31.400 ;
        RECT 45.200 -31.700 45.600 -31.400 ;
        RECT 45.200 -32.000 55.800 -31.700 ;
        RECT 60.250 -31.950 60.650 -30.460 ;
        RECT 63.050 -30.500 63.360 -28.800 ;
        RECT 65.710 -30.300 65.940 -28.790 ;
        RECT 69.450 -28.850 69.730 -27.740 ;
        RECT 69.450 -29.050 69.740 -28.850 ;
        RECT 68.250 -29.500 69.740 -29.050 ;
        RECT 69.510 -29.850 69.740 -29.500 ;
        RECT 73.290 -29.980 73.530 -27.740 ;
        RECT 79.730 -28.100 80.170 -27.360 ;
        RECT 77.090 -28.620 80.170 -28.100 ;
        RECT 76.700 -28.820 76.930 -28.800 ;
        RECT 77.090 -28.820 77.610 -28.620 ;
        RECT 76.700 -29.660 77.610 -28.820 ;
        RECT 79.700 -29.220 79.930 -28.800 ;
        RECT 76.700 -29.800 76.930 -29.660 ;
        RECT 79.700 -29.825 80.650 -29.220 ;
        RECT 73.090 -30.010 73.530 -29.980 ;
        RECT 75.690 -30.000 78.050 -29.980 ;
        RECT 69.790 -30.020 70.250 -30.010 ;
        RECT 72.790 -30.020 73.530 -30.010 ;
        RECT 69.770 -30.220 73.530 -30.020 ;
        RECT 74.550 -30.180 78.050 -30.000 ;
        RECT 69.790 -30.240 70.250 -30.220 ;
        RECT 72.790 -30.240 73.250 -30.220 ;
        RECT 74.550 -30.235 76.650 -30.180 ;
        RECT 74.550 -30.250 76.150 -30.235 ;
        RECT 63.050 -31.100 63.350 -30.500 ;
        RECT 65.650 -31.100 66.050 -30.300 ;
        RECT 74.550 -30.700 74.750 -30.250 ;
        RECT 66.450 -30.900 74.750 -30.700 ;
        RECT 66.450 -31.000 67.350 -30.900 ;
        RECT 77.810 -30.980 78.050 -30.180 ;
        RECT 79.700 -30.460 80.675 -29.825 ;
        RECT 79.700 -30.800 79.930 -30.460 ;
        RECT 79.730 -30.980 79.890 -30.800 ;
        RECT 63.050 -31.150 66.050 -31.100 ;
        RECT 62.400 -31.400 66.050 -31.150 ;
        RECT 77.810 -31.260 79.890 -30.980 ;
        RECT 62.400 -31.900 63.500 -31.400 ;
        RECT 65.050 -31.700 65.450 -31.400 ;
        RECT 45.200 -32.710 45.450 -32.000 ;
        RECT 45.200 -33.000 45.470 -32.710 ;
        RECT 47.800 -32.950 48.050 -32.000 ;
        RECT 48.300 -32.650 48.900 -32.150 ;
        RECT 40.010 -34.800 41.750 -34.500 ;
        RECT 40.010 -35.000 41.200 -34.800 ;
        RECT 40.010 -35.260 40.240 -35.000 ;
        RECT 40.800 -36.000 41.200 -35.000 ;
        RECT 45.240 -35.210 45.470 -33.000 ;
        RECT 47.820 -35.210 48.050 -32.950 ;
        RECT 50.400 -32.950 50.650 -32.000 ;
        RECT 53.000 -32.710 53.250 -32.000 ;
        RECT 52.980 -32.950 53.250 -32.710 ;
        RECT 55.550 -32.900 55.800 -32.000 ;
        RECT 60.100 -32.200 60.800 -31.950 ;
        RECT 65.050 -32.000 75.650 -31.700 ;
        RECT 60.070 -32.900 60.830 -32.200 ;
        RECT 65.050 -32.710 65.300 -32.000 ;
        RECT 50.400 -35.210 50.630 -32.950 ;
        RECT 52.980 -35.210 53.210 -32.950 ;
        RECT 55.560 -35.210 55.790 -32.900 ;
        RECT 65.050 -33.000 65.320 -32.710 ;
        RECT 67.650 -32.950 67.900 -32.000 ;
        RECT 68.150 -32.650 68.750 -32.150 ;
        RECT 65.090 -35.210 65.320 -33.000 ;
        RECT 67.670 -35.210 67.900 -32.950 ;
        RECT 70.250 -32.950 70.500 -32.000 ;
        RECT 72.850 -32.710 73.100 -32.000 ;
        RECT 72.830 -32.950 73.100 -32.710 ;
        RECT 75.400 -32.900 75.650 -32.000 ;
        RECT 70.250 -35.210 70.480 -32.950 ;
        RECT 72.830 -35.210 73.060 -32.950 ;
        RECT 75.410 -35.210 75.640 -32.900 ;
        RECT 80.125 -33.155 80.675 -30.460 ;
        RECT 40.800 -36.400 45.400 -36.000 ;
        RECT 40.800 -36.700 41.200 -36.400 ;
        RECT 39.200 -37.600 41.200 -36.700 ;
        RECT 43.900 -36.900 44.200 -36.400 ;
        RECT 42.000 -38.100 43.000 -37.600 ;
        RECT 43.920 -37.650 44.150 -36.900 ;
        RECT 44.510 -37.400 44.740 -36.650 ;
        RECT 45.100 -36.900 45.400 -36.400 ;
        RECT 46.600 -36.400 48.300 -36.100 ;
        RECT 46.600 -36.650 46.950 -36.400 ;
        RECT 44.500 -38.100 44.800 -37.400 ;
        RECT 45.100 -37.650 45.330 -36.900 ;
        RECT 46.350 -37.650 47.000 -36.650 ;
        RECT 47.360 -37.500 47.590 -36.650 ;
        RECT 47.950 -36.800 48.300 -36.400 ;
        RECT 46.350 -37.700 46.950 -37.650 ;
        RECT 46.350 -37.900 46.750 -37.700 ;
        RECT 42.000 -38.400 44.800 -38.100 ;
        RECT 46.250 -38.400 46.750 -37.900 ;
        RECT 47.350 -38.300 47.600 -37.500 ;
        RECT 47.950 -37.650 48.180 -36.800 ;
        RECT 47.250 -38.700 47.700 -38.300 ;
        RECT 58.475 -38.875 59.025 -38.845 ;
        RECT 58.475 -39.425 61.955 -38.875 ;
        RECT 58.475 -39.455 59.025 -39.425 ;
      LAYER via ;
        RECT -37.850 32.950 -37.550 33.250 ;
        RECT -37.350 32.450 -37.050 32.750 ;
        RECT -21.505 21.795 -21.245 22.055 ;
        RECT -15.105 21.795 -14.845 22.055 ;
        RECT -8.605 21.795 -8.345 22.055 ;
        RECT -2.205 21.795 -1.945 22.055 ;
        RECT 4.295 21.795 4.555 22.055 ;
        RECT 10.695 21.795 10.955 22.055 ;
        RECT 17.195 21.795 17.455 22.055 ;
        RECT 23.595 21.795 23.855 22.055 ;
        RECT 30.095 21.795 30.355 22.055 ;
        RECT 36.495 21.795 36.755 22.055 ;
        RECT 42.995 21.795 43.255 22.055 ;
        RECT 49.395 21.795 49.655 22.055 ;
        RECT 2.700 20.050 3.000 20.350 ;
        RECT -21.505 19.220 -21.245 19.480 ;
        RECT -15.105 19.270 -14.845 19.530 ;
        RECT -8.605 19.270 -8.345 19.530 ;
        RECT -2.205 19.270 -1.945 19.530 ;
        RECT 4.295 19.270 4.555 19.530 ;
        RECT 10.695 19.270 10.955 19.530 ;
        RECT 17.195 19.270 17.455 19.530 ;
        RECT 23.595 19.270 23.855 19.530 ;
        RECT 30.095 19.270 30.355 19.530 ;
        RECT 36.495 19.270 36.755 19.530 ;
        RECT 42.995 19.270 43.255 19.530 ;
        RECT 49.395 19.270 49.655 19.530 ;
        RECT 2.700 17.300 3.000 17.600 ;
        RECT 1.200 11.450 1.600 11.850 ;
        RECT -12.700 10.300 -12.300 10.700 ;
        RECT -17.900 9.600 -17.500 10.000 ;
        RECT -1.750 9.350 -1.050 10.050 ;
        RECT 47.575 10.475 48.025 10.925 ;
        RECT 20.770 6.775 21.225 7.230 ;
        RECT 26.050 6.750 26.450 7.150 ;
        RECT -8.300 1.300 -7.900 1.700 ;
        RECT -6.600 1.500 -6.200 1.900 ;
        RECT 36.325 1.375 36.775 1.825 ;
        RECT -11.450 0.400 -10.950 0.900 ;
        RECT -13.680 -0.880 -13.160 -0.600 ;
        RECT -0.450 -0.400 0.050 0.100 ;
        RECT 3.250 -0.275 3.700 0.175 ;
        RECT 12.575 0.125 12.925 0.475 ;
        RECT -8.560 -0.880 -8.040 -0.600 ;
        RECT -8.000 -5.950 -7.650 -5.600 ;
        RECT -2.700 -8.350 -2.100 -7.750 ;
        RECT -1.500 -8.300 -1.100 -7.900 ;
        RECT -18.700 -8.950 -18.300 -8.550 ;
        RECT -8.050 -9.100 -7.550 -8.750 ;
        RECT 9.820 -0.880 10.340 -0.600 ;
        RECT 14.940 -0.880 15.460 -0.600 ;
        RECT 15.500 -5.950 15.850 -5.600 ;
        RECT 20.800 -8.350 21.400 -7.750 ;
        RECT 30.070 -0.880 30.590 -0.600 ;
        RECT 35.190 -0.880 35.710 -0.600 ;
        RECT 23.300 -6.600 23.700 -6.200 ;
        RECT 35.750 -5.950 36.100 -5.600 ;
        RECT 5.950 -9.050 6.350 -8.650 ;
        RECT 15.450 -9.100 15.950 -8.750 ;
        RECT 41.050 -8.350 41.650 -7.750 ;
        RECT 35.700 -9.100 36.200 -8.750 ;
        RECT -0.450 -19.650 0.050 -19.150 ;
        RECT 22.200 -19.650 22.700 -19.150 ;
        RECT 5.950 -20.450 6.350 -20.050 ;
        RECT 19.350 -20.450 19.750 -20.050 ;
        RECT 19.350 -23.500 19.750 -23.100 ;
        RECT 22.200 -23.950 22.700 -23.450 ;
        RECT 23.300 -24.700 23.700 -24.300 ;
        RECT 20.550 -29.450 21.200 -29.050 ;
        RECT 19.300 -30.950 19.950 -30.550 ;
        RECT 48.840 -24.380 49.360 -24.100 ;
        RECT 69.700 -23.350 70.100 -22.950 ;
        RECT 71.375 -23.600 71.725 -23.250 ;
        RECT 53.960 -24.380 54.480 -24.100 ;
        RECT 68.690 -24.380 69.210 -24.100 ;
        RECT 73.810 -24.380 74.330 -24.100 ;
        RECT 48.450 -29.450 48.800 -29.100 ;
        RECT 42.900 -31.850 43.500 -31.250 ;
        RECT 68.300 -29.450 68.650 -29.100 ;
        RECT 62.750 -31.850 63.350 -31.250 ;
        RECT 48.350 -32.600 48.850 -32.250 ;
        RECT 60.100 -32.900 60.800 -32.200 ;
        RECT 68.200 -32.600 68.700 -32.250 ;
        RECT 80.125 -33.125 80.675 -32.575 ;
        RECT 39.300 -37.500 41.100 -36.800 ;
        RECT 42.100 -38.300 42.900 -37.700 ;
        RECT 46.300 -38.350 46.700 -38.000 ;
        RECT 47.300 -38.650 47.650 -38.350 ;
        RECT 61.375 -39.425 61.925 -38.875 ;
      LAYER met2 ;
        RECT -39.080 34.150 -38.720 34.450 ;
        RECT -39.050 -15.000 -38.750 34.150 ;
        RECT -38.480 33.550 -38.120 33.850 ;
        RECT -38.450 -15.000 -38.150 33.550 ;
        RECT -37.850 -15.000 -37.550 33.280 ;
        RECT -37.350 -15.000 -37.050 32.780 ;
        RECT -21.550 21.750 -21.200 22.100 ;
        RECT -15.150 21.750 -14.800 22.100 ;
        RECT -8.650 21.750 -8.300 22.100 ;
        RECT -2.250 21.750 -1.900 22.100 ;
        RECT 4.250 21.750 4.600 22.100 ;
        RECT 10.650 21.750 11.000 22.100 ;
        RECT 17.150 21.750 17.500 22.100 ;
        RECT 23.550 21.750 23.900 22.100 ;
        RECT 30.050 21.750 30.400 22.100 ;
        RECT 36.450 21.750 36.800 22.100 ;
        RECT 42.950 21.750 43.300 22.100 ;
        RECT 49.350 21.750 49.700 22.100 ;
        RECT -21.500 19.510 -21.250 21.750 ;
        RECT -15.100 19.560 -14.850 21.750 ;
        RECT -8.600 19.560 -8.350 21.750 ;
        RECT -2.200 19.560 -1.950 21.750 ;
        RECT -21.505 19.190 -21.245 19.510 ;
        RECT -15.105 19.240 -14.845 19.560 ;
        RECT -8.605 19.240 -8.345 19.560 ;
        RECT -2.205 19.240 -1.945 19.560 ;
        RECT 2.700 17.600 3.000 20.380 ;
        RECT 4.300 19.560 4.550 21.750 ;
        RECT 4.295 19.240 4.555 19.560 ;
        RECT 10.700 19.530 10.950 21.750 ;
        RECT 17.200 19.560 17.450 21.750 ;
        RECT 23.600 19.560 23.850 21.750 ;
        RECT 30.100 19.560 30.350 21.750 ;
        RECT 10.665 19.270 10.985 19.530 ;
        RECT 17.195 19.240 17.455 19.560 ;
        RECT 23.595 19.240 23.855 19.560 ;
        RECT 30.095 19.240 30.355 19.560 ;
        RECT 36.500 19.530 36.750 21.750 ;
        RECT 43.000 19.560 43.250 21.750 ;
        RECT 49.400 19.560 49.650 21.750 ;
        RECT 36.465 19.270 36.785 19.530 ;
        RECT 42.995 19.240 43.255 19.560 ;
        RECT 49.395 19.240 49.655 19.560 ;
        RECT 2.670 17.300 3.030 17.600 ;
        RECT -12.800 10.200 -12.200 10.800 ;
        RECT -18.000 9.500 -17.400 10.100 ;
        RECT -1.900 9.200 -0.900 10.200 ;
        RECT -8.400 1.200 -7.800 1.800 ;
        RECT -6.700 1.400 -6.100 2.000 ;
        RECT -11.450 0.900 -10.950 0.930 ;
        RECT 1.150 0.900 1.650 11.900 ;
        RECT 47.575 7.600 48.025 10.955 ;
        RECT 20.700 6.700 21.300 7.300 ;
        RECT 25.950 6.650 26.550 7.250 ;
        RECT 47.575 7.025 48.000 7.600 ;
        RECT 43.325 6.575 48.000 7.025 ;
        RECT 36.200 1.300 36.850 1.900 ;
        RECT -11.450 0.400 1.650 0.900 ;
        RECT -11.450 0.370 -10.950 0.400 ;
        RECT -13.760 -0.960 -7.920 -0.480 ;
        RECT -8.050 -6.000 -7.600 -5.550 ;
        RECT -12.700 -7.700 -11.100 -7.600 ;
        RECT -7.950 -7.700 -7.650 -6.000 ;
        RECT -12.700 -8.050 -7.650 -7.700 ;
        RECT -12.700 -8.100 -10.800 -8.050 ;
        RECT -18.700 -20.650 -18.300 -8.520 ;
        RECT -7.950 -8.650 -7.650 -8.050 ;
        RECT -2.850 -8.400 -1.950 -7.650 ;
        RECT -1.600 -8.400 -1.000 -7.750 ;
        RECT -8.100 -9.150 -7.500 -8.650 ;
        RECT -0.450 -19.680 0.050 0.130 ;
        RECT 3.200 -0.300 3.750 0.250 ;
        RECT 12.500 0.050 13.000 0.550 ;
        RECT 9.740 -0.960 15.580 -0.480 ;
        RECT 29.990 -0.960 35.830 -0.480 ;
        RECT 15.450 -6.000 15.900 -5.550 ;
        RECT 35.700 -6.000 36.150 -5.550 ;
        RECT 10.800 -7.700 12.400 -7.600 ;
        RECT 15.550 -7.700 15.850 -6.000 ;
        RECT 10.800 -8.050 15.850 -7.700 ;
        RECT 10.800 -8.100 12.700 -8.050 ;
        RECT 5.950 -20.480 6.350 -8.620 ;
        RECT 15.550 -8.650 15.850 -8.050 ;
        RECT 20.650 -8.400 21.550 -7.650 ;
        RECT 15.400 -9.150 16.000 -8.650 ;
        RECT 22.170 -19.650 22.730 -19.150 ;
        RECT 19.300 -20.500 19.800 -20.000 ;
        RECT -18.730 -21.050 -18.270 -20.650 ;
        RECT 19.350 -23.100 19.750 -20.500 ;
        RECT 19.320 -23.500 19.780 -23.100 ;
        RECT 22.200 -23.980 22.700 -19.650 ;
        RECT 23.300 -24.300 23.700 -6.170 ;
        RECT 31.050 -7.700 32.650 -7.600 ;
        RECT 35.800 -7.700 36.100 -6.000 ;
        RECT 31.050 -8.050 36.100 -7.700 ;
        RECT 31.050 -8.100 32.950 -8.050 ;
        RECT 35.800 -8.650 36.100 -8.050 ;
        RECT 40.900 -7.850 41.800 -7.650 ;
        RECT 43.325 -7.850 43.775 6.575 ;
        RECT 40.900 -8.300 43.775 -7.850 ;
        RECT 40.900 -8.400 41.800 -8.300 ;
        RECT 35.650 -9.150 36.250 -8.650 ;
        RECT 69.600 -23.450 70.200 -22.850 ;
        RECT 71.250 -23.800 71.850 -23.150 ;
        RECT 23.270 -24.700 23.730 -24.300 ;
        RECT 48.720 -24.460 54.560 -23.980 ;
        RECT 68.570 -24.460 74.410 -23.980 ;
        RECT 20.500 -30.000 21.250 -29.000 ;
        RECT 48.400 -29.500 48.850 -29.050 ;
        RECT 68.250 -29.500 68.700 -29.050 ;
        RECT 19.250 -31.650 20.000 -30.500 ;
        RECT 19.250 -39.850 19.950 -31.650 ;
        RECT 20.675 -38.875 21.225 -30.000 ;
        RECT 42.750 -31.900 43.650 -31.150 ;
        RECT 48.450 -31.200 48.750 -29.500 ;
        RECT 51.900 -31.200 53.500 -31.100 ;
        RECT 48.450 -31.550 53.500 -31.200 ;
        RECT 48.450 -32.150 48.750 -31.550 ;
        RECT 51.600 -31.600 53.500 -31.550 ;
        RECT 62.600 -31.900 63.500 -31.150 ;
        RECT 68.300 -31.200 68.600 -29.500 ;
        RECT 71.750 -31.200 73.350 -31.100 ;
        RECT 68.300 -31.550 73.350 -31.200 ;
        RECT 68.300 -32.150 68.600 -31.550 ;
        RECT 71.450 -31.600 73.350 -31.550 ;
        RECT 48.300 -32.650 48.900 -32.150 ;
        RECT 59.205 -34.050 59.695 -33.650 ;
        RECT 39.200 -37.600 41.200 -36.700 ;
        RECT 42.000 -38.100 43.000 -37.600 ;
        RECT 46.250 -38.100 46.750 -37.900 ;
        RECT 50.050 -38.000 50.750 -37.955 ;
        RECT 42.000 -38.400 46.750 -38.100 ;
        RECT 50.000 -38.300 50.750 -38.000 ;
        RECT 59.250 -38.300 59.650 -34.050 ;
        RECT 47.250 -38.700 59.650 -38.300 ;
        RECT 50.050 -38.745 50.750 -38.700 ;
        RECT 20.675 -38.900 49.900 -38.875 ;
        RECT 50.900 -38.900 59.055 -38.875 ;
        RECT 20.675 -39.425 59.055 -38.900 ;
        RECT 60.100 -39.850 60.800 -32.170 ;
        RECT 68.150 -32.650 68.750 -32.150 ;
        RECT 78.375 -33.125 80.705 -32.575 ;
        RECT 78.375 -36.375 78.925 -33.125 ;
        RECT 61.375 -36.925 78.925 -36.375 ;
        RECT 61.375 -39.455 61.925 -36.925 ;
        RECT 19.250 -40.550 60.800 -39.850 ;
      LAYER via2 ;
        RECT -12.700 10.300 -12.300 10.700 ;
        RECT -17.900 9.600 -17.500 10.000 ;
        RECT -1.725 9.375 -1.075 10.025 ;
        RECT -8.300 1.300 -7.900 1.700 ;
        RECT -6.600 1.500 -6.200 1.900 ;
        RECT 20.795 6.800 21.200 7.205 ;
        RECT 26.075 6.775 26.425 7.125 ;
        RECT 36.350 1.400 36.750 1.800 ;
        RECT -12.600 -8.000 -12.100 -7.600 ;
        RECT -2.700 -8.350 -2.100 -7.750 ;
        RECT -1.500 -8.300 -1.100 -7.900 ;
        RECT 3.275 -0.250 3.675 0.150 ;
        RECT 12.575 0.125 12.925 0.475 ;
        RECT 10.900 -8.000 11.400 -7.600 ;
        RECT 20.800 -8.350 21.400 -7.750 ;
        RECT 31.150 -8.000 31.650 -7.600 ;
        RECT 41.050 -8.350 41.650 -7.750 ;
        RECT 69.725 -23.325 70.075 -22.975 ;
        RECT 71.375 -23.600 71.725 -23.250 ;
        RECT 42.900 -31.850 43.500 -31.250 ;
        RECT 52.900 -31.500 53.400 -31.100 ;
        RECT 62.750 -31.850 63.350 -31.250 ;
        RECT 72.750 -31.500 73.250 -31.100 ;
        RECT 59.250 -34.050 59.650 -33.650 ;
        RECT 39.300 -37.500 41.100 -36.800 ;
        RECT 42.100 -38.300 42.900 -37.700 ;
        RECT 50.050 -38.700 50.750 -38.000 ;
      LAYER met3 ;
        RECT -12.800 10.200 -12.200 10.800 ;
        RECT -18.000 9.500 -17.400 10.100 ;
        RECT -14.600 2.500 -6.105 9.500 ;
        RECT -1.900 9.200 -0.900 10.200 ;
        RECT -8.400 1.200 -7.800 1.800 ;
        RECT -6.700 1.400 -6.100 2.000 ;
        RECT 3.100 0.650 12.100 10.145 ;
        RECT 20.700 6.700 21.300 7.300 ;
        RECT 25.950 6.650 26.550 7.250 ;
        RECT 36.200 1.300 36.850 1.900 ;
        RECT 3.200 -0.300 3.750 0.250 ;
        RECT 12.500 0.050 13.000 0.550 ;
        RECT -12.700 -8.100 -12.000 -7.500 ;
        RECT -11.550 -10.800 -4.055 -4.800 ;
        RECT -2.850 -8.400 -1.950 -7.650 ;
        RECT -1.600 -8.400 -1.000 -7.800 ;
        RECT 10.800 -8.100 11.500 -7.500 ;
        RECT 11.950 -10.800 19.445 -4.800 ;
        RECT 20.650 -8.400 21.550 -7.650 ;
        RECT 31.050 -8.100 31.750 -7.500 ;
        RECT 32.200 -10.800 39.695 -4.800 ;
        RECT 40.900 -8.400 41.800 -7.650 ;
        RECT 61.050 -23.350 70.100 -22.950 ;
        RECT 42.750 -31.900 43.650 -31.150 ;
        RECT 44.855 -34.300 52.350 -28.300 ;
        RECT 52.800 -31.600 53.500 -31.000 ;
        RECT 59.225 -33.650 59.675 -33.625 ;
        RECT 61.050 -33.650 61.450 -23.350 ;
        RECT 71.250 -23.800 71.850 -23.150 ;
        RECT 62.600 -31.900 63.500 -31.150 ;
        RECT 59.225 -34.050 61.450 -33.650 ;
        RECT 59.225 -34.075 59.675 -34.050 ;
        RECT 64.705 -34.300 72.200 -28.300 ;
        RECT 72.650 -31.600 73.350 -31.000 ;
        RECT 39.200 -37.600 41.200 -36.700 ;
        RECT 42.000 -38.000 43.000 -37.600 ;
        RECT 21.000 -38.400 43.000 -38.000 ;
        RECT 21.000 -59.000 42.495 -38.400 ;
        RECT 49.900 -38.800 50.850 -37.850 ;
      LAYER via3 ;
        RECT -12.725 10.275 -12.275 10.725 ;
        RECT -17.925 9.575 -17.475 10.025 ;
        RECT -6.525 2.640 -6.205 9.360 ;
        RECT -1.745 9.355 -1.055 10.045 ;
        RECT -8.325 1.275 -7.875 1.725 ;
        RECT -6.625 1.525 -6.175 1.925 ;
        RECT 20.775 6.780 21.220 7.225 ;
        RECT 26.055 6.755 26.445 7.145 ;
        RECT 36.330 1.380 36.770 1.820 ;
        RECT 3.240 0.750 11.960 1.070 ;
        RECT 3.255 -0.270 3.695 0.170 ;
        RECT 12.550 0.100 12.950 0.500 ;
        RECT -12.600 -8.000 -12.100 -7.600 ;
        RECT -11.450 -10.660 -11.130 -4.940 ;
        RECT -2.700 -8.350 -2.100 -7.750 ;
        RECT -1.525 -8.325 -1.075 -7.875 ;
        RECT 10.900 -8.000 11.400 -7.600 ;
        RECT 12.050 -10.660 12.370 -4.940 ;
        RECT 20.800 -8.350 21.400 -7.750 ;
        RECT 31.150 -8.000 31.650 -7.600 ;
        RECT 32.300 -10.660 32.620 -4.940 ;
        RECT 41.050 -8.350 41.650 -7.750 ;
        RECT 42.900 -31.850 43.500 -31.250 ;
        RECT 51.930 -34.160 52.250 -28.440 ;
        RECT 52.900 -31.500 53.400 -31.100 ;
        RECT 71.350 -23.625 71.750 -23.275 ;
        RECT 62.750 -31.850 63.350 -31.250 ;
        RECT 71.780 -34.160 72.100 -28.440 ;
        RECT 72.750 -31.500 73.250 -31.100 ;
        RECT 39.300 -37.500 41.100 -36.800 ;
        RECT 42.075 -58.860 42.395 -38.140 ;
        RECT 50.025 -38.725 50.775 -37.975 ;
      LAYER met4 ;
        RECT -12.730 10.700 -12.270 10.730 ;
        RECT -12.730 10.300 -6.200 10.700 ;
        RECT -12.730 10.270 -12.270 10.300 ;
        RECT -17.930 10.000 -17.470 10.030 ;
        RECT -17.930 9.600 -13.300 10.000 ;
        RECT -17.930 9.570 -17.470 9.600 ;
        RECT -13.700 8.805 -13.300 9.600 ;
        RECT -6.600 9.440 -6.200 10.300 ;
        RECT 1.920 10.620 13.175 11.075 ;
        RECT -1.750 10.040 -0.600 10.050 ;
        RECT 1.920 10.040 2.375 10.620 ;
        RECT -1.750 9.585 2.375 10.040 ;
        RECT -1.750 9.550 -0.600 9.585 ;
        RECT -13.905 3.195 -7.295 8.805 ;
        RECT -8.300 1.730 -7.900 3.195 ;
        RECT -6.605 2.560 -6.125 9.440 ;
        RECT -6.600 1.930 -6.200 2.560 ;
        RECT -8.330 1.270 -7.870 1.730 ;
        RECT -6.630 1.520 -6.170 1.930 ;
        RECT -12.700 -7.600 -12.000 -7.500 ;
        RECT -11.530 -7.600 -11.050 -4.860 ;
        RECT -12.700 -8.100 -11.050 -7.600 ;
        RECT -11.530 -10.740 -11.050 -8.100 ;
        RECT -10.360 -7.650 -4.750 -5.495 ;
        RECT -1.750 -7.100 -1.050 9.550 ;
        RECT 12.720 7.230 13.175 10.620 ;
        RECT 12.720 6.775 21.225 7.230 ;
        RECT 25.950 7.150 26.550 7.250 ;
        RECT 21.900 6.750 26.550 7.150 ;
        RECT 21.900 6.350 22.300 6.750 ;
        RECT 25.950 6.650 26.550 6.750 ;
        RECT 12.550 5.950 22.300 6.350 ;
        RECT 3.160 0.670 12.040 1.150 ;
        RECT 3.250 -0.275 3.700 0.670 ;
        RECT 12.550 0.505 12.950 5.950 ;
        RECT 36.325 1.375 42.925 1.825 ;
        RECT 12.545 0.095 12.955 0.505 ;
        RECT 12.570 -4.020 12.930 0.095 ;
        RECT 12.570 -4.380 13.630 -4.020 ;
        RECT -1.800 -7.600 -1.000 -7.100 ;
        RECT -2.800 -7.650 -1.000 -7.600 ;
        RECT -10.360 -8.450 -1.000 -7.650 ;
        RECT 10.800 -7.600 11.500 -7.500 ;
        RECT 11.970 -7.600 12.450 -4.860 ;
        RECT 13.270 -5.495 13.630 -4.380 ;
        RECT 10.800 -8.100 12.450 -7.600 ;
        RECT -10.360 -10.105 -4.750 -8.450 ;
        RECT -2.800 -8.500 -1.000 -8.450 ;
        RECT 11.970 -10.740 12.450 -8.100 ;
        RECT 13.140 -7.650 18.750 -5.495 ;
        RECT 31.050 -7.600 31.750 -7.500 ;
        RECT 32.220 -7.600 32.700 -4.860 ;
        RECT 13.140 -8.450 21.650 -7.650 ;
        RECT 31.050 -8.100 32.700 -7.600 ;
        RECT 13.140 -10.105 18.750 -8.450 ;
        RECT 32.220 -10.740 32.700 -8.100 ;
        RECT 33.390 -7.650 39.000 -5.495 ;
        RECT 33.390 -8.450 41.900 -7.650 ;
        RECT 33.390 -10.105 39.000 -8.450 ;
        RECT 42.475 -12.025 42.925 1.375 ;
        RECT 42.100 -12.475 42.925 -12.025 ;
        RECT 42.100 -31.150 42.550 -12.475 ;
        RECT 71.345 -23.630 71.755 -23.270 ;
        RECT 71.375 -27.625 71.725 -23.630 ;
        RECT 69.975 -27.975 71.725 -27.625 ;
        RECT 45.550 -31.150 51.160 -28.995 ;
        RECT 42.100 -31.950 51.160 -31.150 ;
        RECT 42.100 -32.400 42.700 -31.950 ;
        RECT 39.200 -37.600 41.200 -36.700 ;
        RECT 39.200 -38.695 39.700 -37.600 ;
        RECT 42.100 -38.060 42.600 -32.400 ;
        RECT 45.550 -33.605 51.160 -31.950 ;
        RECT 51.850 -31.100 52.330 -28.360 ;
        RECT 69.975 -28.995 70.325 -27.975 ;
        RECT 52.800 -31.100 53.500 -31.000 ;
        RECT 51.850 -31.600 53.500 -31.100 ;
        RECT 65.400 -31.150 71.010 -28.995 ;
        RECT 51.850 -34.240 52.330 -31.600 ;
        RECT 62.500 -31.950 71.010 -31.150 ;
        RECT 65.400 -33.605 71.010 -31.950 ;
        RECT 71.700 -31.100 72.180 -28.360 ;
        RECT 72.650 -31.100 73.350 -31.000 ;
        RECT 71.700 -31.600 73.350 -31.100 ;
        RECT 71.700 -34.240 72.180 -31.600 ;
        RECT 21.695 -58.305 41.305 -38.695 ;
        RECT 41.995 -38.700 42.600 -38.060 ;
        RECT 41.995 -58.940 42.475 -38.700 ;
        RECT 49.900 -38.800 50.850 -37.850 ;
        RECT 50.050 -43.795 50.750 -38.800 ;
        RECT 49.645 -51.405 57.255 -43.795 ;
  END
END SystemLevel
END LIBRARY

