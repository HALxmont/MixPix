magic
tech sky130B
magscale 1 2
timestamp 1668274092
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 404998 700408 405004 700460
rect 405056 700448 405062 700460
rect 413646 700448 413652 700460
rect 405056 700420 413652 700448
rect 405056 700408 405062 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 364978 700340 364984 700392
rect 365036 700380 365042 700392
rect 397546 700380 397552 700392
rect 365036 700352 397552 700380
rect 365036 700340 365042 700352
rect 397546 700340 397552 700352
rect 397604 700340 397610 700392
rect 403618 700340 403624 700392
rect 403676 700380 403682 700392
rect 478506 700380 478512 700392
rect 403676 700352 478512 700380
rect 403676 700340 403682 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 292574 700272 292580 700324
rect 292632 700312 292638 700324
rect 300118 700312 300124 700324
rect 292632 700284 300124 700312
rect 292632 700272 292638 700284
rect 300118 700272 300124 700284
rect 300176 700272 300182 700324
rect 348786 700272 348792 700324
rect 348844 700312 348850 700324
rect 396626 700312 396632 700324
rect 348844 700284 396632 700312
rect 348844 700272 348850 700284
rect 396626 700272 396632 700284
rect 396684 700272 396690 700324
rect 400858 700272 400864 700324
rect 400916 700312 400922 700324
rect 543458 700312 543464 700324
rect 400916 700284 543464 700312
rect 400916 700272 400922 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 233878 697552 233884 697604
rect 233936 697592 233942 697604
rect 235166 697592 235172 697604
rect 233936 697564 235172 697592
rect 233936 697552 233942 697564
rect 235166 697552 235172 697564
rect 235224 697552 235230 697604
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 284938 697552 284944 697604
rect 284996 697592 285002 697604
rect 292574 697592 292580 697604
rect 284996 697564 292580 697592
rect 284996 697552 285002 697564
rect 292574 697552 292580 697564
rect 292632 697552 292638 697604
rect 182174 694764 182180 694816
rect 182232 694804 182238 694816
rect 201494 694804 201500 694816
rect 182232 694776 201500 694804
rect 182232 694764 182238 694776
rect 201494 694764 201500 694776
rect 201552 694764 201558 694816
rect 160738 692044 160744 692096
rect 160796 692084 160802 692096
rect 169662 692084 169668 692096
rect 160796 692056 169668 692084
rect 160796 692044 160802 692056
rect 169662 692044 169668 692056
rect 169720 692044 169726 692096
rect 180058 690208 180064 690260
rect 180116 690248 180122 690260
rect 182174 690248 182180 690260
rect 180116 690220 182180 690248
rect 180116 690208 180122 690220
rect 182174 690208 182180 690220
rect 182232 690208 182238 690260
rect 279418 687488 279424 687540
rect 279476 687528 279482 687540
rect 284938 687528 284944 687540
rect 279476 687500 284944 687528
rect 279476 687488 279482 687500
rect 284938 687488 284944 687500
rect 284996 687488 285002 687540
rect 233878 684536 233884 684548
rect 231872 684508 233884 684536
rect 230842 684428 230848 684480
rect 230900 684468 230906 684480
rect 231872 684468 231900 684508
rect 233878 684496 233884 684508
rect 233936 684496 233942 684548
rect 230900 684440 231900 684468
rect 230900 684428 230906 684440
rect 2774 683680 2780 683732
rect 2832 683720 2838 683732
rect 4798 683720 4804 683732
rect 2832 683692 4804 683720
rect 2832 683680 2838 683692
rect 4798 683680 4804 683692
rect 4856 683680 4862 683732
rect 399478 683136 399484 683188
rect 399536 683176 399542 683188
rect 580166 683176 580172 683188
rect 399536 683148 580172 683176
rect 399536 683136 399542 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 229738 681708 229744 681760
rect 229796 681748 229802 681760
rect 230842 681748 230848 681760
rect 229796 681720 230848 681748
rect 229796 681708 229802 681720
rect 230842 681708 230848 681720
rect 230900 681708 230906 681760
rect 147766 678036 147772 678088
rect 147824 678076 147830 678088
rect 153194 678076 153200 678088
rect 147824 678048 153200 678076
rect 147824 678036 147830 678048
rect 153194 678036 153200 678048
rect 153252 678036 153258 678088
rect 147030 675520 147036 675572
rect 147088 675560 147094 675572
rect 147766 675560 147772 675572
rect 147088 675532 147772 675560
rect 147088 675520 147094 675532
rect 147766 675520 147772 675532
rect 147824 675520 147830 675572
rect 272518 674840 272524 674892
rect 272576 674880 272582 674892
rect 279418 674880 279424 674892
rect 272576 674852 279424 674880
rect 272576 674840 272582 674852
rect 279418 674840 279424 674852
rect 279476 674840 279482 674892
rect 159450 674772 159456 674824
rect 159508 674812 159514 674824
rect 160738 674812 160744 674824
rect 159508 674784 160744 674812
rect 159508 674772 159514 674784
rect 160738 674772 160744 674784
rect 160796 674772 160802 674824
rect 266354 674092 266360 674144
rect 266412 674132 266418 674144
rect 275278 674132 275284 674144
rect 266412 674104 275284 674132
rect 266412 674092 266418 674104
rect 275278 674092 275284 674104
rect 275336 674092 275342 674144
rect 413278 670692 413284 670744
rect 413336 670732 413342 670744
rect 580166 670732 580172 670744
rect 413336 670704 580172 670732
rect 413336 670692 413342 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 157334 668584 157340 668636
rect 157392 668624 157398 668636
rect 159450 668624 159456 668636
rect 157392 668596 159456 668624
rect 157392 668584 157398 668596
rect 159450 668584 159456 668596
rect 159508 668584 159514 668636
rect 145558 667836 145564 667888
rect 145616 667876 145622 667888
rect 147030 667876 147036 667888
rect 145616 667848 147036 667876
rect 145616 667836 145622 667848
rect 147030 667836 147036 667848
rect 147088 667836 147094 667888
rect 150434 665796 150440 665848
rect 150492 665836 150498 665848
rect 157334 665836 157340 665848
rect 150492 665808 157340 665836
rect 150492 665796 150498 665808
rect 157334 665796 157340 665808
rect 157392 665796 157398 665848
rect 228358 663756 228364 663808
rect 228416 663796 228422 663808
rect 229738 663796 229744 663808
rect 228416 663768 229744 663796
rect 228416 663756 228422 663768
rect 229738 663756 229744 663768
rect 229796 663756 229802 663808
rect 146938 662396 146944 662448
rect 146996 662436 147002 662448
rect 150434 662436 150440 662448
rect 146996 662408 150440 662436
rect 146996 662396 147002 662408
rect 150434 662396 150440 662408
rect 150492 662396 150498 662448
rect 173158 662396 173164 662448
rect 173216 662436 173222 662448
rect 180058 662436 180064 662448
rect 173216 662408 180064 662436
rect 173216 662396 173222 662408
rect 180058 662396 180064 662408
rect 180116 662396 180122 662448
rect 275278 661852 275284 661904
rect 275336 661892 275342 661904
rect 278038 661892 278044 661904
rect 275336 661864 278044 661892
rect 275336 661852 275342 661864
rect 278038 661852 278044 661864
rect 278096 661852 278102 661904
rect 260098 658928 260104 658980
rect 260156 658968 260162 658980
rect 272518 658968 272524 658980
rect 260156 658940 272524 658968
rect 260156 658928 260162 658940
rect 272518 658928 272524 658940
rect 272576 658928 272582 658980
rect 215938 658180 215944 658232
rect 215996 658220 216002 658232
rect 218054 658220 218060 658232
rect 215996 658192 218060 658220
rect 215996 658180 216002 658192
rect 218054 658180 218060 658192
rect 218112 658180 218118 658232
rect 142798 657976 142804 658028
rect 142856 658016 142862 658028
rect 145558 658016 145564 658028
rect 142856 657988 145564 658016
rect 142856 657976 142862 657988
rect 145558 657976 145564 657988
rect 145616 657976 145622 658028
rect 331214 655732 331220 655784
rect 331272 655772 331278 655784
rect 335354 655772 335360 655784
rect 331272 655744 335360 655772
rect 331272 655732 331278 655744
rect 335354 655732 335360 655744
rect 335412 655732 335418 655784
rect 282914 653692 282920 653744
rect 282972 653732 282978 653744
rect 286318 653732 286324 653744
rect 282972 653704 286324 653732
rect 282972 653692 282978 653704
rect 286318 653692 286324 653704
rect 286376 653692 286382 653744
rect 142798 652780 142804 652792
rect 139412 652752 142804 652780
rect 138382 652672 138388 652724
rect 138440 652712 138446 652724
rect 139412 652712 139440 652752
rect 142798 652740 142804 652752
rect 142856 652740 142862 652792
rect 166994 652740 167000 652792
rect 167052 652780 167058 652792
rect 173158 652780 173164 652792
rect 167052 652752 173164 652780
rect 167052 652740 167058 652752
rect 173158 652740 173164 652752
rect 173216 652740 173222 652792
rect 222838 652740 222844 652792
rect 222896 652780 222902 652792
rect 228358 652780 228364 652792
rect 222896 652752 228364 652780
rect 222896 652740 222902 652752
rect 228358 652740 228364 652752
rect 228416 652740 228422 652792
rect 335354 652740 335360 652792
rect 335412 652780 335418 652792
rect 341518 652780 341524 652792
rect 335412 652752 341524 652780
rect 335412 652740 335418 652752
rect 341518 652740 341524 652752
rect 341576 652740 341582 652792
rect 138440 652684 139440 652712
rect 138440 652672 138446 652684
rect 278038 652060 278044 652112
rect 278096 652100 278102 652112
rect 281442 652100 281448 652112
rect 278096 652072 281448 652100
rect 278096 652060 278102 652072
rect 281442 652060 281448 652072
rect 281500 652060 281506 652112
rect 165338 650020 165344 650072
rect 165396 650060 165402 650072
rect 166994 650060 167000 650072
rect 165396 650032 167000 650060
rect 165396 650020 165402 650032
rect 166994 650020 167000 650032
rect 167052 650020 167058 650072
rect 213178 650020 213184 650072
rect 213236 650060 213242 650072
rect 215938 650060 215944 650072
rect 213236 650032 215944 650060
rect 213236 650020 213242 650032
rect 215938 650020 215944 650032
rect 215996 650020 216002 650072
rect 281442 647164 281448 647216
rect 281500 647204 281506 647216
rect 285674 647204 285680 647216
rect 281500 647176 285680 647204
rect 281500 647164 281506 647176
rect 285674 647164 285680 647176
rect 285732 647164 285738 647216
rect 159358 646484 159364 646536
rect 159416 646524 159422 646536
rect 165338 646524 165344 646536
rect 159416 646496 165344 646524
rect 159416 646484 159422 646496
rect 165338 646484 165344 646496
rect 165396 646484 165402 646536
rect 138382 644484 138388 644496
rect 136652 644456 138388 644484
rect 135898 644376 135904 644428
rect 135956 644416 135962 644428
rect 136652 644416 136680 644456
rect 138382 644444 138388 644456
rect 138440 644444 138446 644496
rect 135956 644388 136680 644416
rect 135956 644376 135962 644388
rect 285674 642404 285680 642456
rect 285732 642444 285738 642456
rect 289078 642444 289084 642456
rect 285732 642416 289084 642444
rect 285732 642404 285738 642416
rect 289078 642404 289084 642416
rect 289136 642404 289142 642456
rect 286318 642336 286324 642388
rect 286376 642376 286382 642388
rect 294598 642376 294604 642388
rect 286376 642348 294604 642376
rect 286376 642336 286382 642348
rect 294598 642336 294604 642348
rect 294656 642336 294662 642388
rect 221550 640296 221556 640348
rect 221608 640336 221614 640348
rect 222838 640336 222844 640348
rect 221608 640308 222844 640336
rect 221608 640296 221614 640308
rect 222838 640296 222844 640308
rect 222896 640296 222902 640348
rect 133138 639548 133144 639600
rect 133196 639588 133202 639600
rect 159358 639588 159364 639600
rect 133196 639560 159364 639588
rect 133196 639548 133202 639560
rect 159358 639548 159364 639560
rect 159416 639548 159422 639600
rect 210418 638596 210424 638648
rect 210476 638636 210482 638648
rect 213178 638636 213184 638648
rect 210476 638608 213184 638636
rect 210476 638596 210482 638608
rect 213178 638596 213184 638608
rect 213236 638596 213242 638648
rect 220078 638392 220084 638444
rect 220136 638432 220142 638444
rect 221550 638432 221556 638444
rect 220136 638404 221556 638432
rect 220136 638392 220142 638404
rect 221550 638392 221556 638404
rect 221608 638392 221614 638444
rect 3326 632068 3332 632120
rect 3384 632108 3390 632120
rect 7558 632108 7564 632120
rect 3384 632080 7564 632108
rect 3384 632068 3390 632080
rect 7558 632068 7564 632080
rect 7616 632068 7622 632120
rect 133230 630640 133236 630692
rect 133288 630680 133294 630692
rect 135898 630680 135904 630692
rect 133288 630652 135904 630680
rect 133288 630640 133294 630652
rect 135898 630640 135904 630652
rect 135956 630640 135962 630692
rect 531958 630640 531964 630692
rect 532016 630680 532022 630692
rect 579982 630680 579988 630692
rect 532016 630652 579988 630680
rect 532016 630640 532022 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 289078 630164 289084 630216
rect 289136 630204 289142 630216
rect 295334 630204 295340 630216
rect 289136 630176 295340 630204
rect 289136 630164 289142 630176
rect 295334 630164 295340 630176
rect 295392 630164 295398 630216
rect 254578 626560 254584 626612
rect 254636 626600 254642 626612
rect 260098 626600 260104 626612
rect 254636 626572 260104 626600
rect 254636 626560 254642 626572
rect 260098 626560 260104 626572
rect 260156 626560 260162 626612
rect 341518 626560 341524 626612
rect 341576 626600 341582 626612
rect 347038 626600 347044 626612
rect 341576 626572 347044 626600
rect 341576 626560 341582 626572
rect 347038 626560 347044 626572
rect 347096 626560 347102 626612
rect 295334 625540 295340 625592
rect 295392 625580 295398 625592
rect 298094 625580 298100 625592
rect 295392 625552 298100 625580
rect 295392 625540 295398 625552
rect 298094 625540 298100 625552
rect 298152 625540 298158 625592
rect 129734 623772 129740 623824
rect 129792 623812 129798 623824
rect 133230 623812 133236 623824
rect 129792 623784 133236 623812
rect 129792 623772 129798 623784
rect 133230 623772 133236 623784
rect 133288 623772 133294 623824
rect 113818 623024 113824 623076
rect 113876 623064 113882 623076
rect 133138 623064 133144 623076
rect 113876 623036 133144 623064
rect 113876 623024 113882 623036
rect 133138 623024 133144 623036
rect 133196 623024 133202 623076
rect 128998 620984 129004 621036
rect 129056 621024 129062 621036
rect 129734 621024 129740 621036
rect 129056 620996 129740 621024
rect 129056 620984 129062 620996
rect 129734 620984 129740 620996
rect 129792 620984 129798 621036
rect 298094 620304 298100 620356
rect 298152 620344 298158 620356
rect 305638 620344 305644 620356
rect 298152 620316 305644 620344
rect 298152 620304 298158 620316
rect 305638 620304 305644 620316
rect 305696 620304 305702 620356
rect 145558 618876 145564 618928
rect 145616 618916 145622 618928
rect 146938 618916 146944 618928
rect 145616 618888 146944 618916
rect 145616 618876 145622 618888
rect 146938 618876 146944 618888
rect 146996 618876 147002 618928
rect 108298 611940 108304 611992
rect 108356 611980 108362 611992
rect 113818 611980 113824 611992
rect 108356 611952 113824 611980
rect 108356 611940 108362 611952
rect 113818 611940 113824 611952
rect 113876 611940 113882 611992
rect 143534 608472 143540 608524
rect 143592 608512 143598 608524
rect 145558 608512 145564 608524
rect 143592 608484 145564 608512
rect 143592 608472 143598 608484
rect 145558 608472 145564 608484
rect 145616 608472 145622 608524
rect 294598 607860 294604 607912
rect 294656 607900 294662 607912
rect 300118 607900 300124 607912
rect 294656 607872 300124 607900
rect 294656 607860 294662 607872
rect 300118 607860 300124 607872
rect 300176 607860 300182 607912
rect 305638 606432 305644 606484
rect 305696 606472 305702 606484
rect 310882 606472 310888 606484
rect 305696 606444 310888 606472
rect 305696 606432 305702 606444
rect 310882 606432 310888 606444
rect 310940 606432 310946 606484
rect 142798 604460 142804 604512
rect 142856 604500 142862 604512
rect 143534 604500 143540 604512
rect 142856 604472 143540 604500
rect 142856 604460 142862 604472
rect 143534 604460 143540 604472
rect 143592 604460 143598 604512
rect 310882 600244 310888 600296
rect 310940 600284 310946 600296
rect 315298 600284 315304 600296
rect 310940 600256 315304 600284
rect 310940 600244 310946 600256
rect 315298 600244 315304 600256
rect 315356 600244 315362 600296
rect 79318 592628 79324 592680
rect 79376 592668 79382 592680
rect 108298 592668 108304 592680
rect 79376 592640 108304 592668
rect 79376 592628 79382 592640
rect 108298 592628 108304 592640
rect 108356 592628 108362 592680
rect 347038 592560 347044 592612
rect 347096 592600 347102 592612
rect 353938 592600 353944 592612
rect 347096 592572 353944 592600
rect 347096 592560 347102 592572
rect 353938 592560 353944 592572
rect 353996 592560 354002 592612
rect 249058 587188 249064 587240
rect 249116 587228 249122 587240
rect 254578 587228 254584 587240
rect 249116 587200 254584 587228
rect 249116 587188 249122 587200
rect 254578 587188 254584 587200
rect 254636 587188 254642 587240
rect 315298 587120 315304 587172
rect 315356 587160 315362 587172
rect 319070 587160 319076 587172
rect 315356 587132 319076 587160
rect 315356 587120 315362 587132
rect 319070 587120 319076 587132
rect 319128 587120 319134 587172
rect 141418 586508 141424 586560
rect 141476 586548 141482 586560
rect 142798 586548 142804 586560
rect 141476 586520 142804 586548
rect 141476 586508 141482 586520
rect 142798 586508 142804 586520
rect 142856 586508 142862 586560
rect 319070 582972 319076 583024
rect 319128 583012 319134 583024
rect 333974 583012 333980 583024
rect 319128 582984 333980 583012
rect 319128 582972 319134 582984
rect 333974 582972 333980 582984
rect 334032 582972 334038 583024
rect 218698 580932 218704 580984
rect 218756 580972 218762 580984
rect 220078 580972 220084 580984
rect 218756 580944 220084 580972
rect 218756 580932 218762 580944
rect 220078 580932 220084 580944
rect 220136 580932 220142 580984
rect 3326 579776 3332 579828
rect 3384 579816 3390 579828
rect 8938 579816 8944 579828
rect 3384 579788 8944 579816
rect 3384 579776 3390 579788
rect 8938 579776 8944 579788
rect 8996 579776 9002 579828
rect 333974 577464 333980 577516
rect 334032 577504 334038 577516
rect 340138 577504 340144 577516
rect 334032 577476 340144 577504
rect 334032 577464 334038 577476
rect 340138 577464 340144 577476
rect 340196 577464 340202 577516
rect 353938 577464 353944 577516
rect 353996 577504 354002 577516
rect 360838 577504 360844 577516
rect 353996 577476 360844 577504
rect 353996 577464 354002 577476
rect 360838 577464 360844 577476
rect 360896 577464 360902 577516
rect 530578 576852 530584 576904
rect 530636 576892 530642 576904
rect 580166 576892 580172 576904
rect 530636 576864 580172 576892
rect 530636 576852 530642 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 109678 576104 109684 576156
rect 109736 576144 109742 576156
rect 141418 576144 141424 576156
rect 109736 576116 141424 576144
rect 109736 576104 109742 576116
rect 141418 576104 141424 576116
rect 141476 576104 141482 576156
rect 204898 573248 204904 573300
rect 204956 573288 204962 573300
rect 210418 573288 210424 573300
rect 204956 573260 210424 573288
rect 204956 573248 204962 573260
rect 210418 573248 210424 573260
rect 210476 573248 210482 573300
rect 300118 572908 300124 572960
rect 300176 572948 300182 572960
rect 302878 572948 302884 572960
rect 300176 572920 302884 572948
rect 300176 572908 300182 572920
rect 302878 572908 302884 572920
rect 302936 572908 302942 572960
rect 340138 569168 340144 569220
rect 340196 569208 340202 569220
rect 352558 569208 352564 569220
rect 340196 569180 352564 569208
rect 340196 569168 340202 569180
rect 352558 569168 352564 569180
rect 352616 569168 352622 569220
rect 302878 562980 302884 563032
rect 302936 563020 302942 563032
rect 307018 563020 307024 563032
rect 302936 562992 307024 563020
rect 302936 562980 302942 562992
rect 307018 562980 307024 562992
rect 307076 562980 307082 563032
rect 202138 562300 202144 562352
rect 202196 562340 202202 562352
rect 204898 562340 204904 562352
rect 202196 562312 204904 562340
rect 202196 562300 202202 562312
rect 204898 562300 204904 562312
rect 204956 562300 204962 562352
rect 108298 561008 108304 561060
rect 108356 561048 108362 561060
rect 109678 561048 109684 561060
rect 108356 561020 109684 561048
rect 108356 561008 108362 561020
rect 109678 561008 109684 561020
rect 109736 561008 109742 561060
rect 239398 560940 239404 560992
rect 239456 560980 239462 560992
rect 249058 560980 249064 560992
rect 239456 560952 249064 560980
rect 239456 560940 239462 560952
rect 249058 560940 249064 560952
rect 249116 560940 249122 560992
rect 106274 556180 106280 556232
rect 106332 556220 106338 556232
rect 108298 556220 108304 556232
rect 106332 556192 108304 556220
rect 106332 556180 106338 556192
rect 108298 556180 108304 556192
rect 108356 556180 108362 556232
rect 195974 556180 195980 556232
rect 196032 556220 196038 556232
rect 202138 556220 202144 556232
rect 196032 556192 202144 556220
rect 196032 556180 196038 556192
rect 202138 556180 202144 556192
rect 202196 556180 202202 556232
rect 104158 551488 104164 551540
rect 104216 551528 104222 551540
rect 106274 551528 106280 551540
rect 104216 551500 106280 551528
rect 104216 551488 104222 551500
rect 106274 551488 106280 551500
rect 106332 551488 106338 551540
rect 191190 550808 191196 550860
rect 191248 550848 191254 550860
rect 195974 550848 195980 550860
rect 191248 550820 195980 550848
rect 191248 550808 191254 550820
rect 195974 550808 195980 550820
rect 196032 550808 196038 550860
rect 188338 547884 188344 547936
rect 188396 547924 188402 547936
rect 191190 547924 191196 547936
rect 188396 547896 191196 547924
rect 188396 547884 188402 547896
rect 191190 547884 191196 547896
rect 191248 547884 191254 547936
rect 352558 547136 352564 547188
rect 352616 547176 352622 547188
rect 364978 547176 364984 547188
rect 352616 547148 364984 547176
rect 352616 547136 352622 547148
rect 364978 547136 364984 547148
rect 365036 547136 365042 547188
rect 217410 545096 217416 545148
rect 217468 545136 217474 545148
rect 218698 545136 218704 545148
rect 217468 545108 218704 545136
rect 217468 545096 217474 545108
rect 218698 545096 218704 545108
rect 218756 545096 218762 545148
rect 215938 542988 215944 543040
rect 215996 543028 216002 543040
rect 217410 543028 217416 543040
rect 215996 543000 217416 543028
rect 215996 542988 216002 543000
rect 217410 542988 217416 543000
rect 217468 542988 217474 543040
rect 233878 542308 233884 542360
rect 233936 542348 233942 542360
rect 239398 542348 239404 542360
rect 233936 542320 239404 542348
rect 233936 542308 233942 542320
rect 239398 542308 239404 542320
rect 239456 542308 239462 542360
rect 127618 540880 127624 540932
rect 127676 540920 127682 540932
rect 128998 540920 129004 540932
rect 127676 540892 129004 540920
rect 127676 540880 127682 540892
rect 128998 540880 129004 540892
rect 129056 540880 129062 540932
rect 214558 535440 214564 535492
rect 214616 535480 214622 535492
rect 215938 535480 215944 535492
rect 214616 535452 215944 535480
rect 214616 535440 214622 535452
rect 215938 535440 215944 535452
rect 215996 535440 216002 535492
rect 307018 534692 307024 534744
rect 307076 534732 307082 534744
rect 344278 534732 344284 534744
rect 307076 534704 344284 534732
rect 307076 534692 307082 534704
rect 344278 534692 344284 534704
rect 344336 534692 344342 534744
rect 126238 529864 126244 529916
rect 126296 529904 126302 529916
rect 127618 529904 127624 529916
rect 126296 529876 127624 529904
rect 126296 529864 126302 529876
rect 127618 529864 127624 529876
rect 127676 529864 127682 529916
rect 360838 528572 360844 528624
rect 360896 528612 360902 528624
rect 366358 528612 366364 528624
rect 360896 528584 366364 528612
rect 360896 528572 360902 528584
rect 366358 528572 366364 528584
rect 366416 528572 366422 528624
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 10318 527184 10324 527196
rect 3016 527156 10324 527184
rect 3016 527144 3022 527156
rect 10318 527144 10324 527156
rect 10376 527144 10382 527196
rect 101398 527144 101404 527196
rect 101456 527184 101462 527196
rect 104158 527184 104164 527196
rect 101456 527156 104164 527184
rect 101456 527144 101462 527156
rect 104158 527144 104164 527156
rect 104216 527144 104222 527196
rect 526438 524424 526444 524476
rect 526496 524464 526502 524476
rect 580166 524464 580172 524476
rect 526496 524436 580172 524464
rect 526496 524424 526502 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 185578 523472 185584 523524
rect 185636 523512 185642 523524
rect 188338 523512 188344 523524
rect 185636 523484 188344 523512
rect 185636 523472 185642 523484
rect 188338 523472 188344 523484
rect 188396 523472 188402 523524
rect 124214 520208 124220 520260
rect 124272 520248 124278 520260
rect 126238 520248 126244 520260
rect 124272 520220 126244 520248
rect 124272 520208 124278 520220
rect 126238 520208 126244 520220
rect 126296 520208 126302 520260
rect 225598 519528 225604 519580
rect 225656 519568 225662 519580
rect 233878 519568 233884 519580
rect 225656 519540 233884 519568
rect 225656 519528 225662 519540
rect 233878 519528 233884 519540
rect 233936 519528 233942 519580
rect 344278 519528 344284 519580
rect 344336 519568 344342 519580
rect 349706 519568 349712 519580
rect 344336 519540 349712 519568
rect 344336 519528 344342 519540
rect 349706 519528 349712 519540
rect 349764 519528 349770 519580
rect 176654 518168 176660 518220
rect 176712 518208 176718 518220
rect 185578 518208 185584 518220
rect 176712 518180 185584 518208
rect 176712 518168 176718 518180
rect 185578 518168 185584 518180
rect 185636 518168 185642 518220
rect 98638 516128 98644 516180
rect 98696 516168 98702 516180
rect 101398 516168 101404 516180
rect 98696 516140 101404 516168
rect 98696 516128 98702 516140
rect 101398 516128 101404 516140
rect 101456 516128 101462 516180
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 25498 514808 25504 514820
rect 3384 514780 25504 514808
rect 3384 514768 3390 514780
rect 25498 514768 25504 514780
rect 25556 514768 25562 514820
rect 123478 514768 123484 514820
rect 123536 514808 123542 514820
rect 124214 514808 124220 514820
rect 123536 514780 124220 514808
rect 123536 514768 123542 514780
rect 124214 514768 124220 514780
rect 124272 514768 124278 514820
rect 349706 514700 349712 514752
rect 349764 514740 349770 514752
rect 355318 514740 355324 514752
rect 349764 514712 355324 514740
rect 349764 514700 349770 514712
rect 355318 514700 355324 514712
rect 355376 514700 355382 514752
rect 163498 514020 163504 514072
rect 163556 514060 163562 514072
rect 176654 514060 176660 514072
rect 163556 514032 176660 514060
rect 163556 514020 163562 514032
rect 176654 514020 176660 514032
rect 176712 514020 176718 514072
rect 211798 513272 211804 513324
rect 211856 513312 211862 513324
rect 214558 513312 214564 513324
rect 211856 513284 214564 513312
rect 211856 513272 211862 513284
rect 214558 513272 214564 513284
rect 214616 513272 214622 513324
rect 210418 508512 210424 508564
rect 210476 508552 210482 508564
rect 225598 508552 225604 508564
rect 210476 508524 225604 508552
rect 210476 508512 210482 508524
rect 225598 508512 225604 508524
rect 225656 508512 225662 508564
rect 157978 507832 157984 507884
rect 158036 507872 158042 507884
rect 163498 507872 163504 507884
rect 158036 507844 163504 507872
rect 158036 507832 158042 507844
rect 163498 507832 163504 507844
rect 163556 507832 163562 507884
rect 3234 500964 3240 501016
rect 3292 501004 3298 501016
rect 43438 501004 43444 501016
rect 3292 500976 43444 501004
rect 3292 500964 3298 500976
rect 43438 500964 43444 500976
rect 43496 500964 43502 501016
rect 203518 498176 203524 498228
rect 203576 498216 203582 498228
rect 210418 498216 210424 498228
rect 203576 498188 210424 498216
rect 203576 498176 203582 498188
rect 210418 498176 210424 498188
rect 210476 498176 210482 498228
rect 366358 494708 366364 494760
rect 366416 494748 366422 494760
rect 374638 494748 374644 494760
rect 366416 494720 374644 494748
rect 366416 494708 366422 494720
rect 374638 494708 374644 494720
rect 374696 494708 374702 494760
rect 73154 487772 73160 487824
rect 73212 487812 73218 487824
rect 79318 487812 79324 487824
rect 73212 487784 79324 487812
rect 73212 487772 73218 487784
rect 79318 487772 79324 487784
rect 79376 487772 79382 487824
rect 355318 485800 355324 485852
rect 355376 485840 355382 485852
rect 359826 485840 359832 485852
rect 355376 485812 359832 485840
rect 355376 485800 355382 485812
rect 359826 485800 359832 485812
rect 359884 485800 359890 485852
rect 149698 485052 149704 485104
rect 149756 485092 149762 485104
rect 157978 485092 157984 485104
rect 149756 485064 157984 485092
rect 149756 485052 149762 485064
rect 157978 485052 157984 485064
rect 158036 485052 158042 485104
rect 374638 485052 374644 485104
rect 374696 485092 374702 485104
rect 384022 485092 384028 485104
rect 374696 485064 384028 485092
rect 374696 485052 374702 485064
rect 384022 485052 384028 485064
rect 384080 485052 384086 485104
rect 65518 484372 65524 484424
rect 65576 484412 65582 484424
rect 73154 484412 73160 484424
rect 65576 484384 73160 484412
rect 65576 484372 65582 484384
rect 73154 484372 73160 484384
rect 73212 484372 73218 484424
rect 384022 480904 384028 480956
rect 384080 480944 384086 480956
rect 393958 480944 393964 480956
rect 384080 480916 393964 480944
rect 384080 480904 384086 480916
rect 393958 480904 393964 480916
rect 394016 480904 394022 480956
rect 359826 480700 359832 480752
rect 359884 480740 359890 480752
rect 364334 480740 364340 480752
rect 359884 480712 364340 480740
rect 359884 480700 359890 480712
rect 364334 480700 364340 480712
rect 364392 480700 364398 480752
rect 364334 476076 364340 476128
rect 364392 476116 364398 476128
rect 370590 476116 370596 476128
rect 364392 476088 370596 476116
rect 364392 476076 364398 476088
rect 370590 476076 370596 476088
rect 370648 476076 370654 476128
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 18598 474756 18604 474768
rect 3108 474728 18604 474756
rect 3108 474716 3114 474728
rect 18598 474716 18604 474728
rect 18656 474716 18662 474768
rect 97258 473016 97264 473068
rect 97316 473056 97322 473068
rect 98638 473056 98644 473068
rect 97316 473028 98644 473056
rect 97316 473016 97322 473028
rect 98638 473016 98644 473028
rect 98696 473016 98702 473068
rect 525058 470568 525064 470620
rect 525116 470608 525122 470620
rect 579982 470608 579988 470620
rect 525116 470580 579988 470608
rect 525116 470568 525122 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 364978 469820 364984 469872
rect 365036 469860 365042 469872
rect 370498 469860 370504 469872
rect 365036 469832 370504 469860
rect 365036 469820 365042 469832
rect 370498 469820 370504 469832
rect 370556 469820 370562 469872
rect 95878 469208 95884 469260
rect 95936 469248 95942 469260
rect 97258 469248 97264 469260
rect 95936 469220 97264 469248
rect 95936 469208 95942 469220
rect 97258 469208 97264 469220
rect 97316 469208 97322 469260
rect 393958 469208 393964 469260
rect 394016 469248 394022 469260
rect 396534 469248 396540 469260
rect 394016 469220 396540 469248
rect 394016 469208 394022 469220
rect 396534 469208 396540 469220
rect 396592 469208 396598 469260
rect 370590 465944 370596 465996
rect 370648 465984 370654 465996
rect 373258 465984 373264 465996
rect 370648 465956 373264 465984
rect 370648 465944 370654 465956
rect 373258 465944 373264 465956
rect 373316 465944 373322 465996
rect 210418 463360 210424 463412
rect 210476 463400 210482 463412
rect 211798 463400 211804 463412
rect 210476 463372 211804 463400
rect 210476 463360 210482 463372
rect 211798 463360 211804 463372
rect 211856 463360 211862 463412
rect 3326 462340 3332 462392
rect 3384 462380 3390 462392
rect 28258 462380 28264 462392
rect 3384 462352 28264 462380
rect 3384 462340 3390 462352
rect 28258 462340 28264 462352
rect 28316 462340 28322 462392
rect 141418 461592 141424 461644
rect 141476 461632 141482 461644
rect 149698 461632 149704 461644
rect 141476 461604 149704 461632
rect 141476 461592 141482 461604
rect 149698 461592 149704 461604
rect 149756 461592 149762 461644
rect 373258 453296 373264 453348
rect 373316 453336 373322 453348
rect 393958 453336 393964 453348
rect 373316 453308 393964 453336
rect 373316 453296 373322 453308
rect 393958 453296 393964 453308
rect 394016 453296 394022 453348
rect 62114 452616 62120 452668
rect 62172 452656 62178 452668
rect 65518 452656 65524 452668
rect 62172 452628 65524 452656
rect 62172 452616 62178 452628
rect 65518 452616 65524 452628
rect 65576 452616 65582 452668
rect 49602 449148 49608 449200
rect 49660 449188 49666 449200
rect 62114 449188 62120 449200
rect 49660 449160 62120 449188
rect 49660 449148 49666 449160
rect 62114 449148 62120 449160
rect 62172 449148 62178 449200
rect 3326 448536 3332 448588
rect 3384 448576 3390 448588
rect 37918 448576 37924 448588
rect 3384 448548 37924 448576
rect 3384 448536 3390 448548
rect 37918 448536 37924 448548
rect 37976 448536 37982 448588
rect 45002 446360 45008 446412
rect 45060 446400 45066 446412
rect 49602 446400 49608 446412
rect 45060 446372 49608 446400
rect 45060 446360 45066 446372
rect 49602 446360 49608 446372
rect 49660 446360 49666 446412
rect 94498 445680 94504 445732
rect 94556 445720 94562 445732
rect 95878 445720 95884 445732
rect 94556 445692 95884 445720
rect 94556 445680 94562 445692
rect 95878 445680 95884 445692
rect 95936 445680 95942 445732
rect 208394 438880 208400 438932
rect 208452 438920 208458 438932
rect 210418 438920 210424 438932
rect 208452 438892 210424 438920
rect 208452 438880 208458 438892
rect 210418 438880 210424 438892
rect 210476 438880 210482 438932
rect 207658 435344 207664 435396
rect 207716 435384 207722 435396
rect 208394 435384 208400 435396
rect 207716 435356 208400 435384
rect 207716 435344 207722 435356
rect 208394 435344 208400 435356
rect 208452 435344 208458 435396
rect 396718 430584 396724 430636
rect 396776 430624 396782 430636
rect 580074 430624 580080 430636
rect 396776 430596 580080 430624
rect 396776 430584 396782 430596
rect 580074 430584 580080 430596
rect 580132 430584 580138 430636
rect 200666 429156 200672 429208
rect 200724 429196 200730 429208
rect 203518 429196 203524 429208
rect 200724 429168 203524 429196
rect 200724 429156 200730 429168
rect 203518 429156 203524 429168
rect 203576 429156 203582 429208
rect 370498 424328 370504 424380
rect 370556 424368 370562 424380
rect 389818 424368 389824 424380
rect 370556 424340 389824 424368
rect 370556 424328 370562 424340
rect 389818 424328 389824 424340
rect 389876 424328 389882 424380
rect 2958 422288 2964 422340
rect 3016 422328 3022 422340
rect 13078 422328 13084 422340
rect 3016 422300 13084 422328
rect 3016 422288 3022 422300
rect 13078 422288 13084 422300
rect 13136 422288 13142 422340
rect 93118 422288 93124 422340
rect 93176 422328 93182 422340
rect 94498 422328 94504 422340
rect 93176 422300 94504 422328
rect 93176 422288 93182 422300
rect 94498 422288 94504 422300
rect 94556 422288 94562 422340
rect 197998 422288 198004 422340
rect 198056 422328 198062 422340
rect 200666 422328 200672 422340
rect 198056 422300 200672 422328
rect 198056 422288 198062 422300
rect 200666 422288 200672 422300
rect 200724 422288 200730 422340
rect 122098 420180 122104 420232
rect 122156 420220 122162 420232
rect 123478 420220 123484 420232
rect 122156 420192 123484 420220
rect 122156 420180 122162 420192
rect 123478 420180 123484 420192
rect 123536 420180 123542 420232
rect 410518 418140 410524 418192
rect 410576 418180 410582 418192
rect 580074 418180 580080 418192
rect 410576 418152 580080 418180
rect 410576 418140 410582 418152
rect 580074 418140 580080 418152
rect 580132 418140 580138 418192
rect 193858 415352 193864 415404
rect 193916 415392 193922 415404
rect 197998 415392 198004 415404
rect 193916 415364 198004 415392
rect 193916 415352 193922 415364
rect 197998 415352 198004 415364
rect 198056 415352 198062 415404
rect 91094 413924 91100 413976
rect 91152 413964 91158 413976
rect 93118 413964 93124 413976
rect 91152 413936 93124 413964
rect 91152 413924 91158 413936
rect 93118 413924 93124 413936
rect 93176 413924 93182 413976
rect 3326 409844 3332 409896
rect 3384 409884 3390 409896
rect 32398 409884 32404 409896
rect 3384 409856 32404 409884
rect 3384 409844 3390 409856
rect 32398 409844 32404 409856
rect 32456 409844 32462 409896
rect 91094 408524 91100 408536
rect 88352 408496 91100 408524
rect 87690 408416 87696 408468
rect 87748 408456 87754 408468
rect 88352 408456 88380 408496
rect 91094 408484 91100 408496
rect 91152 408484 91158 408536
rect 87748 408428 88380 408456
rect 87748 408416 87754 408428
rect 87690 405736 87696 405748
rect 85592 405708 87696 405736
rect 84194 405628 84200 405680
rect 84252 405668 84258 405680
rect 85592 405668 85620 405708
rect 87690 405696 87696 405708
rect 87748 405696 87754 405748
rect 84252 405640 85620 405668
rect 84252 405628 84258 405640
rect 207658 404376 207664 404388
rect 204272 404348 207664 404376
rect 203886 404268 203892 404320
rect 203944 404308 203950 404320
rect 204272 404308 204300 404348
rect 207658 404336 207664 404348
rect 207716 404336 207722 404388
rect 417418 404336 417424 404388
rect 417476 404376 417482 404388
rect 580074 404376 580080 404388
rect 417476 404348 580080 404376
rect 417476 404336 417482 404348
rect 580074 404336 580080 404348
rect 580132 404336 580138 404388
rect 203944 404280 204300 404308
rect 203944 404268 203950 404280
rect 393958 404268 393964 404320
rect 394016 404308 394022 404320
rect 396994 404308 397000 404320
rect 394016 404280 397000 404308
rect 394016 404268 394022 404280
rect 396994 404268 397000 404280
rect 397052 404268 397058 404320
rect 131758 402228 131764 402280
rect 131816 402268 131822 402280
rect 141418 402268 141424 402280
rect 131816 402240 141424 402268
rect 131816 402228 131822 402240
rect 141418 402228 141424 402240
rect 141476 402228 141482 402280
rect 84194 401656 84200 401668
rect 84166 401616 84200 401656
rect 84252 401616 84258 401668
rect 119338 401616 119344 401668
rect 119396 401656 119402 401668
rect 122098 401656 122104 401668
rect 119396 401628 122104 401656
rect 119396 401616 119402 401628
rect 122098 401616 122104 401628
rect 122156 401616 122162 401668
rect 82446 401548 82452 401600
rect 82504 401588 82510 401600
rect 84166 401588 84194 401616
rect 82504 401560 84194 401588
rect 82504 401548 82510 401560
rect 389818 399100 389824 399152
rect 389876 399140 389882 399152
rect 392578 399140 392584 399152
rect 389876 399112 392584 399140
rect 389876 399100 389882 399112
rect 392578 399100 392584 399112
rect 392636 399100 392642 399152
rect 116578 398828 116584 398880
rect 116636 398868 116642 398880
rect 119338 398868 119344 398880
rect 116636 398840 119344 398868
rect 116636 398828 116642 398840
rect 119338 398828 119344 398840
rect 119396 398828 119402 398880
rect 201402 397672 201408 397724
rect 201460 397712 201466 397724
rect 203886 397712 203892 397724
rect 201460 397684 203892 397712
rect 201460 397672 201466 397684
rect 203886 397672 203892 397684
rect 203944 397672 203950 397724
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 39298 397508 39304 397520
rect 3384 397480 39304 397508
rect 3384 397468 3390 397480
rect 39298 397468 39304 397480
rect 39356 397468 39362 397520
rect 80698 397468 80704 397520
rect 80756 397508 80762 397520
rect 82446 397508 82452 397520
rect 80756 397480 82452 397508
rect 80756 397468 80762 397480
rect 82446 397468 82452 397480
rect 82504 397468 82510 397520
rect 69658 396720 69664 396772
rect 69716 396760 69722 396772
rect 136634 396760 136640 396772
rect 69716 396732 136640 396760
rect 69716 396720 69722 396732
rect 136634 396720 136640 396732
rect 136692 396720 136698 396772
rect 198734 393320 198740 393372
rect 198792 393360 198798 393372
rect 201402 393360 201408 393372
rect 198792 393332 201408 393360
rect 198792 393320 198798 393332
rect 201402 393320 201408 393332
rect 201460 393320 201466 393372
rect 194502 389172 194508 389224
rect 194560 389212 194566 389224
rect 198734 389212 198740 389224
rect 194560 389184 198740 389212
rect 194560 389172 194566 389184
rect 198734 389172 198740 389184
rect 198792 389172 198798 389224
rect 73798 388424 73804 388476
rect 73856 388464 73862 388476
rect 80698 388464 80704 388476
rect 73856 388436 80704 388464
rect 73856 388424 73862 388436
rect 80698 388424 80704 388436
rect 80756 388424 80762 388476
rect 68278 384956 68284 385008
rect 68336 384996 68342 385008
rect 69658 384996 69664 385008
rect 68336 384968 69664 384996
rect 68336 384956 68342 384968
rect 69658 384956 69664 384968
rect 69716 384956 69722 385008
rect 191834 384616 191840 384668
rect 191892 384656 191898 384668
rect 194502 384656 194508 384668
rect 191892 384628 194508 384656
rect 191892 384616 191898 384628
rect 194502 384616 194508 384628
rect 194560 384616 194566 384668
rect 177298 384276 177304 384328
rect 177356 384316 177362 384328
rect 193858 384316 193864 384328
rect 177356 384288 193864 384316
rect 177356 384276 177362 384288
rect 193858 384276 193864 384288
rect 193916 384276 193922 384328
rect 189718 382236 189724 382288
rect 189776 382276 189782 382288
rect 191834 382276 191840 382288
rect 189776 382248 191840 382276
rect 189776 382236 189782 382248
rect 191834 382236 191840 382248
rect 191892 382236 191898 382288
rect 396810 378156 396816 378208
rect 396868 378196 396874 378208
rect 580074 378196 580080 378208
rect 396868 378168 580080 378196
rect 396868 378156 396874 378168
rect 580074 378156 580080 378168
rect 580132 378156 580138 378208
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 14458 371260 14464 371272
rect 3384 371232 14464 371260
rect 3384 371220 3390 371232
rect 14458 371220 14464 371232
rect 14516 371220 14522 371272
rect 392578 371152 392584 371204
rect 392636 371192 392642 371204
rect 395338 371192 395344 371204
rect 392636 371164 395344 371192
rect 392636 371152 392642 371164
rect 395338 371152 395344 371164
rect 395396 371152 395402 371204
rect 114922 370744 114928 370796
rect 114980 370784 114986 370796
rect 116578 370784 116584 370796
rect 114980 370756 116584 370784
rect 114980 370744 114986 370756
rect 116578 370744 116584 370756
rect 116636 370744 116642 370796
rect 71038 369860 71044 369912
rect 71096 369900 71102 369912
rect 73798 369900 73804 369912
rect 71096 369872 73804 369900
rect 71096 369860 71102 369872
rect 73798 369860 73804 369872
rect 73856 369860 73862 369912
rect 112438 367752 112444 367804
rect 112496 367792 112502 367804
rect 114922 367792 114928 367804
rect 112496 367764 114928 367792
rect 112496 367752 112502 367764
rect 114922 367752 114928 367764
rect 114980 367752 114986 367804
rect 409138 364352 409144 364404
rect 409196 364392 409202 364404
rect 579798 364392 579804 364404
rect 409196 364364 579804 364392
rect 409196 364352 409202 364364
rect 579798 364352 579804 364364
rect 579856 364352 579862 364404
rect 69658 362924 69664 362976
rect 69716 362964 69722 362976
rect 71038 362964 71044 362976
rect 69716 362936 71044 362964
rect 69716 362924 69722 362936
rect 71038 362924 71044 362936
rect 71096 362924 71102 362976
rect 189718 362964 189724 362976
rect 187712 362936 189724 362964
rect 186314 362856 186320 362908
rect 186372 362896 186378 362908
rect 187712 362896 187740 362936
rect 189718 362924 189724 362936
rect 189776 362924 189782 362976
rect 186372 362868 187740 362896
rect 186372 362856 186378 362868
rect 186314 360244 186320 360256
rect 184952 360216 186320 360244
rect 182358 360136 182364 360188
rect 182416 360176 182422 360188
rect 184952 360176 184980 360216
rect 186314 360204 186320 360216
rect 186372 360204 186378 360256
rect 182416 360148 184980 360176
rect 182416 360136 182422 360148
rect 65426 358776 65432 358828
rect 65484 358816 65490 358828
rect 68278 358816 68284 358828
rect 65484 358788 68284 358816
rect 65484 358776 65490 358788
rect 68278 358776 68284 358788
rect 68336 358776 68342 358828
rect 64138 358096 64144 358148
rect 64196 358136 64202 358148
rect 65426 358136 65432 358148
rect 64196 358108 65432 358136
rect 64196 358096 64202 358108
rect 65426 358096 65432 358108
rect 65484 358096 65490 358148
rect 3326 357416 3332 357468
rect 3384 357456 3390 357468
rect 26878 357456 26884 357468
rect 3384 357428 26884 357456
rect 3384 357416 3390 357428
rect 26878 357416 26884 357428
rect 26936 357416 26942 357468
rect 123478 357008 123484 357060
rect 123536 357048 123542 357060
rect 131758 357048 131764 357060
rect 123536 357020 131764 357048
rect 123536 357008 123542 357020
rect 131758 357008 131764 357020
rect 131816 357008 131822 357060
rect 182358 354736 182364 354748
rect 180812 354708 182364 354736
rect 179414 354628 179420 354680
rect 179472 354668 179478 354680
rect 180812 354668 180840 354708
rect 182358 354696 182364 354708
rect 182416 354696 182422 354748
rect 179472 354640 180840 354668
rect 179472 354628 179478 354640
rect 111058 353268 111064 353320
rect 111116 353308 111122 353320
rect 112438 353308 112444 353320
rect 111116 353280 112444 353308
rect 111116 353268 111122 353280
rect 112438 353268 112444 353280
rect 112496 353268 112502 353320
rect 414658 351908 414664 351960
rect 414716 351948 414722 351960
rect 580074 351948 580080 351960
rect 414716 351920 580080 351948
rect 414716 351908 414722 351920
rect 580074 351908 580080 351920
rect 580132 351908 580138 351960
rect 179414 346440 179420 346452
rect 178052 346412 179420 346440
rect 174998 346332 175004 346384
rect 175056 346372 175062 346384
rect 178052 346372 178080 346412
rect 179414 346400 179420 346412
rect 179472 346400 179478 346452
rect 175056 346344 178080 346372
rect 175056 346332 175062 346344
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 43530 345080 43536 345092
rect 3384 345052 43536 345080
rect 3384 345040 3390 345052
rect 43530 345040 43536 345052
rect 43588 345040 43594 345092
rect 66254 343612 66260 343664
rect 66312 343652 66318 343664
rect 69658 343652 69664 343664
rect 66312 343624 69664 343652
rect 66312 343612 66318 343624
rect 69658 343612 69664 343624
rect 69716 343612 69722 343664
rect 109770 343612 109776 343664
rect 109828 343652 109834 343664
rect 111058 343652 111064 343664
rect 109828 343624 111064 343652
rect 109828 343612 109834 343624
rect 111058 343612 111064 343624
rect 111116 343612 111122 343664
rect 117958 343612 117964 343664
rect 118016 343652 118022 343664
rect 123478 343652 123484 343664
rect 118016 343624 123484 343652
rect 118016 343612 118022 343624
rect 123478 343612 123484 343624
rect 123536 343612 123542 343664
rect 108298 340008 108304 340060
rect 108356 340048 108362 340060
rect 109770 340048 109776 340060
rect 108356 340020 109776 340048
rect 108356 340008 108362 340020
rect 109770 340008 109776 340020
rect 109828 340008 109834 340060
rect 171870 339464 171876 339516
rect 171928 339504 171934 339516
rect 174998 339504 175004 339516
rect 171928 339476 175004 339504
rect 171928 339464 171934 339476
rect 174998 339464 175004 339476
rect 175056 339464 175062 339516
rect 64230 336744 64236 336796
rect 64288 336784 64294 336796
rect 66162 336784 66168 336796
rect 64288 336756 66168 336784
rect 64288 336744 64294 336756
rect 66162 336744 66168 336756
rect 66220 336744 66226 336796
rect 165430 335452 165436 335504
rect 165488 335492 165494 335504
rect 171870 335492 171876 335504
rect 165488 335464 171876 335492
rect 165488 335452 165494 335464
rect 171870 335452 171876 335464
rect 171928 335452 171934 335504
rect 162854 332596 162860 332648
rect 162912 332636 162918 332648
rect 165430 332636 165436 332648
rect 162912 332608 165436 332636
rect 162912 332596 162918 332608
rect 165430 332596 165436 332608
rect 165488 332596 165494 332648
rect 79318 331848 79324 331900
rect 79376 331888 79382 331900
rect 117958 331888 117964 331900
rect 79376 331860 117964 331888
rect 79376 331848 79382 331860
rect 117958 331848 117964 331860
rect 118016 331848 118022 331900
rect 162854 331276 162860 331288
rect 161446 331248 162860 331276
rect 157978 331168 157984 331220
rect 158036 331208 158042 331220
rect 161446 331208 161474 331248
rect 162854 331236 162860 331248
rect 162912 331236 162918 331288
rect 158036 331180 161474 331208
rect 158036 331168 158042 331180
rect 68278 320832 68284 320884
rect 68336 320872 68342 320884
rect 79318 320872 79324 320884
rect 68336 320844 79324 320872
rect 68336 320832 68342 320844
rect 79318 320832 79324 320844
rect 79376 320832 79382 320884
rect 157978 320192 157984 320204
rect 155972 320164 157984 320192
rect 154758 320084 154764 320136
rect 154816 320124 154822 320136
rect 155972 320124 156000 320164
rect 157978 320152 157984 320164
rect 158036 320152 158042 320204
rect 154816 320096 156000 320124
rect 154816 320084 154822 320096
rect 166258 319404 166264 319456
rect 166316 319444 166322 319456
rect 177298 319444 177304 319456
rect 166316 319416 177304 319444
rect 166316 319404 166322 319416
rect 177298 319404 177304 319416
rect 177356 319404 177362 319456
rect 62758 318860 62764 318912
rect 62816 318900 62822 318912
rect 64138 318900 64144 318912
rect 62816 318872 64144 318900
rect 62816 318860 62822 318872
rect 64138 318860 64144 318872
rect 64196 318860 64202 318912
rect 3142 318792 3148 318844
rect 3200 318832 3206 318844
rect 17218 318832 17224 318844
rect 3200 318804 17224 318832
rect 3200 318792 3206 318804
rect 17218 318792 17224 318804
rect 17276 318792 17282 318844
rect 153194 318384 153200 318436
rect 153252 318424 153258 318436
rect 154758 318424 154764 318436
rect 153252 318396 154764 318424
rect 153252 318384 153258 318396
rect 154758 318384 154764 318396
rect 154816 318384 154822 318436
rect 152458 314644 152464 314696
rect 152516 314684 152522 314696
rect 153194 314684 153200 314696
rect 152516 314656 153200 314684
rect 152516 314644 152522 314656
rect 153194 314644 153200 314656
rect 153252 314644 153258 314696
rect 407758 311856 407764 311908
rect 407816 311896 407822 311908
rect 580074 311896 580080 311908
rect 407816 311868 580080 311896
rect 407816 311856 407822 311868
rect 580074 311856 580080 311868
rect 580132 311856 580138 311908
rect 153838 311108 153844 311160
rect 153896 311148 153902 311160
rect 166258 311148 166264 311160
rect 153896 311120 166264 311148
rect 153896 311108 153902 311120
rect 166258 311108 166264 311120
rect 166316 311108 166322 311160
rect 102778 305600 102784 305652
rect 102836 305640 102842 305652
rect 108298 305640 108304 305652
rect 102836 305612 108304 305640
rect 102836 305600 102842 305612
rect 108298 305600 108304 305612
rect 108356 305600 108362 305652
rect 61378 303628 61384 303680
rect 61436 303668 61442 303680
rect 64230 303668 64236 303680
rect 61436 303640 64236 303668
rect 61436 303628 61442 303640
rect 64230 303628 64236 303640
rect 64288 303628 64294 303680
rect 133138 302880 133144 302932
rect 133196 302920 133202 302932
rect 153838 302920 153844 302932
rect 133196 302892 153844 302920
rect 133196 302880 133202 302892
rect 153838 302880 153844 302892
rect 153896 302880 153902 302932
rect 61470 299412 61476 299464
rect 61528 299452 61534 299464
rect 62758 299452 62764 299464
rect 61528 299424 62764 299452
rect 61528 299412 61534 299424
rect 62758 299412 62764 299424
rect 62816 299412 62822 299464
rect 400950 298120 400956 298172
rect 401008 298160 401014 298172
rect 580074 298160 580080 298172
rect 401008 298132 580080 298160
rect 401008 298120 401014 298132
rect 580074 298120 580080 298132
rect 580132 298120 580138 298172
rect 60090 297712 60096 297764
rect 60148 297752 60154 297764
rect 61378 297752 61384 297764
rect 60148 297724 61384 297752
rect 60148 297712 60154 297724
rect 61378 297712 61384 297724
rect 61436 297712 61442 297764
rect 59998 293972 60004 294024
rect 60056 294012 60062 294024
rect 61470 294012 61476 294024
rect 60056 293984 61476 294012
rect 60056 293972 60062 293984
rect 61470 293972 61476 293984
rect 61528 293972 61534 294024
rect 124490 293224 124496 293276
rect 124548 293264 124554 293276
rect 133138 293264 133144 293276
rect 124548 293236 133144 293264
rect 124548 293224 124554 293236
rect 133138 293224 133144 293236
rect 133196 293224 133202 293276
rect 65610 292544 65616 292596
rect 65668 292584 65674 292596
rect 68278 292584 68284 292596
rect 65668 292556 68284 292584
rect 65668 292544 65674 292556
rect 68278 292544 68284 292556
rect 68336 292544 68342 292596
rect 58618 290504 58624 290556
rect 58676 290544 58682 290556
rect 60090 290544 60096 290556
rect 58676 290516 60096 290544
rect 58676 290504 58682 290516
rect 60090 290504 60096 290516
rect 60148 290504 60154 290556
rect 65518 290436 65524 290488
rect 65576 290476 65582 290488
rect 104894 290476 104900 290488
rect 65576 290448 104900 290476
rect 65576 290436 65582 290448
rect 104894 290436 104900 290448
rect 104952 290436 104958 290488
rect 101398 290368 101404 290420
rect 101456 290408 101462 290420
rect 102778 290408 102784 290420
rect 101456 290380 102784 290408
rect 101456 290368 101462 290380
rect 102778 290368 102784 290380
rect 102836 290368 102842 290420
rect 122098 288396 122104 288448
rect 122156 288436 122162 288448
rect 124490 288436 124496 288448
rect 122156 288408 124496 288436
rect 122156 288396 122162 288408
rect 124490 288396 124496 288408
rect 124548 288396 124554 288448
rect 50522 286288 50528 286340
rect 50580 286328 50586 286340
rect 65610 286328 65616 286340
rect 50580 286300 65616 286328
rect 50580 286288 50586 286300
rect 65610 286288 65616 286300
rect 65668 286288 65674 286340
rect 56594 285676 56600 285728
rect 56652 285716 56658 285728
rect 58618 285716 58624 285728
rect 56652 285688 58624 285716
rect 56652 285676 56658 285688
rect 58618 285676 58624 285688
rect 58676 285676 58682 285728
rect 57974 282888 57980 282940
rect 58032 282928 58038 282940
rect 59998 282928 60004 282940
rect 58032 282900 60004 282928
rect 58032 282888 58038 282900
rect 59998 282888 60004 282900
rect 60056 282888 60062 282940
rect 55858 282072 55864 282124
rect 55916 282112 55922 282124
rect 56594 282112 56600 282124
rect 55916 282084 56600 282112
rect 55916 282072 55922 282084
rect 56594 282072 56600 282084
rect 56652 282072 56658 282124
rect 45830 279216 45836 279268
rect 45888 279256 45894 279268
rect 50522 279256 50528 279268
rect 45888 279228 50528 279256
rect 45888 279216 45894 279228
rect 50522 279216 50528 279228
rect 50580 279216 50586 279268
rect 54478 278740 54484 278792
rect 54536 278780 54542 278792
rect 57882 278780 57888 278792
rect 54536 278752 57888 278780
rect 54536 278740 54542 278752
rect 57882 278740 57888 278752
rect 57940 278740 57946 278792
rect 62758 277992 62764 278044
rect 62816 278032 62822 278044
rect 101398 278032 101404 278044
rect 62816 278004 101404 278032
rect 62816 277992 62822 278004
rect 101398 277992 101404 278004
rect 101456 277992 101462 278044
rect 118878 277584 118884 277636
rect 118936 277624 118942 277636
rect 122098 277624 122104 277636
rect 118936 277596 122104 277624
rect 118936 277584 118942 277596
rect 122098 277584 122104 277596
rect 122156 277584 122162 277636
rect 63494 276020 63500 276072
rect 63552 276060 63558 276072
rect 65518 276060 65524 276072
rect 63552 276032 65524 276060
rect 63552 276020 63558 276032
rect 65518 276020 65524 276032
rect 65576 276020 65582 276072
rect 53834 275272 53840 275324
rect 53892 275312 53898 275324
rect 55858 275312 55864 275324
rect 53892 275284 55864 275312
rect 53892 275272 53898 275284
rect 55858 275272 55864 275284
rect 55916 275272 55922 275324
rect 112438 273912 112444 273964
rect 112496 273952 112502 273964
rect 118878 273952 118884 273964
rect 112496 273924 118884 273952
rect 112496 273912 112502 273924
rect 118878 273912 118884 273924
rect 118936 273912 118942 273964
rect 50982 271872 50988 271924
rect 51040 271912 51046 271924
rect 53834 271912 53840 271924
rect 51040 271884 53840 271912
rect 51040 271872 51046 271884
rect 53834 271872 53840 271884
rect 53892 271872 53898 271924
rect 396902 271872 396908 271924
rect 396960 271912 396966 271924
rect 579798 271912 579804 271924
rect 396960 271884 579804 271912
rect 396960 271872 396966 271884
rect 579798 271872 579804 271884
rect 579856 271872 579862 271924
rect 58526 268608 58532 268660
rect 58584 268648 58590 268660
rect 63402 268648 63408 268660
rect 58584 268620 63408 268648
rect 58584 268608 58590 268620
rect 63402 268608 63408 268620
rect 63460 268608 63466 268660
rect 46934 268064 46940 268116
rect 46992 268104 46998 268116
rect 50982 268104 50988 268116
rect 46992 268076 50988 268104
rect 46992 268064 46998 268076
rect 50982 268064 50988 268076
rect 51040 268064 51046 268116
rect 3234 266364 3240 266416
rect 3292 266404 3298 266416
rect 21358 266404 21364 266416
rect 3292 266376 21364 266404
rect 3292 266364 3298 266376
rect 21358 266364 21364 266376
rect 21416 266364 21422 266416
rect 53098 266364 53104 266416
rect 53156 266404 53162 266416
rect 54478 266404 54484 266416
rect 53156 266376 54484 266404
rect 53156 266364 53162 266376
rect 54478 266364 54484 266376
rect 54536 266364 54542 266416
rect 56134 266364 56140 266416
rect 56192 266404 56198 266416
rect 58526 266404 58532 266416
rect 56192 266376 58532 266404
rect 56192 266364 56198 266376
rect 58526 266364 58532 266376
rect 58584 266364 58590 266416
rect 45186 264120 45192 264172
rect 45244 264160 45250 264172
rect 46842 264160 46848 264172
rect 45244 264132 46848 264160
rect 45244 264120 45250 264132
rect 46842 264120 46848 264132
rect 46900 264120 46906 264172
rect 151078 263236 151084 263288
rect 151136 263276 151142 263288
rect 152458 263276 152464 263288
rect 151136 263248 152464 263276
rect 151136 263236 151142 263248
rect 152458 263236 152464 263248
rect 152516 263236 152522 263288
rect 54478 262760 54484 262812
rect 54536 262800 54542 262812
rect 56134 262800 56140 262812
rect 54536 262772 56140 262800
rect 54536 262760 54542 262772
rect 56134 262760 56140 262772
rect 56192 262760 56198 262812
rect 59998 262760 60004 262812
rect 60056 262800 60062 262812
rect 62758 262800 62764 262812
rect 60056 262772 62764 262800
rect 60056 262760 60062 262772
rect 62758 262760 62764 262772
rect 62816 262760 62822 262812
rect 93118 261468 93124 261520
rect 93176 261508 93182 261520
rect 112438 261508 112444 261520
rect 93176 261480 112444 261508
rect 93176 261468 93182 261480
rect 112438 261468 112444 261480
rect 112496 261468 112502 261520
rect 406378 258068 406384 258120
rect 406436 258108 406442 258120
rect 579982 258108 579988 258120
rect 406436 258080 579988 258108
rect 406436 258068 406442 258080
rect 579982 258068 579988 258080
rect 580040 258068 580046 258120
rect 57606 255280 57612 255332
rect 57664 255320 57670 255332
rect 59998 255320 60004 255332
rect 57664 255292 60004 255320
rect 57664 255280 57670 255292
rect 59998 255280 60004 255292
rect 60056 255280 60062 255332
rect 143074 255280 143080 255332
rect 143132 255320 143138 255332
rect 151078 255320 151084 255332
rect 143132 255292 151084 255320
rect 143132 255280 143138 255292
rect 151078 255280 151084 255292
rect 151136 255280 151142 255332
rect 3326 253920 3332 253972
rect 3384 253960 3390 253972
rect 35158 253960 35164 253972
rect 3384 253932 35164 253960
rect 3384 253920 3390 253932
rect 35158 253920 35164 253932
rect 35216 253920 35222 253972
rect 49602 253920 49608 253972
rect 49660 253960 49666 253972
rect 53098 253960 53104 253972
rect 49660 253932 53104 253960
rect 49660 253920 49666 253932
rect 53098 253920 53104 253932
rect 53156 253920 53162 253972
rect 140038 252288 140044 252340
rect 140096 252328 140102 252340
rect 143074 252328 143080 252340
rect 140096 252300 143080 252328
rect 140096 252288 140102 252300
rect 143074 252288 143080 252300
rect 143132 252288 143138 252340
rect 54478 251240 54484 251252
rect 52472 251212 54484 251240
rect 50246 251132 50252 251184
rect 50304 251172 50310 251184
rect 52472 251172 52500 251212
rect 54478 251200 54484 251212
rect 54536 251200 54542 251252
rect 50304 251144 52500 251172
rect 50304 251132 50310 251144
rect 46198 249296 46204 249348
rect 46256 249336 46262 249348
rect 49602 249336 49608 249348
rect 46256 249308 49608 249336
rect 46256 249296 46262 249308
rect 49602 249296 49608 249308
rect 49660 249296 49666 249348
rect 57606 248452 57612 248464
rect 55232 248424 57612 248452
rect 51074 248344 51080 248396
rect 51132 248384 51138 248396
rect 55232 248384 55260 248424
rect 57606 248412 57612 248424
rect 57664 248412 57670 248464
rect 51132 248356 55260 248384
rect 51132 248344 51138 248356
rect 45370 244876 45376 244928
rect 45428 244916 45434 244928
rect 50982 244916 50988 244928
rect 45428 244888 50988 244916
rect 45428 244876 45434 244888
rect 50982 244876 50988 244888
rect 51040 244876 51046 244928
rect 80054 244876 80060 244928
rect 80112 244916 80118 244928
rect 93118 244916 93124 244928
rect 80112 244888 93124 244916
rect 80112 244876 80118 244888
rect 93118 244876 93124 244888
rect 93176 244876 93182 244928
rect 138014 244400 138020 244452
rect 138072 244440 138078 244452
rect 140038 244440 140044 244452
rect 138072 244412 140044 244440
rect 138072 244400 138078 244412
rect 140038 244400 140044 244412
rect 140096 244400 140102 244452
rect 399570 244264 399576 244316
rect 399628 244304 399634 244316
rect 579982 244304 579988 244316
rect 399628 244276 579988 244304
rect 399628 244264 399634 244276
rect 579982 244264 579988 244276
rect 580040 244264 580046 244316
rect 47486 243176 47492 243228
rect 47544 243216 47550 243228
rect 50246 243216 50252 243228
rect 47544 243188 50252 243216
rect 47544 243176 47550 243188
rect 50246 243176 50252 243188
rect 50304 243176 50310 243228
rect 44910 240864 44916 240916
rect 44968 240904 44974 240916
rect 71774 240904 71780 240916
rect 44968 240876 71780 240904
rect 44968 240864 44974 240876
rect 71774 240864 71780 240876
rect 71832 240864 71838 240916
rect 45278 240796 45284 240848
rect 45336 240836 45342 240848
rect 88334 240836 88340 240848
rect 45336 240808 88340 240836
rect 45336 240796 45342 240808
rect 88334 240796 88340 240808
rect 88392 240796 88398 240848
rect 45830 240728 45836 240780
rect 45888 240768 45894 240780
rect 138014 240768 138020 240780
rect 45888 240740 138020 240768
rect 45888 240728 45894 240740
rect 138014 240728 138020 240740
rect 138072 240728 138078 240780
rect 45646 240592 45652 240644
rect 45704 240632 45710 240644
rect 47486 240632 47492 240644
rect 45704 240604 47492 240632
rect 45704 240592 45710 240604
rect 47486 240592 47492 240604
rect 47544 240592 47550 240644
rect 2774 240320 2780 240372
rect 2832 240360 2838 240372
rect 4890 240360 4896 240372
rect 2832 240332 4896 240360
rect 2832 240320 2838 240332
rect 4890 240320 4896 240332
rect 4948 240320 4954 240372
rect 45462 240184 45468 240236
rect 45520 240224 45526 240236
rect 46198 240224 46204 240236
rect 45520 240196 46204 240224
rect 45520 240184 45526 240196
rect 46198 240184 46204 240196
rect 46256 240184 46262 240236
rect 395338 240048 395344 240100
rect 395396 240088 395402 240100
rect 396442 240088 396448 240100
rect 395396 240060 396448 240088
rect 395396 240048 395402 240060
rect 396442 240048 396448 240060
rect 396500 240048 396506 240100
rect 80054 239816 80060 239828
rect 64846 239788 80060 239816
rect 45554 239368 45560 239420
rect 45612 239408 45618 239420
rect 64846 239408 64874 239788
rect 80054 239776 80060 239788
rect 80112 239776 80118 239828
rect 45612 239380 64874 239408
rect 45612 239368 45618 239380
rect 44818 238824 44824 238876
rect 44876 238864 44882 238876
rect 45738 238864 45744 238876
rect 44876 238836 45744 238864
rect 44876 238824 44882 238836
rect 45738 238824 45744 238836
rect 45796 238824 45802 238876
rect 45094 238756 45100 238808
rect 45152 238796 45158 238808
rect 45830 238796 45836 238808
rect 45152 238768 45836 238796
rect 45152 238756 45158 238768
rect 45830 238756 45836 238768
rect 45888 238756 45894 238808
rect 45186 233180 45192 233232
rect 45244 233220 45250 233232
rect 45830 233220 45836 233232
rect 45244 233192 45836 233220
rect 45244 233180 45250 233192
rect 45830 233180 45836 233192
rect 45888 233180 45894 233232
rect 45462 232908 45468 232960
rect 45520 232948 45526 232960
rect 45520 232920 64874 232948
rect 45520 232908 45526 232920
rect 64846 232404 64874 232920
rect 86218 232404 86224 232416
rect 64846 232376 86224 232404
rect 86218 232364 86224 232376
rect 86276 232364 86282 232416
rect 394142 232364 394148 232416
rect 394200 232404 394206 232416
rect 396994 232404 397000 232416
rect 394200 232376 397000 232404
rect 394200 232364 394206 232376
rect 396994 232364 397000 232376
rect 397052 232364 397058 232416
rect 393958 231820 393964 231872
rect 394016 231860 394022 231872
rect 580074 231860 580080 231872
rect 394016 231832 580080 231860
rect 394016 231820 394022 231832
rect 580074 231820 580080 231832
rect 580132 231820 580138 231872
rect 3694 231140 3700 231192
rect 3752 231180 3758 231192
rect 180794 231180 180800 231192
rect 3752 231152 180800 231180
rect 3752 231140 3758 231152
rect 180794 231140 180800 231152
rect 180852 231140 180858 231192
rect 384390 231140 384396 231192
rect 384448 231180 384454 231192
rect 396442 231180 396448 231192
rect 384448 231152 396448 231180
rect 384448 231140 384454 231152
rect 396442 231140 396448 231152
rect 396500 231140 396506 231192
rect 45830 231072 45836 231124
rect 45888 231112 45894 231124
rect 49694 231112 49700 231124
rect 45888 231084 49700 231112
rect 45888 231072 45894 231084
rect 49694 231072 49700 231084
rect 49752 231072 49758 231124
rect 118602 231072 118608 231124
rect 118660 231112 118666 231124
rect 397546 231112 397552 231124
rect 118660 231084 397552 231112
rect 118660 231072 118666 231084
rect 397546 231072 397552 231084
rect 397604 231072 397610 231124
rect 45370 231004 45376 231056
rect 45428 231044 45434 231056
rect 150434 231044 150440 231056
rect 45428 231016 150440 231044
rect 45428 231004 45434 231016
rect 150434 231004 150440 231016
rect 150492 231004 150498 231056
rect 86218 230800 86224 230852
rect 86276 230840 86282 230852
rect 88886 230840 88892 230852
rect 86276 230812 88892 230840
rect 86276 230800 86282 230812
rect 88886 230800 88892 230812
rect 88944 230800 88950 230852
rect 45554 230460 45560 230512
rect 45612 230500 45618 230512
rect 45612 230472 48360 230500
rect 45612 230460 45618 230472
rect 48332 230432 48360 230472
rect 390554 230460 390560 230512
rect 390612 230500 390618 230512
rect 394142 230500 394148 230512
rect 390612 230472 394148 230500
rect 390612 230460 390618 230472
rect 394142 230460 394148 230472
rect 394200 230460 394206 230512
rect 54478 230432 54484 230444
rect 48332 230404 54484 230432
rect 54478 230392 54484 230404
rect 54536 230392 54542 230444
rect 163498 229780 163504 229832
rect 163556 229820 163562 229832
rect 176654 229820 176660 229832
rect 163556 229792 176660 229820
rect 163556 229780 163562 229792
rect 176654 229780 176660 229792
rect 176712 229780 176718 229832
rect 45094 229712 45100 229764
rect 45152 229752 45158 229764
rect 53098 229752 53104 229764
rect 45152 229724 53104 229752
rect 45152 229712 45158 229724
rect 53098 229712 53104 229724
rect 53156 229712 53162 229764
rect 120810 229712 120816 229764
rect 120868 229752 120874 229764
rect 580718 229752 580724 229764
rect 120868 229724 580724 229752
rect 120868 229712 120874 229724
rect 580718 229712 580724 229724
rect 580776 229712 580782 229764
rect 150434 229440 150440 229492
rect 150492 229480 150498 229492
rect 153194 229480 153200 229492
rect 150492 229452 153200 229480
rect 150492 229440 150498 229452
rect 153194 229440 153200 229452
rect 153252 229440 153258 229492
rect 49694 229100 49700 229152
rect 49752 229140 49758 229152
rect 49752 229112 51120 229140
rect 49752 229100 49758 229112
rect 51092 229072 51120 229112
rect 52454 229072 52460 229084
rect 51092 229044 52460 229072
rect 52454 229032 52460 229044
rect 52512 229032 52518 229084
rect 166258 228420 166264 228472
rect 166316 228460 166322 228472
rect 296714 228460 296720 228472
rect 166316 228432 296720 228460
rect 166316 228420 166322 228432
rect 296714 228420 296720 228432
rect 296772 228420 296778 228472
rect 53098 228352 53104 228404
rect 53156 228392 53162 228404
rect 58894 228392 58900 228404
rect 53156 228364 58900 228392
rect 53156 228352 53162 228364
rect 58894 228352 58900 228364
rect 58952 228352 58958 228404
rect 117222 228352 117228 228404
rect 117280 228392 117286 228404
rect 143534 228392 143540 228404
rect 117280 228364 143540 228392
rect 117280 228352 117286 228364
rect 143534 228352 143540 228364
rect 143592 228352 143598 228404
rect 161382 228352 161388 228404
rect 161440 228392 161446 228404
rect 386506 228392 386512 228404
rect 161440 228364 386512 228392
rect 161440 228352 161446 228364
rect 386506 228352 386512 228364
rect 386564 228352 386570 228404
rect 391934 228352 391940 228404
rect 391992 228392 391998 228404
rect 396534 228392 396540 228404
rect 391992 228364 396540 228392
rect 391992 228352 391998 228364
rect 396534 228352 396540 228364
rect 396592 228352 396598 228404
rect 3050 227740 3056 227792
rect 3108 227780 3114 227792
rect 140038 227780 140044 227792
rect 3108 227752 140044 227780
rect 3108 227740 3114 227752
rect 140038 227740 140044 227752
rect 140096 227740 140102 227792
rect 144914 227740 144920 227792
rect 144972 227780 144978 227792
rect 146478 227780 146484 227792
rect 144972 227752 146484 227780
rect 144972 227740 144978 227752
rect 146478 227740 146484 227752
rect 146536 227740 146542 227792
rect 44818 227196 44824 227248
rect 44876 227236 44882 227248
rect 47394 227236 47400 227248
rect 44876 227208 47400 227236
rect 44876 227196 44882 227208
rect 47394 227196 47400 227208
rect 47452 227196 47458 227248
rect 120718 226992 120724 227044
rect 120776 227032 120782 227044
rect 580166 227032 580172 227044
rect 120776 227004 580172 227032
rect 120776 226992 120782 227004
rect 580166 226992 580172 227004
rect 580224 226992 580230 227044
rect 153194 226516 153200 226568
rect 153252 226556 153258 226568
rect 155954 226556 155960 226568
rect 153252 226528 155960 226556
rect 153252 226516 153258 226528
rect 155954 226516 155960 226528
rect 156012 226516 156018 226568
rect 52454 226312 52460 226364
rect 52512 226352 52518 226364
rect 52512 226324 55214 226352
rect 52512 226312 52518 226324
rect 55186 226284 55214 226324
rect 56686 226284 56692 226296
rect 55186 226256 56692 226284
rect 56686 226244 56692 226256
rect 56744 226244 56750 226296
rect 387794 225020 387800 225072
rect 387852 225060 387858 225072
rect 390462 225060 390468 225072
rect 387852 225032 390468 225060
rect 387852 225020 387858 225032
rect 390462 225020 390468 225032
rect 390520 225020 390526 225072
rect 88886 224952 88892 225004
rect 88944 224992 88950 225004
rect 88944 224964 89760 224992
rect 88944 224952 88950 224964
rect 45002 224884 45008 224936
rect 45060 224924 45066 224936
rect 47578 224924 47584 224936
rect 45060 224896 47584 224924
rect 45060 224884 45066 224896
rect 47578 224884 47584 224896
rect 47636 224884 47642 224936
rect 89732 224924 89760 224964
rect 387058 224952 387064 225004
rect 387116 224992 387122 225004
rect 391934 224992 391940 225004
rect 387116 224964 391940 224992
rect 387116 224952 387122 224964
rect 391934 224952 391940 224964
rect 391992 224952 391998 225004
rect 91094 224924 91100 224936
rect 89732 224896 91100 224924
rect 91094 224884 91100 224896
rect 91152 224884 91158 224936
rect 58894 224204 58900 224256
rect 58952 224244 58958 224256
rect 63494 224244 63500 224256
rect 58952 224216 63500 224244
rect 58952 224204 58958 224216
rect 63494 224204 63500 224216
rect 63552 224204 63558 224256
rect 118694 224204 118700 224256
rect 118752 224244 118758 224256
rect 580810 224244 580816 224256
rect 118752 224216 580816 224244
rect 118752 224204 118758 224216
rect 580810 224204 580816 224216
rect 580868 224204 580874 224256
rect 155954 223524 155960 223576
rect 156012 223564 156018 223576
rect 157978 223564 157984 223576
rect 156012 223536 157984 223564
rect 156012 223524 156018 223536
rect 157978 223524 157984 223536
rect 158036 223524 158042 223576
rect 56686 222164 56692 222216
rect 56744 222204 56750 222216
rect 56744 222176 58020 222204
rect 56744 222164 56750 222176
rect 57992 222136 58020 222176
rect 60642 222136 60648 222148
rect 57992 222108 60648 222136
rect 60642 222096 60648 222108
rect 60700 222096 60706 222148
rect 383654 221824 383660 221876
rect 383712 221864 383718 221876
rect 387794 221864 387800 221876
rect 383712 221836 387800 221864
rect 383712 221824 383718 221836
rect 387794 221824 387800 221836
rect 387852 221824 387858 221876
rect 47394 220736 47400 220788
rect 47452 220776 47458 220788
rect 49602 220776 49608 220788
rect 47452 220748 49608 220776
rect 47452 220736 47458 220748
rect 49602 220736 49608 220748
rect 49660 220736 49666 220788
rect 63494 220124 63500 220176
rect 63552 220164 63558 220176
rect 68278 220164 68284 220176
rect 63552 220136 68284 220164
rect 63552 220124 63558 220136
rect 68278 220124 68284 220136
rect 68336 220124 68342 220176
rect 3878 220056 3884 220108
rect 3936 220096 3942 220108
rect 179506 220096 179512 220108
rect 3936 220068 179512 220096
rect 3936 220056 3942 220068
rect 179506 220056 179512 220068
rect 179564 220056 179570 220108
rect 91094 219444 91100 219496
rect 91152 219484 91158 219496
rect 91152 219456 92520 219484
rect 91152 219444 91158 219456
rect 92492 219416 92520 219456
rect 95142 219416 95148 219428
rect 92492 219388 95148 219416
rect 95142 219376 95148 219388
rect 95200 219376 95206 219428
rect 54478 218220 54484 218272
rect 54536 218260 54542 218272
rect 56686 218260 56692 218272
rect 54536 218232 56692 218260
rect 54536 218220 54542 218232
rect 56686 218220 56692 218232
rect 56744 218220 56750 218272
rect 382274 218084 382280 218136
rect 382332 218124 382338 218136
rect 383654 218124 383660 218136
rect 382332 218096 383660 218124
rect 382332 218084 382338 218096
rect 383654 218084 383660 218096
rect 383712 218084 383718 218136
rect 192478 218016 192484 218068
rect 192536 218056 192542 218068
rect 580166 218056 580172 218068
rect 192536 218028 580172 218056
rect 192536 218016 192542 218028
rect 580166 218016 580172 218028
rect 580224 218016 580230 218068
rect 60642 217744 60648 217796
rect 60700 217784 60706 217796
rect 64138 217784 64144 217796
rect 60700 217756 64144 217784
rect 60700 217744 60706 217756
rect 64138 217744 64144 217756
rect 64196 217744 64202 217796
rect 95142 216588 95148 216640
rect 95200 216628 95206 216640
rect 98086 216628 98092 216640
rect 95200 216600 98092 216628
rect 95200 216588 95206 216600
rect 98086 216588 98092 216600
rect 98144 216588 98150 216640
rect 49694 214752 49700 214804
rect 49752 214792 49758 214804
rect 53098 214792 53104 214804
rect 49752 214764 53104 214792
rect 49752 214752 49758 214764
rect 53098 214752 53104 214764
rect 53156 214752 53162 214804
rect 3326 213936 3332 213988
rect 3384 213976 3390 213988
rect 22738 213976 22744 213988
rect 3384 213948 22744 213976
rect 3384 213936 3390 213948
rect 22738 213936 22744 213948
rect 22796 213936 22802 213988
rect 98086 213868 98092 213920
rect 98144 213908 98150 213920
rect 104158 213908 104164 213920
rect 98144 213880 104164 213908
rect 98144 213868 98150 213880
rect 104158 213868 104164 213880
rect 104216 213868 104222 213920
rect 56686 212440 56692 212492
rect 56744 212480 56750 212492
rect 58710 212480 58716 212492
rect 56744 212452 58716 212480
rect 56744 212440 56750 212452
rect 58710 212440 58716 212452
rect 58768 212440 58774 212492
rect 104158 211760 104164 211812
rect 104216 211800 104222 211812
rect 108298 211800 108304 211812
rect 104216 211772 108304 211800
rect 104216 211760 104222 211772
rect 108298 211760 108304 211772
rect 108356 211760 108362 211812
rect 382274 209828 382280 209840
rect 380912 209800 382280 209828
rect 378778 209720 378784 209772
rect 378836 209760 378842 209772
rect 380912 209760 380940 209800
rect 382274 209788 382280 209800
rect 382332 209788 382338 209840
rect 378836 209732 380940 209760
rect 378836 209720 378842 209732
rect 4062 209040 4068 209092
rect 4120 209080 4126 209092
rect 180886 209080 180892 209092
rect 4120 209052 180892 209080
rect 4120 209040 4126 209052
rect 180886 209040 180892 209052
rect 180944 209040 180950 209092
rect 58710 208360 58716 208412
rect 58768 208400 58774 208412
rect 61378 208400 61384 208412
rect 58768 208372 61384 208400
rect 58768 208360 58774 208372
rect 61378 208360 61384 208372
rect 61436 208360 61442 208412
rect 157978 208360 157984 208412
rect 158036 208400 158042 208412
rect 158036 208372 161474 208400
rect 158036 208360 158042 208372
rect 161446 208332 161474 208372
rect 162118 208332 162124 208344
rect 161446 208304 162124 208332
rect 162118 208292 162124 208304
rect 162176 208292 162182 208344
rect 53098 207000 53104 207052
rect 53156 207040 53162 207052
rect 53156 207012 55214 207040
rect 53156 207000 53162 207012
rect 55186 206972 55214 207012
rect 55858 206972 55864 206984
rect 55186 206944 55864 206972
rect 55858 206932 55864 206944
rect 55916 206932 55922 206984
rect 384298 205708 384304 205760
rect 384356 205748 384362 205760
rect 387058 205748 387064 205760
rect 384356 205720 387064 205748
rect 384356 205708 384362 205720
rect 387058 205708 387064 205720
rect 387116 205708 387122 205760
rect 122098 205640 122104 205692
rect 122156 205680 122162 205692
rect 580166 205680 580172 205692
rect 122156 205652 580172 205680
rect 122156 205640 122162 205652
rect 580166 205640 580172 205652
rect 580224 205640 580230 205692
rect 45646 205164 45652 205216
rect 45704 205204 45710 205216
rect 49602 205204 49608 205216
rect 45704 205176 49608 205204
rect 45704 205164 45710 205176
rect 49602 205164 49608 205176
rect 49660 205164 49666 205216
rect 64138 204212 64144 204264
rect 64196 204252 64202 204264
rect 65518 204252 65524 204264
rect 64196 204224 65524 204252
rect 64196 204212 64202 204224
rect 65518 204212 65524 204224
rect 65576 204212 65582 204264
rect 155218 203532 155224 203584
rect 155276 203572 155282 203584
rect 266354 203572 266360 203584
rect 155276 203544 266360 203572
rect 155276 203532 155282 203544
rect 266354 203532 266360 203544
rect 266412 203532 266418 203584
rect 49602 202784 49608 202836
rect 49660 202824 49666 202836
rect 53834 202824 53840 202836
rect 49660 202796 53840 202824
rect 49660 202784 49666 202796
rect 53834 202784 53840 202796
rect 53892 202784 53898 202836
rect 153194 202104 153200 202156
rect 153252 202144 153258 202156
rect 235994 202144 236000 202156
rect 153252 202116 236000 202144
rect 153252 202104 153258 202116
rect 235994 202104 236000 202116
rect 236052 202104 236058 202156
rect 47578 201424 47584 201476
rect 47636 201464 47642 201476
rect 50338 201464 50344 201476
rect 47636 201436 50344 201464
rect 47636 201424 47642 201436
rect 50338 201424 50344 201436
rect 50396 201424 50402 201476
rect 155954 200744 155960 200796
rect 156012 200784 156018 200796
rect 166258 200784 166264 200796
rect 156012 200756 166264 200784
rect 156012 200744 156018 200756
rect 166258 200744 166264 200756
rect 166316 200744 166322 200796
rect 140038 199384 140044 199436
rect 140096 199424 140102 199436
rect 164234 199424 164240 199436
rect 140096 199396 164240 199424
rect 140096 199384 140102 199396
rect 164234 199384 164240 199396
rect 164292 199384 164298 199436
rect 148962 198024 148968 198076
rect 149020 198064 149026 198076
rect 207014 198064 207020 198076
rect 149020 198036 207020 198064
rect 149020 198024 149026 198036
rect 207014 198024 207020 198036
rect 207072 198024 207078 198076
rect 159818 197956 159824 198008
rect 159876 197996 159882 198008
rect 356054 197996 356060 198008
rect 159876 197968 356060 197996
rect 159876 197956 159882 197968
rect 356054 197956 356060 197968
rect 356112 197956 356118 198008
rect 376018 197344 376024 197396
rect 376076 197384 376082 197396
rect 378778 197384 378784 197396
rect 376076 197356 378784 197384
rect 376076 197344 376082 197356
rect 378778 197344 378784 197356
rect 378836 197344 378842 197396
rect 53834 197276 53840 197328
rect 53892 197316 53898 197328
rect 57698 197316 57704 197328
rect 53892 197288 57704 197316
rect 53892 197276 53898 197288
rect 57698 197276 57704 197288
rect 57756 197276 57762 197328
rect 65518 196664 65524 196716
rect 65576 196704 65582 196716
rect 66898 196704 66904 196716
rect 65576 196676 66904 196704
rect 65576 196664 65582 196676
rect 66898 196664 66904 196676
rect 66956 196664 66962 196716
rect 158254 196596 158260 196648
rect 158312 196636 158318 196648
rect 327074 196636 327080 196648
rect 158312 196608 327080 196636
rect 158312 196596 158318 196608
rect 327074 196596 327080 196608
rect 327132 196596 327138 196648
rect 162118 195984 162124 196036
rect 162176 196024 162182 196036
rect 162176 195996 164280 196024
rect 162176 195984 162182 195996
rect 56594 195916 56600 195968
rect 56652 195956 56658 195968
rect 138106 195956 138112 195968
rect 56652 195928 138112 195956
rect 56652 195916 56658 195928
rect 138106 195916 138112 195928
rect 138164 195916 138170 195968
rect 164252 195956 164280 195996
rect 166258 195956 166264 195968
rect 164252 195928 166264 195956
rect 166258 195916 166264 195928
rect 166316 195916 166322 195968
rect 86954 195848 86960 195900
rect 87012 195888 87018 195900
rect 139394 195888 139400 195900
rect 87012 195860 139400 195888
rect 87012 195848 87018 195860
rect 139394 195848 139400 195860
rect 139452 195848 139458 195900
rect 150342 195644 150348 195696
rect 150400 195684 150406 195696
rect 165430 195684 165436 195696
rect 150400 195656 165436 195684
rect 150400 195644 150406 195656
rect 165430 195644 165436 195656
rect 165488 195644 165494 195696
rect 379514 193740 379520 193792
rect 379572 193780 379578 193792
rect 384390 193780 384396 193792
rect 379572 193752 384396 193780
rect 379572 193740 379578 193752
rect 384390 193740 384396 193752
rect 384448 193740 384454 193792
rect 57698 193128 57704 193180
rect 57756 193168 57762 193180
rect 61746 193168 61752 193180
rect 57756 193140 61752 193168
rect 57756 193128 57762 193140
rect 61746 193128 61752 193140
rect 61804 193128 61810 193180
rect 151630 191088 151636 191140
rect 151688 191088 151694 191140
rect 371878 191088 371884 191140
rect 371936 191128 371942 191140
rect 379514 191128 379520 191140
rect 371936 191100 379520 191128
rect 371936 191088 371942 191100
rect 379514 191088 379520 191100
rect 379572 191088 379578 191140
rect 50338 190884 50344 190936
rect 50396 190924 50402 190936
rect 57238 190924 57244 190936
rect 50396 190896 57244 190924
rect 50396 190884 50402 190896
rect 57238 190884 57244 190896
rect 57296 190884 57302 190936
rect 2958 187688 2964 187740
rect 3016 187728 3022 187740
rect 119338 187728 119344 187740
rect 3016 187700 119344 187728
rect 3016 187688 3022 187700
rect 119338 187688 119344 187700
rect 119396 187688 119402 187740
rect 61746 184832 61752 184884
rect 61804 184872 61810 184884
rect 64966 184872 64972 184884
rect 61804 184844 64972 184872
rect 61804 184832 61810 184844
rect 64966 184832 64972 184844
rect 65024 184832 65030 184884
rect 68278 184832 68284 184884
rect 68336 184872 68342 184884
rect 72418 184872 72424 184884
rect 68336 184844 72424 184872
rect 68336 184832 68342 184844
rect 72418 184832 72424 184844
rect 72476 184832 72482 184884
rect 66898 183472 66904 183524
rect 66956 183512 66962 183524
rect 68278 183512 68284 183524
rect 66956 183484 68284 183512
rect 66956 183472 66962 183484
rect 68278 183472 68284 183484
rect 68336 183472 68342 183524
rect 55858 182112 55864 182164
rect 55916 182152 55922 182164
rect 58618 182152 58624 182164
rect 55916 182124 58624 182152
rect 55916 182112 55922 182124
rect 58618 182112 58624 182124
rect 58676 182112 58682 182164
rect 64966 181432 64972 181484
rect 65024 181472 65030 181484
rect 75178 181472 75184 181484
rect 65024 181444 75184 181472
rect 65024 181432 65030 181444
rect 75178 181432 75184 181444
rect 75236 181432 75242 181484
rect 162118 180928 162124 180940
rect 161676 180900 162124 180928
rect 144454 180684 144460 180736
rect 144512 180724 144518 180736
rect 146110 180724 146116 180736
rect 144512 180696 146116 180724
rect 144512 180684 144518 180696
rect 146110 180684 146116 180696
rect 146168 180684 146174 180736
rect 161676 180600 161704 180900
rect 162118 180888 162124 180900
rect 162176 180888 162182 180940
rect 161658 180548 161664 180600
rect 161716 180548 161722 180600
rect 136818 180316 136824 180328
rect 122806 180288 136824 180316
rect 9582 180072 9588 180124
rect 9640 180112 9646 180124
rect 122806 180112 122834 180288
rect 136818 180276 136824 180288
rect 136876 180276 136882 180328
rect 9640 180084 122834 180112
rect 9640 180072 9646 180084
rect 136634 180072 136640 180124
rect 136692 180112 136698 180124
rect 141234 180112 141240 180124
rect 136692 180084 141240 180112
rect 136692 180072 136698 180084
rect 141234 180072 141240 180084
rect 141292 180072 141298 180124
rect 143534 179596 143540 179648
rect 143592 179596 143598 179648
rect 72418 179324 72424 179376
rect 72476 179364 72482 179376
rect 75730 179364 75736 179376
rect 72476 179336 75736 179364
rect 72476 179324 72482 179336
rect 75730 179324 75736 179336
rect 75788 179324 75794 179376
rect 122834 178780 122840 178832
rect 122892 178820 122898 178832
rect 136634 178820 136640 178832
rect 122892 178792 136640 178820
rect 122892 178780 122898 178792
rect 136634 178780 136640 178792
rect 136692 178780 136698 178832
rect 121454 178644 121460 178696
rect 121512 178684 121518 178696
rect 137002 178684 137008 178696
rect 121512 178656 137008 178684
rect 121512 178644 121518 178656
rect 137002 178644 137008 178656
rect 137060 178644 137066 178696
rect 143552 178684 143580 179596
rect 144178 178684 144184 178696
rect 143552 178656 144184 178684
rect 144178 178644 144184 178656
rect 144236 178644 144242 178696
rect 159082 178508 159088 178560
rect 159140 178548 159146 178560
rect 161658 178548 161664 178560
rect 159140 178520 161664 178548
rect 159140 178508 159146 178520
rect 161658 178508 161664 178520
rect 161716 178508 161722 178560
rect 166258 178236 166264 178288
rect 166316 178276 166322 178288
rect 167638 178276 167644 178288
rect 166316 178248 167644 178276
rect 166316 178236 166322 178248
rect 167638 178236 167644 178248
rect 167696 178236 167702 178288
rect 189718 178032 189724 178084
rect 189776 178072 189782 178084
rect 580166 178072 580172 178084
rect 189776 178044 580172 178072
rect 189776 178032 189782 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 61378 177964 61384 178016
rect 61436 178004 61442 178016
rect 65886 178004 65892 178016
rect 61436 177976 65892 178004
rect 61436 177964 61442 177976
rect 65886 177964 65892 177976
rect 65944 177964 65950 178016
rect 140774 177828 140780 177880
rect 140832 177868 140838 177880
rect 141602 177868 141608 177880
rect 140832 177840 141608 177868
rect 140832 177828 140838 177840
rect 141602 177828 141608 177840
rect 141660 177828 141666 177880
rect 124214 177284 124220 177336
rect 124272 177324 124278 177336
rect 137094 177324 137100 177336
rect 124272 177296 137100 177324
rect 124272 177284 124278 177296
rect 137094 177284 137100 177296
rect 137152 177284 137158 177336
rect 75730 176944 75736 176996
rect 75788 176984 75794 176996
rect 77294 176984 77300 176996
rect 75788 176956 77300 176984
rect 75788 176944 75794 176956
rect 77294 176944 77300 176956
rect 77352 176944 77358 176996
rect 159082 176196 159088 176248
rect 159140 176196 159146 176248
rect 3326 176060 3332 176112
rect 3384 176100 3390 176112
rect 9582 176100 9588 176112
rect 3384 176072 9588 176100
rect 3384 176060 3390 176072
rect 9582 176060 9588 176072
rect 9640 176060 9646 176112
rect 125594 175992 125600 176044
rect 125652 176032 125658 176044
rect 137186 176032 137192 176044
rect 125652 176004 137192 176032
rect 125652 175992 125658 176004
rect 137186 175992 137192 176004
rect 137244 175992 137250 176044
rect 128354 175924 128360 175976
rect 128412 175964 128418 175976
rect 137278 175964 137284 175976
rect 128412 175936 137284 175964
rect 128412 175924 128418 175936
rect 137278 175924 137284 175936
rect 137336 175924 137342 175976
rect 159100 175636 159128 176196
rect 355318 175924 355324 175976
rect 355376 175964 355382 175976
rect 371878 175964 371884 175976
rect 355376 175936 371884 175964
rect 355376 175924 355382 175936
rect 371878 175924 371884 175936
rect 371936 175924 371942 175976
rect 159082 175584 159088 175636
rect 159140 175584 159146 175636
rect 165522 174972 165528 175024
rect 165580 174972 165586 175024
rect 163148 174752 163176 174866
rect 165540 174752 165568 174972
rect 163130 174700 163136 174752
rect 163188 174700 163194 174752
rect 165522 174700 165528 174752
rect 165580 174700 165586 174752
rect 3694 174088 3700 174140
rect 3752 174128 3758 174140
rect 179414 174128 179420 174140
rect 3752 174100 179420 174128
rect 3752 174088 3758 174100
rect 179414 174088 179420 174100
rect 179472 174088 179478 174140
rect 77294 173884 77300 173936
rect 77352 173924 77358 173936
rect 77352 173896 78720 173924
rect 77352 173884 77358 173896
rect 65886 173816 65892 173868
rect 65944 173856 65950 173868
rect 66898 173856 66904 173868
rect 65944 173828 66904 173856
rect 65944 173816 65950 173828
rect 66898 173816 66904 173828
rect 66956 173816 66962 173868
rect 78692 173856 78720 173896
rect 133874 173884 133880 173936
rect 133932 173924 133938 173936
rect 135254 173924 135260 173936
rect 133932 173896 135260 173924
rect 133932 173884 133938 173896
rect 135254 173884 135260 173896
rect 135312 173884 135318 173936
rect 81342 173856 81348 173868
rect 78692 173828 81348 173856
rect 81342 173816 81348 173828
rect 81400 173816 81406 173868
rect 140774 173816 140780 173868
rect 140832 173856 140838 173868
rect 141602 173856 141608 173868
rect 140832 173828 141608 173856
rect 140832 173816 140838 173828
rect 141602 173816 141608 173828
rect 141660 173816 141666 173868
rect 131114 173204 131120 173256
rect 131172 173244 131178 173256
rect 137370 173244 137376 173256
rect 131172 173216 137376 173244
rect 131172 173204 131178 173216
rect 137370 173204 137376 173216
rect 137428 173204 137434 173256
rect 126974 173136 126980 173188
rect 127032 173176 127038 173188
rect 140774 173176 140780 173188
rect 127032 173148 140780 173176
rect 127032 173136 127038 173148
rect 140774 173136 140780 173148
rect 140832 173136 140838 173188
rect 135254 172388 135260 172440
rect 135312 172428 135318 172440
rect 138934 172428 138940 172440
rect 135312 172400 138940 172428
rect 135312 172388 135318 172400
rect 138934 172388 138940 172400
rect 138992 172388 138998 172440
rect 132494 172184 132500 172236
rect 132552 172224 132558 172236
rect 137462 172224 137468 172236
rect 132552 172196 137468 172224
rect 132552 172184 132558 172196
rect 137462 172184 137468 172196
rect 137520 172184 137526 172236
rect 138014 171912 138020 171964
rect 138072 171952 138078 171964
rect 140958 171952 140964 171964
rect 138072 171924 140964 171952
rect 138072 171912 138078 171924
rect 140958 171912 140964 171924
rect 141016 171912 141022 171964
rect 160002 171028 160008 171080
rect 160060 171068 160066 171080
rect 163866 171068 163872 171080
rect 160060 171040 163872 171068
rect 160060 171028 160066 171040
rect 163866 171028 163872 171040
rect 163924 171028 163930 171080
rect 57238 170076 57244 170128
rect 57296 170116 57302 170128
rect 60642 170116 60648 170128
rect 57296 170088 60648 170116
rect 57296 170076 57302 170088
rect 60642 170076 60648 170088
rect 60700 170076 60706 170128
rect 35158 168988 35164 169040
rect 35216 169028 35222 169040
rect 182266 169028 182272 169040
rect 35216 169000 182272 169028
rect 35216 168988 35222 169000
rect 182266 168988 182272 169000
rect 182324 168988 182330 169040
rect 68278 168580 68284 168632
rect 68336 168620 68342 168632
rect 69750 168620 69756 168632
rect 68336 168592 69756 168620
rect 68336 168580 68342 168592
rect 69750 168580 69756 168592
rect 69808 168580 69814 168632
rect 60642 166608 60648 166660
rect 60700 166648 60706 166660
rect 62114 166648 62120 166660
rect 60700 166620 62120 166648
rect 60700 166608 60706 166620
rect 62114 166608 62120 166620
rect 62172 166608 62178 166660
rect 130378 165588 130384 165640
rect 130436 165628 130442 165640
rect 580166 165628 580172 165640
rect 130436 165600 580172 165628
rect 130436 165588 130442 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 69750 165520 69756 165572
rect 69808 165560 69814 165572
rect 71038 165560 71044 165572
rect 69808 165532 71044 165560
rect 69808 165520 69814 165532
rect 71038 165520 71044 165532
rect 71096 165520 71102 165572
rect 81434 165520 81440 165572
rect 81492 165560 81498 165572
rect 83458 165560 83464 165572
rect 81492 165532 83464 165560
rect 81492 165520 81498 165532
rect 83458 165520 83464 165532
rect 83516 165520 83522 165572
rect 163866 165520 163872 165572
rect 163924 165560 163930 165572
rect 166258 165560 166264 165572
rect 163924 165532 166264 165560
rect 163924 165520 163930 165532
rect 166258 165520 166264 165532
rect 166316 165520 166322 165572
rect 167638 165520 167644 165572
rect 167696 165560 167702 165572
rect 169018 165560 169024 165572
rect 167696 165532 169024 165560
rect 167696 165520 167702 165532
rect 169018 165520 169024 165532
rect 169076 165520 169082 165572
rect 26878 164840 26884 164892
rect 26936 164880 26942 164892
rect 182358 164880 182364 164892
rect 26936 164852 182364 164880
rect 26936 164840 26942 164852
rect 182358 164840 182364 164852
rect 182416 164840 182422 164892
rect 162854 164772 162860 164824
rect 162912 164812 162918 164824
rect 163590 164812 163596 164824
rect 162912 164784 163596 164812
rect 162912 164772 162918 164784
rect 163590 164772 163596 164784
rect 163648 164772 163654 164824
rect 75178 163480 75184 163532
rect 75236 163520 75242 163532
rect 86218 163520 86224 163532
rect 75236 163492 86224 163520
rect 75236 163480 75242 163492
rect 86218 163480 86224 163492
rect 86276 163480 86282 163532
rect 345658 163480 345664 163532
rect 345716 163520 345722 163532
rect 355318 163520 355324 163532
rect 345716 163492 355324 163520
rect 345716 163480 345722 163492
rect 355318 163480 355324 163492
rect 355376 163480 355382 163532
rect 3326 162868 3332 162920
rect 3384 162908 3390 162920
rect 108390 162908 108396 162920
rect 3384 162880 108396 162908
rect 3384 162868 3390 162880
rect 108390 162868 108396 162880
rect 108448 162868 108454 162920
rect 66898 162800 66904 162852
rect 66956 162840 66962 162852
rect 68278 162840 68284 162852
rect 66956 162812 68284 162840
rect 66956 162800 66962 162812
rect 68278 162800 68284 162812
rect 68336 162800 68342 162852
rect 62114 162188 62120 162240
rect 62172 162228 62178 162240
rect 87598 162228 87604 162240
rect 62172 162200 87604 162228
rect 62172 162188 62178 162200
rect 87598 162188 87604 162200
rect 87656 162188 87662 162240
rect 32398 162120 32404 162172
rect 32456 162160 32462 162172
rect 182726 162160 182732 162172
rect 32456 162132 182732 162160
rect 32456 162120 32462 162132
rect 182726 162120 182732 162132
rect 182784 162120 182790 162172
rect 3510 160692 3516 160744
rect 3568 160732 3574 160744
rect 179598 160732 179604 160744
rect 3568 160704 179604 160732
rect 3568 160692 3574 160704
rect 179598 160692 179604 160704
rect 179656 160692 179662 160744
rect 376018 160120 376024 160132
rect 373966 160092 376024 160120
rect 373258 160012 373264 160064
rect 373316 160052 373322 160064
rect 373966 160052 373994 160092
rect 376018 160080 376024 160092
rect 376076 160080 376082 160132
rect 373316 160024 373994 160052
rect 373316 160012 373322 160024
rect 58618 159400 58624 159452
rect 58676 159440 58682 159452
rect 81434 159440 81440 159452
rect 58676 159412 81440 159440
rect 58676 159400 58682 159412
rect 81434 159400 81440 159412
rect 81492 159400 81498 159452
rect 23474 159332 23480 159384
rect 23532 159372 23538 159384
rect 180978 159372 180984 159384
rect 23532 159344 180984 159372
rect 23532 159332 23538 159344
rect 180978 159332 180984 159344
rect 181036 159332 181042 159384
rect 81434 157972 81440 158024
rect 81492 158012 81498 158024
rect 84746 158012 84752 158024
rect 81492 157984 84752 158012
rect 81492 157972 81498 157984
rect 84746 157972 84752 157984
rect 84804 157972 84810 158024
rect 83458 157292 83464 157344
rect 83516 157332 83522 157344
rect 84838 157332 84844 157344
rect 83516 157304 84844 157332
rect 83516 157292 83522 157304
rect 84838 157292 84844 157304
rect 84896 157292 84902 157344
rect 84746 156612 84752 156664
rect 84804 156652 84810 156664
rect 89070 156652 89076 156664
rect 84804 156624 89076 156652
rect 84804 156612 84810 156624
rect 89070 156612 89076 156624
rect 89128 156612 89134 156664
rect 118234 156612 118240 156664
rect 118292 156652 118298 156664
rect 417418 156652 417424 156664
rect 118292 156624 417424 156652
rect 118292 156612 118298 156624
rect 417418 156612 417424 156624
rect 417476 156612 417482 156664
rect 118326 155184 118332 155236
rect 118384 155224 118390 155236
rect 414658 155224 414664 155236
rect 118384 155196 414664 155224
rect 118384 155184 118390 155196
rect 414658 155184 414664 155196
rect 414716 155184 414722 155236
rect 87598 154504 87604 154556
rect 87656 154544 87662 154556
rect 90358 154544 90364 154556
rect 87656 154516 90364 154544
rect 87656 154504 87662 154516
rect 90358 154504 90364 154516
rect 90416 154504 90422 154556
rect 118510 153824 118516 153876
rect 118568 153864 118574 153876
rect 400950 153864 400956 153876
rect 118568 153836 400956 153864
rect 118568 153824 118574 153836
rect 400950 153824 400956 153836
rect 401008 153824 401014 153876
rect 71038 153144 71044 153196
rect 71096 153184 71102 153196
rect 73798 153184 73804 153196
rect 71096 153156 73804 153184
rect 71096 153144 71102 153156
rect 73798 153144 73804 153156
rect 73856 153144 73862 153196
rect 118418 152464 118424 152516
rect 118476 152504 118482 152516
rect 399570 152504 399576 152516
rect 118476 152476 399576 152504
rect 118476 152464 118482 152476
rect 399570 152464 399576 152476
rect 399628 152464 399634 152516
rect 381538 151852 381544 151904
rect 381596 151892 381602 151904
rect 384298 151892 384304 151904
rect 381596 151864 384304 151892
rect 381596 151852 381602 151864
rect 384298 151852 384304 151864
rect 384356 151852 384362 151904
rect 181438 151784 181444 151836
rect 181496 151824 181502 151836
rect 579982 151824 579988 151836
rect 181496 151796 579988 151824
rect 181496 151784 181502 151796
rect 579982 151784 579988 151796
rect 580040 151784 580046 151836
rect 118786 151036 118792 151088
rect 118844 151076 118850 151088
rect 580534 151076 580540 151088
rect 118844 151048 580540 151076
rect 118844 151036 118850 151048
rect 580534 151036 580540 151048
rect 580592 151036 580598 151088
rect 165430 150900 165436 150952
rect 165488 150940 165494 150952
rect 167730 150940 167736 150952
rect 165488 150912 167736 150940
rect 165488 150900 165494 150912
rect 167730 150900 167736 150912
rect 167788 150900 167794 150952
rect 89070 149812 89076 149864
rect 89128 149852 89134 149864
rect 91002 149852 91008 149864
rect 89128 149824 91008 149852
rect 89128 149812 89134 149824
rect 91002 149812 91008 149824
rect 91060 149812 91066 149864
rect 319438 149744 319444 149796
rect 319496 149784 319502 149796
rect 345658 149784 345664 149796
rect 319496 149756 345664 149784
rect 319496 149744 319502 149756
rect 345658 149744 345664 149756
rect 345716 149744 345722 149796
rect 120994 149676 121000 149728
rect 121052 149716 121058 149728
rect 429194 149716 429200 149728
rect 121052 149688 429200 149716
rect 121052 149676 121058 149688
rect 429194 149676 429200 149688
rect 429252 149676 429258 149728
rect 86218 149200 86224 149252
rect 86276 149240 86282 149252
rect 88978 149240 88984 149252
rect 86276 149212 88984 149240
rect 86276 149200 86282 149212
rect 88978 149200 88984 149212
rect 89036 149200 89042 149252
rect 3510 149064 3516 149116
rect 3568 149104 3574 149116
rect 178678 149104 178684 149116
rect 3568 149076 178684 149104
rect 3568 149064 3574 149076
rect 178678 149064 178684 149076
rect 178736 149064 178742 149116
rect 91002 148996 91008 149048
rect 91060 149036 91066 149048
rect 92474 149036 92480 149048
rect 91060 149008 92480 149036
rect 91060 148996 91066 149008
rect 92474 148996 92480 149008
rect 92532 148996 92538 149048
rect 166258 147296 166264 147348
rect 166316 147336 166322 147348
rect 168374 147336 168380 147348
rect 166316 147308 168380 147336
rect 166316 147296 166322 147308
rect 168374 147296 168380 147308
rect 168432 147296 168438 147348
rect 169018 146888 169024 146940
rect 169076 146928 169082 146940
rect 175182 146928 175188 146940
rect 169076 146900 175188 146928
rect 169076 146888 169082 146900
rect 175182 146888 175188 146900
rect 175240 146888 175246 146940
rect 108298 146208 108304 146260
rect 108356 146248 108362 146260
rect 109678 146248 109684 146260
rect 108356 146220 109684 146248
rect 108356 146208 108362 146220
rect 109678 146208 109684 146220
rect 109736 146208 109742 146260
rect 118970 145528 118976 145580
rect 119028 145568 119034 145580
rect 494054 145568 494060 145580
rect 119028 145540 494060 145568
rect 119028 145528 119034 145540
rect 494054 145528 494060 145540
rect 494112 145528 494118 145580
rect 373350 144236 373356 144288
rect 373408 144276 373414 144288
rect 381538 144276 381544 144288
rect 373408 144248 381544 144276
rect 373408 144236 373414 144248
rect 381538 144236 381544 144248
rect 381596 144236 381602 144288
rect 118878 144168 118884 144220
rect 118936 144208 118942 144220
rect 558914 144208 558920 144220
rect 118936 144180 558920 144208
rect 118936 144168 118942 144180
rect 558914 144168 558920 144180
rect 558972 144168 558978 144220
rect 175274 143556 175280 143608
rect 175332 143596 175338 143608
rect 175332 143568 176700 143596
rect 175332 143556 175338 143568
rect 151814 143488 151820 143540
rect 151872 143528 151878 143540
rect 157426 143528 157432 143540
rect 151872 143500 157432 143528
rect 151872 143488 151878 143500
rect 157426 143488 157432 143500
rect 157484 143488 157490 143540
rect 167730 143488 167736 143540
rect 167788 143528 167794 143540
rect 169938 143528 169944 143540
rect 167788 143500 169944 143528
rect 167788 143488 167794 143500
rect 169938 143488 169944 143500
rect 169996 143488 170002 143540
rect 176672 143528 176700 143568
rect 178218 143528 178224 143540
rect 176672 143500 178224 143528
rect 178218 143488 178224 143500
rect 178276 143488 178282 143540
rect 164050 143420 164056 143472
rect 164108 143460 164114 143472
rect 166074 143460 166080 143472
rect 164108 143432 166080 143460
rect 164108 143420 164114 143432
rect 166074 143420 166080 143432
rect 166132 143420 166138 143472
rect 137738 143148 137744 143200
rect 137796 143188 137802 143200
rect 139394 143188 139400 143200
rect 137796 143160 139400 143188
rect 137796 143148 137802 143160
rect 139394 143148 139400 143160
rect 139452 143148 139458 143200
rect 162762 143080 162768 143132
rect 162820 143120 162826 143132
rect 166166 143120 166172 143132
rect 162820 143092 166172 143120
rect 162820 143080 162826 143092
rect 166166 143080 166172 143092
rect 166224 143080 166230 143132
rect 162854 142944 162860 142996
rect 162912 142984 162918 142996
rect 174630 142984 174636 142996
rect 162912 142956 174636 142984
rect 162912 142944 162918 142956
rect 174630 142944 174636 142956
rect 174688 142944 174694 142996
rect 150434 142876 150440 142928
rect 150492 142916 150498 142928
rect 154574 142916 154580 142928
rect 150492 142888 154580 142916
rect 150492 142876 150498 142888
rect 154574 142876 154580 142888
rect 154632 142876 154638 142928
rect 164234 142876 164240 142928
rect 164292 142916 164298 142928
rect 176194 142916 176200 142928
rect 164292 142888 176200 142916
rect 164292 142876 164298 142888
rect 176194 142876 176200 142888
rect 176252 142876 176258 142928
rect 92474 142808 92480 142860
rect 92532 142848 92538 142860
rect 104894 142848 104900 142860
rect 92532 142820 104900 142848
rect 92532 142808 92538 142820
rect 104894 142808 104900 142820
rect 104952 142808 104958 142860
rect 118142 142808 118148 142860
rect 118200 142848 118206 142860
rect 130378 142848 130384 142860
rect 118200 142820 130384 142848
rect 118200 142808 118206 142820
rect 130378 142808 130384 142820
rect 130436 142808 130442 142860
rect 163130 142808 163136 142860
rect 163188 142848 163194 142860
rect 178034 142848 178040 142860
rect 163188 142820 178040 142848
rect 163188 142808 163194 142820
rect 178034 142808 178040 142820
rect 178092 142808 178098 142860
rect 149054 142128 149060 142180
rect 149112 142168 149118 142180
rect 152734 142168 152740 142180
rect 149112 142140 152740 142168
rect 149112 142128 149118 142140
rect 152734 142128 152740 142140
rect 152792 142128 152798 142180
rect 45278 141516 45284 141568
rect 45336 141556 45342 141568
rect 182450 141556 182456 141568
rect 45336 141528 182456 141556
rect 45336 141516 45342 141528
rect 182450 141516 182456 141528
rect 182508 141516 182514 141568
rect 28258 141448 28264 141500
rect 28316 141488 28322 141500
rect 182542 141488 182548 141500
rect 28316 141460 182548 141488
rect 28316 141448 28322 141460
rect 182542 141448 182548 141460
rect 182600 141448 182606 141500
rect 104894 141380 104900 141432
rect 104952 141420 104958 141432
rect 107654 141420 107660 141432
rect 104952 141392 107660 141420
rect 104952 141380 104958 141392
rect 107654 141380 107660 141392
rect 107712 141380 107718 141432
rect 117958 141380 117964 141432
rect 118016 141420 118022 141432
rect 413278 141420 413284 141432
rect 118016 141392 413284 141420
rect 118016 141380 118022 141392
rect 413278 141380 413284 141392
rect 413336 141380 413342 141432
rect 107654 140088 107660 140140
rect 107712 140128 107718 140140
rect 181530 140128 181536 140140
rect 107712 140100 181536 140128
rect 107712 140088 107718 140100
rect 181530 140088 181536 140100
rect 181588 140088 181594 140140
rect 25498 140020 25504 140072
rect 25556 140060 25562 140072
rect 182634 140060 182640 140072
rect 25556 140032 182640 140060
rect 25556 140020 25562 140032
rect 182634 140020 182640 140032
rect 182692 140020 182698 140072
rect 88978 139476 88984 139528
rect 89036 139516 89042 139528
rect 91370 139516 91376 139528
rect 89036 139488 91376 139516
rect 89036 139476 89042 139488
rect 91370 139476 91376 139488
rect 91428 139476 91434 139528
rect 118050 139476 118056 139528
rect 118108 139516 118114 139528
rect 122098 139516 122104 139528
rect 118108 139488 122104 139516
rect 118108 139476 118114 139488
rect 122098 139476 122104 139488
rect 122156 139476 122162 139528
rect 3694 139408 3700 139460
rect 3752 139448 3758 139460
rect 181070 139448 181076 139460
rect 3752 139420 181076 139448
rect 3752 139408 3758 139420
rect 181070 139408 181076 139420
rect 181128 139408 181134 139460
rect 316678 139408 316684 139460
rect 316736 139448 316742 139460
rect 319438 139448 319444 139460
rect 316736 139420 319444 139448
rect 316736 139408 316742 139420
rect 319438 139408 319444 139420
rect 319496 139408 319502 139460
rect 178218 139340 178224 139392
rect 178276 139380 178282 139392
rect 180150 139380 180156 139392
rect 178276 139352 180156 139380
rect 178276 139340 178282 139352
rect 180150 139340 180156 139352
rect 180208 139340 180214 139392
rect 178678 139272 178684 139324
rect 178736 139312 178742 139324
rect 182174 139312 182180 139324
rect 178736 139284 182180 139312
rect 178736 139272 178742 139284
rect 182174 139272 182180 139284
rect 182232 139272 182238 139324
rect 188338 137980 188344 138032
rect 188396 138020 188402 138032
rect 580166 138020 580172 138032
rect 188396 137992 580172 138020
rect 188396 137980 188402 137992
rect 580166 137980 580172 137992
rect 580224 137980 580230 138032
rect 21450 136688 21456 136740
rect 21508 136728 21514 136740
rect 117314 136728 117320 136740
rect 21508 136700 117320 136728
rect 21508 136688 21514 136700
rect 117314 136688 117320 136700
rect 117372 136688 117378 136740
rect 3510 136620 3516 136672
rect 3568 136660 3574 136672
rect 120902 136660 120908 136672
rect 3568 136632 120908 136660
rect 3568 136620 3574 136632
rect 120902 136620 120908 136632
rect 120960 136620 120966 136672
rect 3510 135940 3516 135992
rect 3568 135980 3574 135992
rect 3694 135980 3700 135992
rect 3568 135952 3700 135980
rect 3568 135940 3574 135952
rect 3694 135940 3700 135952
rect 3752 135940 3758 135992
rect 90358 135872 90364 135924
rect 90416 135912 90422 135924
rect 105538 135912 105544 135924
rect 90416 135884 105544 135912
rect 90416 135872 90422 135884
rect 105538 135872 105544 135884
rect 105596 135872 105602 135924
rect 97258 135260 97264 135312
rect 97316 135300 97322 135312
rect 117314 135300 117320 135312
rect 97316 135272 117320 135300
rect 97316 135260 97322 135272
rect 117314 135260 117320 135272
rect 117372 135260 117378 135312
rect 18690 133900 18696 133952
rect 18748 133940 18754 133952
rect 117314 133940 117320 133952
rect 18748 133912 117320 133940
rect 18748 133900 18754 133912
rect 117314 133900 117320 133912
rect 117372 133900 117378 133952
rect 108390 133832 108396 133884
rect 108448 133872 108454 133884
rect 117406 133872 117412 133884
rect 108448 133844 117412 133872
rect 108448 133832 108454 133844
rect 117406 133832 117412 133844
rect 117464 133832 117470 133884
rect 91370 132812 91376 132864
rect 91428 132852 91434 132864
rect 94222 132852 94228 132864
rect 91428 132824 94228 132852
rect 91428 132812 91434 132824
rect 94222 132812 94228 132824
rect 94280 132812 94286 132864
rect 22738 132404 22744 132456
rect 22796 132444 22802 132456
rect 117314 132444 117320 132456
rect 22796 132416 117320 132444
rect 22796 132404 22802 132416
rect 117314 132404 117320 132416
rect 117372 132404 117378 132456
rect 84838 131724 84844 131776
rect 84896 131764 84902 131776
rect 86310 131764 86316 131776
rect 84896 131736 86316 131764
rect 84896 131724 84902 131736
rect 86310 131724 86316 131736
rect 86368 131724 86374 131776
rect 369854 131112 369860 131164
rect 369912 131152 369918 131164
rect 373258 131152 373264 131164
rect 369912 131124 373264 131152
rect 369912 131112 369918 131124
rect 373258 131112 373264 131124
rect 373316 131112 373322 131164
rect 21358 131044 21364 131096
rect 21416 131084 21422 131096
rect 117314 131084 117320 131096
rect 21416 131056 117320 131084
rect 21416 131044 21422 131056
rect 117314 131044 117320 131056
rect 117372 131044 117378 131096
rect 86310 130840 86316 130892
rect 86368 130880 86374 130892
rect 87598 130880 87604 130892
rect 86368 130852 87604 130880
rect 86368 130840 86374 130852
rect 87598 130840 87604 130852
rect 87656 130840 87662 130892
rect 109678 129752 109684 129804
rect 109736 129792 109742 129804
rect 111058 129792 111064 129804
rect 109736 129764 111064 129792
rect 109736 129752 109742 129764
rect 111058 129752 111064 129764
rect 111116 129752 111122 129804
rect 17218 129684 17224 129736
rect 17276 129724 17282 129736
rect 117314 129724 117320 129736
rect 17276 129696 117320 129724
rect 17276 129684 17282 129696
rect 117314 129684 117320 129696
rect 117372 129684 117378 129736
rect 355962 129004 355968 129056
rect 356020 129044 356026 129056
rect 369854 129044 369860 129056
rect 356020 129016 369860 129044
rect 356020 129004 356026 129016
rect 369854 129004 369860 129016
rect 369912 129004 369918 129056
rect 14458 128256 14464 128308
rect 14516 128296 14522 128308
rect 117314 128296 117320 128308
rect 14516 128268 117320 128296
rect 14516 128256 14522 128268
rect 117314 128256 117320 128268
rect 117372 128256 117378 128308
rect 68278 127576 68284 127628
rect 68336 127616 68342 127628
rect 71038 127616 71044 127628
rect 68336 127588 71044 127616
rect 68336 127576 68342 127588
rect 71038 127576 71044 127588
rect 71096 127576 71102 127628
rect 328914 127576 328920 127628
rect 328972 127616 328978 127628
rect 355962 127616 355968 127628
rect 328972 127588 355968 127616
rect 328972 127576 328978 127588
rect 355962 127576 355968 127588
rect 356020 127576 356026 127628
rect 13078 126896 13084 126948
rect 13136 126936 13142 126948
rect 117314 126936 117320 126948
rect 13136 126908 117320 126936
rect 13136 126896 13142 126908
rect 117314 126896 117320 126908
rect 117372 126896 117378 126948
rect 94222 126828 94228 126880
rect 94280 126868 94286 126880
rect 100018 126868 100024 126880
rect 94280 126840 100024 126868
rect 94280 126828 94286 126840
rect 100018 126828 100024 126840
rect 100076 126828 100082 126880
rect 105538 126828 105544 126880
rect 105596 126868 105602 126880
rect 109678 126868 109684 126880
rect 105596 126840 109684 126868
rect 105596 126828 105602 126840
rect 109678 126828 109684 126840
rect 109736 126828 109742 126880
rect 326706 126012 326712 126064
rect 326764 126052 326770 126064
rect 328914 126052 328920 126064
rect 326764 126024 328920 126052
rect 326764 126012 326770 126024
rect 328914 126012 328920 126024
rect 328972 126012 328978 126064
rect 180058 125604 180064 125656
rect 180116 125644 180122 125656
rect 579798 125644 579804 125656
rect 180116 125616 579804 125644
rect 180116 125604 180122 125616
rect 579798 125604 579804 125616
rect 579856 125604 579862 125656
rect 73798 124788 73804 124840
rect 73856 124828 73862 124840
rect 75822 124828 75828 124840
rect 73856 124800 75828 124828
rect 73856 124788 73862 124800
rect 75822 124788 75828 124800
rect 75880 124788 75886 124840
rect 322934 124448 322940 124500
rect 322992 124488 322998 124500
rect 326706 124488 326712 124500
rect 322992 124460 326712 124488
rect 322992 124448 322998 124460
rect 326706 124448 326712 124460
rect 326764 124448 326770 124500
rect 18598 124108 18604 124160
rect 18656 124148 18662 124160
rect 117314 124148 117320 124160
rect 18656 124120 117320 124148
rect 18656 124108 18662 124120
rect 117314 124108 117320 124120
rect 117372 124108 117378 124160
rect 367738 123632 367744 123684
rect 367796 123672 367802 123684
rect 373350 123672 373356 123684
rect 367796 123644 373356 123672
rect 367796 123632 367802 123644
rect 373350 123632 373356 123644
rect 373408 123632 373414 123684
rect 304258 123428 304264 123480
rect 304316 123468 304322 123480
rect 322934 123468 322940 123480
rect 304316 123440 322940 123468
rect 304316 123428 304322 123440
rect 322934 123428 322940 123440
rect 322992 123428 322998 123480
rect 10318 122748 10324 122800
rect 10376 122788 10382 122800
rect 117314 122788 117320 122800
rect 10376 122760 117320 122788
rect 10376 122748 10382 122760
rect 117314 122748 117320 122760
rect 117372 122748 117378 122800
rect 109678 122476 109684 122528
rect 109736 122516 109742 122528
rect 113818 122516 113824 122528
rect 109736 122488 113824 122516
rect 109736 122476 109742 122488
rect 113818 122476 113824 122488
rect 113876 122476 113882 122528
rect 87598 121796 87604 121848
rect 87656 121836 87662 121848
rect 91002 121836 91008 121848
rect 87656 121808 91008 121836
rect 87656 121796 87662 121808
rect 91002 121796 91008 121808
rect 91060 121796 91066 121848
rect 8938 121388 8944 121440
rect 8996 121428 9002 121440
rect 117314 121428 117320 121440
rect 8996 121400 117320 121428
rect 8996 121388 9002 121400
rect 117314 121388 117320 121400
rect 117372 121388 117378 121440
rect 7558 120028 7564 120080
rect 7616 120068 7622 120080
rect 117314 120068 117320 120080
rect 7616 120040 117320 120068
rect 7616 120028 7622 120040
rect 117314 120028 117320 120040
rect 117372 120028 117378 120080
rect 91094 119892 91100 119944
rect 91152 119932 91158 119944
rect 93118 119932 93124 119944
rect 91152 119904 93124 119932
rect 91152 119892 91158 119904
rect 93118 119892 93124 119904
rect 93176 119892 93182 119944
rect 181530 119824 181536 119876
rect 181588 119864 181594 119876
rect 182266 119864 182272 119876
rect 181588 119836 182272 119864
rect 181588 119824 181594 119836
rect 182266 119824 182272 119836
rect 182324 119824 182330 119876
rect 75914 119076 75920 119128
rect 75972 119116 75978 119128
rect 78582 119116 78588 119128
rect 75972 119088 78588 119116
rect 75972 119076 75978 119088
rect 78582 119076 78588 119088
rect 78640 119076 78646 119128
rect 4798 118600 4804 118652
rect 4856 118640 4862 118652
rect 117314 118640 117320 118652
rect 4856 118612 117320 118640
rect 4856 118600 4862 118612
rect 117314 118600 117320 118612
rect 117372 118600 117378 118652
rect 71038 117920 71044 117972
rect 71096 117960 71102 117972
rect 77294 117960 77300 117972
rect 71096 117932 77300 117960
rect 71096 117920 71102 117932
rect 77294 117920 77300 117932
rect 77352 117920 77358 117972
rect 40034 117240 40040 117292
rect 40092 117280 40098 117292
rect 117314 117280 117320 117292
rect 40092 117252 117320 117280
rect 40092 117240 40098 117252
rect 117314 117240 117320 117252
rect 117372 117240 117378 117292
rect 77294 116016 77300 116068
rect 77352 116056 77358 116068
rect 79318 116056 79324 116068
rect 77352 116028 79324 116056
rect 77352 116016 77358 116028
rect 79318 116016 79324 116028
rect 79376 116016 79382 116068
rect 100018 115880 100024 115932
rect 100076 115920 100082 115932
rect 117314 115920 117320 115932
rect 100076 115892 117320 115920
rect 100076 115880 100082 115892
rect 117314 115880 117320 115892
rect 117372 115880 117378 115932
rect 180150 114520 180156 114572
rect 180208 114560 180214 114572
rect 180208 114532 180794 114560
rect 180208 114520 180214 114532
rect 78582 114452 78588 114504
rect 78640 114492 78646 114504
rect 117314 114492 117320 114504
rect 78640 114464 117320 114492
rect 78640 114452 78646 114464
rect 117314 114452 117320 114464
rect 117372 114452 117378 114504
rect 180766 114492 180794 114532
rect 182174 114492 182180 114504
rect 180766 114464 182180 114492
rect 182174 114452 182180 114464
rect 182232 114452 182238 114504
rect 93118 113092 93124 113144
rect 93176 113132 93182 113144
rect 117314 113132 117320 113144
rect 93176 113104 117320 113132
rect 93176 113092 93182 113104
rect 117314 113092 117320 113104
rect 117372 113092 117378 113144
rect 79318 112412 79324 112464
rect 79376 112452 79382 112464
rect 88242 112452 88248 112464
rect 79376 112424 88248 112452
rect 79376 112412 79382 112424
rect 88242 112412 88248 112424
rect 88300 112412 88306 112464
rect 180150 111800 180156 111852
rect 180208 111840 180214 111852
rect 580166 111840 580172 111852
rect 180208 111812 580172 111840
rect 180208 111800 180214 111812
rect 580166 111800 580172 111812
rect 580224 111800 580230 111852
rect 2958 111732 2964 111784
rect 3016 111772 3022 111784
rect 18690 111772 18696 111784
rect 3016 111744 18696 111772
rect 3016 111732 3022 111744
rect 18690 111732 18696 111744
rect 18748 111732 18754 111784
rect 88242 111732 88248 111784
rect 88300 111772 88306 111784
rect 117314 111772 117320 111784
rect 88300 111744 117320 111772
rect 88300 111732 88306 111744
rect 117314 111732 117320 111744
rect 117372 111732 117378 111784
rect 111058 109012 111064 109064
rect 111116 109052 111122 109064
rect 112438 109052 112444 109064
rect 111116 109024 112444 109052
rect 111116 109012 111122 109024
rect 112438 109012 112444 109024
rect 112496 109012 112502 109064
rect 113818 109012 113824 109064
rect 113876 109052 113882 109064
rect 120626 109052 120632 109064
rect 113876 109024 120632 109052
rect 113876 109012 113882 109024
rect 120626 109012 120632 109024
rect 120684 109012 120690 109064
rect 183278 107584 183284 107636
rect 183336 107624 183342 107636
rect 304258 107624 304264 107636
rect 183336 107596 304264 107624
rect 183336 107584 183342 107596
rect 304258 107584 304264 107596
rect 304316 107584 304322 107636
rect 183278 106224 183284 106276
rect 183336 106264 183342 106276
rect 396626 106264 396632 106276
rect 183336 106236 396632 106264
rect 183336 106224 183342 106236
rect 396626 106224 396632 106236
rect 396684 106224 396690 106276
rect 183278 104796 183284 104848
rect 183336 104836 183342 104848
rect 404998 104836 405004 104848
rect 183336 104808 405004 104836
rect 183336 104796 183342 104808
rect 404998 104796 405004 104808
rect 405056 104796 405062 104848
rect 183278 103436 183284 103488
rect 183336 103476 183342 103488
rect 403618 103476 403624 103488
rect 183336 103448 403624 103476
rect 183336 103436 183342 103448
rect 403618 103436 403624 103448
rect 403676 103436 403682 103488
rect 112438 103096 112444 103148
rect 112496 103136 112502 103148
rect 115382 103136 115388 103148
rect 112496 103108 115388 103136
rect 112496 103096 112502 103108
rect 115382 103096 115388 103108
rect 115440 103096 115446 103148
rect 183278 102076 183284 102128
rect 183336 102116 183342 102128
rect 400858 102116 400864 102128
rect 183336 102088 400864 102116
rect 183336 102076 183342 102088
rect 400858 102076 400864 102088
rect 400916 102076 400922 102128
rect 183186 100648 183192 100700
rect 183244 100688 183250 100700
rect 399478 100688 399484 100700
rect 183244 100660 399484 100688
rect 183244 100648 183250 100660
rect 399478 100648 399484 100660
rect 399536 100648 399542 100700
rect 115382 100308 115388 100360
rect 115440 100348 115446 100360
rect 117314 100348 117320 100360
rect 115440 100320 117320 100348
rect 115440 100308 115446 100320
rect 117314 100308 117320 100320
rect 117372 100308 117378 100360
rect 182818 99356 182824 99408
rect 182876 99396 182882 99408
rect 580166 99396 580172 99408
rect 182876 99368 580172 99396
rect 182876 99356 182882 99368
rect 580166 99356 580172 99368
rect 580224 99356 580230 99408
rect 183186 99288 183192 99340
rect 183244 99328 183250 99340
rect 531958 99328 531964 99340
rect 183244 99300 531964 99328
rect 183244 99288 183250 99300
rect 531958 99288 531964 99300
rect 532016 99288 532022 99340
rect 117314 97928 117320 97980
rect 117372 97968 117378 97980
rect 120810 97968 120816 97980
rect 117372 97940 120816 97968
rect 117372 97928 117378 97940
rect 120810 97928 120816 97940
rect 120868 97928 120874 97980
rect 183186 97928 183192 97980
rect 183244 97968 183250 97980
rect 530578 97968 530584 97980
rect 183244 97940 530584 97968
rect 183244 97928 183250 97940
rect 530578 97928 530584 97940
rect 530636 97928 530642 97980
rect 183186 96568 183192 96620
rect 183244 96608 183250 96620
rect 526438 96608 526444 96620
rect 183244 96580 526444 96608
rect 183244 96568 183250 96580
rect 526438 96568 526444 96580
rect 526496 96568 526502 96620
rect 183462 95140 183468 95192
rect 183520 95180 183526 95192
rect 525058 95180 525064 95192
rect 183520 95152 525064 95180
rect 183520 95140 183526 95152
rect 525058 95140 525064 95152
rect 525116 95140 525122 95192
rect 183462 93780 183468 93832
rect 183520 93820 183526 93832
rect 410518 93820 410524 93832
rect 183520 93792 410524 93820
rect 183520 93780 183526 93792
rect 410518 93780 410524 93792
rect 410576 93780 410582 93832
rect 183462 92420 183468 92472
rect 183520 92460 183526 92472
rect 409138 92460 409144 92472
rect 183520 92432 409144 92460
rect 183520 92420 183526 92432
rect 409138 92420 409144 92432
rect 409196 92420 409202 92472
rect 183462 90992 183468 91044
rect 183520 91032 183526 91044
rect 407758 91032 407764 91044
rect 183520 91004 407764 91032
rect 183520 90992 183526 91004
rect 407758 90992 407764 91004
rect 407816 90992 407822 91044
rect 183462 89632 183468 89684
rect 183520 89672 183526 89684
rect 406378 89672 406384 89684
rect 183520 89644 406384 89672
rect 183520 89632 183526 89644
rect 406378 89632 406384 89644
rect 406436 89632 406442 89684
rect 305638 88952 305644 89004
rect 305696 88992 305702 89004
rect 316678 88992 316684 89004
rect 305696 88964 316684 88992
rect 305696 88952 305702 88964
rect 316678 88952 316684 88964
rect 316736 88952 316742 89004
rect 183462 88272 183468 88324
rect 183520 88312 183526 88324
rect 192478 88312 192484 88324
rect 183520 88284 192484 88312
rect 183520 88272 183526 88284
rect 192478 88272 192484 88284
rect 192536 88272 192542 88324
rect 182542 86504 182548 86556
rect 182600 86544 182606 86556
rect 189718 86544 189724 86556
rect 182600 86516 189724 86544
rect 182600 86504 182606 86516
rect 189718 86504 189724 86516
rect 189776 86504 189782 86556
rect 182726 84872 182732 84924
rect 182784 84912 182790 84924
rect 188338 84912 188344 84924
rect 182784 84884 188344 84912
rect 182784 84872 182790 84884
rect 188338 84872 188344 84884
rect 188396 84872 188402 84924
rect 3326 84192 3332 84244
rect 3384 84232 3390 84244
rect 120258 84232 120264 84244
rect 3384 84204 120264 84232
rect 3384 84192 3390 84204
rect 120258 84192 120264 84204
rect 120316 84192 120322 84244
rect 293954 83444 293960 83496
rect 294012 83484 294018 83496
rect 305638 83484 305644 83496
rect 294012 83456 305644 83484
rect 294012 83444 294018 83456
rect 305638 83444 305644 83456
rect 305696 83444 305702 83496
rect 178954 82084 178960 82136
rect 179012 82124 179018 82136
rect 580258 82124 580264 82136
rect 179012 82096 580264 82124
rect 179012 82084 179018 82096
rect 580258 82084 580264 82096
rect 580316 82084 580322 82136
rect 179414 80792 179420 80844
rect 179472 80832 179478 80844
rect 580442 80832 580448 80844
rect 179472 80804 580448 80832
rect 179472 80792 179478 80804
rect 580442 80792 580448 80804
rect 580500 80792 580506 80844
rect 118602 80724 118608 80776
rect 118660 80764 118666 80776
rect 579982 80764 579988 80776
rect 118660 80736 579988 80764
rect 118660 80724 118666 80736
rect 579982 80724 579988 80736
rect 580040 80724 580046 80776
rect 580718 80696 580724 80708
rect 166966 80668 174492 80696
rect 120810 80588 120816 80640
rect 120868 80628 120874 80640
rect 121822 80628 121828 80640
rect 120868 80600 121828 80628
rect 120868 80588 120874 80600
rect 121822 80588 121828 80600
rect 121880 80588 121886 80640
rect 166966 80628 166994 80668
rect 174464 80640 174492 80668
rect 176626 80668 580724 80696
rect 158778 80600 166994 80628
rect 143506 80464 146432 80492
rect 125134 80316 125140 80368
rect 125192 80356 125198 80368
rect 143506 80356 143534 80464
rect 125192 80328 143534 80356
rect 125192 80316 125198 80328
rect 124766 80248 124772 80300
rect 124824 80288 124830 80300
rect 124824 80260 132494 80288
rect 124824 80248 124830 80260
rect 124950 80180 124956 80232
rect 125008 80220 125014 80232
rect 125008 80192 130378 80220
rect 125008 80180 125014 80192
rect 123570 80112 123576 80164
rect 123628 80152 123634 80164
rect 123628 80124 129274 80152
rect 123628 80112 123634 80124
rect 123294 80044 123300 80096
rect 123352 80084 123358 80096
rect 123352 80056 126790 80084
rect 123352 80044 123358 80056
rect 123202 79976 123208 80028
rect 123260 80016 123266 80028
rect 123260 79988 126698 80016
rect 123260 79976 123266 79988
rect 122190 79908 122196 79960
rect 122248 79948 122254 79960
rect 125732 79948 125738 79960
rect 122248 79920 125738 79948
rect 122248 79908 122254 79920
rect 125732 79908 125738 79920
rect 125790 79908 125796 79960
rect 126100 79948 126106 79960
rect 126072 79908 126106 79948
rect 126158 79908 126164 79960
rect 126284 79908 126290 79960
rect 126342 79908 126348 79960
rect 126468 79948 126474 79960
rect 126440 79908 126474 79948
rect 126526 79908 126532 79960
rect 124858 79772 124864 79824
rect 124916 79812 124922 79824
rect 125640 79812 125646 79824
rect 124916 79784 125646 79812
rect 124916 79772 124922 79784
rect 125640 79772 125646 79784
rect 125698 79772 125704 79824
rect 43530 79704 43536 79756
rect 43588 79744 43594 79756
rect 116854 79744 116860 79756
rect 43588 79716 116860 79744
rect 43588 79704 43594 79716
rect 116854 79704 116860 79716
rect 116912 79704 116918 79756
rect 123018 79704 123024 79756
rect 123076 79744 123082 79756
rect 126072 79744 126100 79908
rect 126192 79880 126198 79892
rect 123076 79716 126100 79744
rect 126164 79840 126198 79880
rect 126250 79840 126256 79892
rect 123076 79704 123082 79716
rect 126164 79620 126192 79840
rect 126302 79756 126330 79908
rect 126238 79704 126244 79756
rect 126296 79716 126330 79756
rect 126296 79704 126302 79716
rect 126440 79676 126468 79908
rect 126670 79892 126698 79988
rect 126762 79960 126790 80056
rect 129246 79960 129274 80124
rect 130350 79960 130378 80192
rect 130442 79988 131022 80016
rect 126744 79908 126750 79960
rect 126802 79908 126808 79960
rect 127204 79948 127210 79960
rect 126946 79920 127210 79948
rect 126560 79880 126566 79892
rect 126532 79840 126566 79880
rect 126618 79840 126624 79892
rect 126652 79840 126658 79892
rect 126710 79840 126716 79892
rect 126532 79756 126560 79840
rect 126514 79704 126520 79756
rect 126572 79704 126578 79756
rect 126606 79676 126612 79688
rect 126440 79648 126612 79676
rect 126606 79636 126612 79648
rect 126664 79636 126670 79688
rect 39298 79568 39304 79620
rect 39356 79608 39362 79620
rect 125134 79608 125140 79620
rect 39356 79580 125140 79608
rect 39356 79568 39362 79580
rect 125134 79568 125140 79580
rect 125192 79568 125198 79620
rect 126146 79568 126152 79620
rect 126204 79568 126210 79620
rect 126330 79568 126336 79620
rect 126388 79568 126394 79620
rect 120902 79500 120908 79552
rect 120960 79540 120966 79552
rect 125594 79540 125600 79552
rect 120960 79512 125600 79540
rect 120960 79500 120966 79512
rect 125594 79500 125600 79512
rect 125652 79500 125658 79552
rect 125686 79500 125692 79552
rect 125744 79540 125750 79552
rect 126348 79540 126376 79568
rect 125744 79512 126376 79540
rect 125744 79500 125750 79512
rect 126790 79500 126796 79552
rect 126848 79540 126854 79552
rect 126946 79540 126974 79920
rect 127204 79908 127210 79920
rect 127262 79908 127268 79960
rect 127480 79908 127486 79960
rect 127538 79908 127544 79960
rect 127940 79948 127946 79960
rect 127866 79920 127946 79948
rect 127296 79880 127302 79892
rect 127268 79840 127302 79880
rect 127354 79840 127360 79892
rect 127388 79840 127394 79892
rect 127446 79840 127452 79892
rect 127112 79772 127118 79824
rect 127170 79772 127176 79824
rect 127130 79688 127158 79772
rect 127066 79636 127072 79688
rect 127124 79648 127158 79688
rect 127124 79636 127130 79648
rect 127268 79608 127296 79840
rect 127406 79812 127434 79840
rect 127360 79784 127434 79812
rect 127360 79688 127388 79784
rect 127498 79756 127526 79908
rect 127756 79840 127762 79892
rect 127814 79840 127820 79892
rect 127434 79704 127440 79756
rect 127492 79716 127526 79756
rect 127492 79704 127498 79716
rect 127342 79636 127348 79688
rect 127400 79636 127406 79688
rect 127774 79620 127802 79840
rect 127618 79608 127624 79620
rect 127268 79580 127624 79608
rect 127618 79568 127624 79580
rect 127676 79568 127682 79620
rect 127710 79568 127716 79620
rect 127768 79580 127802 79620
rect 127768 79568 127774 79580
rect 126848 79512 126974 79540
rect 126848 79500 126854 79512
rect 116854 79432 116860 79484
rect 116912 79472 116918 79484
rect 116912 79444 126284 79472
rect 116912 79432 116918 79444
rect 120258 79364 120264 79416
rect 120316 79404 120322 79416
rect 126256 79404 126284 79444
rect 126330 79432 126336 79484
rect 126388 79472 126394 79484
rect 127866 79472 127894 79920
rect 127940 79908 127946 79920
rect 127998 79908 128004 79960
rect 128124 79908 128130 79960
rect 128182 79908 128188 79960
rect 128492 79948 128498 79960
rect 128464 79908 128498 79948
rect 128550 79908 128556 79960
rect 128768 79908 128774 79960
rect 128826 79908 128832 79960
rect 129228 79908 129234 79960
rect 129286 79908 129292 79960
rect 130332 79908 130338 79960
rect 130390 79908 130396 79960
rect 128142 79756 128170 79908
rect 128308 79840 128314 79892
rect 128366 79880 128372 79892
rect 128366 79840 128400 79880
rect 128372 79756 128400 79840
rect 128464 79756 128492 79908
rect 128786 79756 128814 79908
rect 128860 79840 128866 79892
rect 128918 79840 128924 79892
rect 129136 79880 129142 79892
rect 128970 79852 129142 79880
rect 128078 79704 128084 79756
rect 128136 79716 128170 79756
rect 128136 79704 128142 79716
rect 128354 79704 128360 79756
rect 128412 79704 128418 79756
rect 128446 79704 128452 79756
rect 128504 79704 128510 79756
rect 128722 79704 128728 79756
rect 128780 79716 128814 79756
rect 128780 79704 128786 79716
rect 127986 79636 127992 79688
rect 128044 79676 128050 79688
rect 128878 79676 128906 79840
rect 128044 79648 128906 79676
rect 128044 79636 128050 79648
rect 128262 79568 128268 79620
rect 128320 79608 128326 79620
rect 128970 79608 128998 79852
rect 129136 79840 129142 79852
rect 129194 79840 129200 79892
rect 129412 79840 129418 79892
rect 129470 79840 129476 79892
rect 129596 79840 129602 79892
rect 129654 79840 129660 79892
rect 129688 79840 129694 79892
rect 129746 79840 129752 79892
rect 129182 79704 129188 79756
rect 129240 79744 129246 79756
rect 129430 79744 129458 79840
rect 129614 79756 129642 79840
rect 129240 79716 129458 79744
rect 129240 79704 129246 79716
rect 129550 79704 129556 79756
rect 129608 79716 129642 79756
rect 129608 79704 129614 79716
rect 129090 79636 129096 79688
rect 129148 79676 129154 79688
rect 129706 79676 129734 79840
rect 129872 79772 129878 79824
rect 129930 79772 129936 79824
rect 129148 79648 129734 79676
rect 129148 79636 129154 79648
rect 128320 79580 128998 79608
rect 128320 79568 128326 79580
rect 128814 79500 128820 79552
rect 128872 79540 128878 79552
rect 129550 79540 129556 79552
rect 128872 79512 129556 79540
rect 128872 79500 128878 79512
rect 129550 79500 129556 79512
rect 129608 79500 129614 79552
rect 129642 79500 129648 79552
rect 129700 79540 129706 79552
rect 129890 79540 129918 79772
rect 130442 79744 130470 79988
rect 130994 79960 131022 79988
rect 132466 79960 132494 80260
rect 132558 80056 133506 80084
rect 130516 79908 130522 79960
rect 130574 79908 130580 79960
rect 130608 79908 130614 79960
rect 130666 79908 130672 79960
rect 130976 79908 130982 79960
rect 131034 79908 131040 79960
rect 131252 79908 131258 79960
rect 131310 79908 131316 79960
rect 131344 79908 131350 79960
rect 131402 79908 131408 79960
rect 131436 79908 131442 79960
rect 131494 79908 131500 79960
rect 131988 79908 131994 79960
rect 132046 79908 132052 79960
rect 132448 79908 132454 79960
rect 132506 79908 132512 79960
rect 130028 79716 130470 79744
rect 130028 79552 130056 79716
rect 130534 79676 130562 79908
rect 130120 79648 130562 79676
rect 129700 79512 129918 79540
rect 129700 79500 129706 79512
rect 130010 79500 130016 79552
rect 130068 79500 130074 79552
rect 126388 79444 127894 79472
rect 126388 79432 126394 79444
rect 128998 79404 129004 79416
rect 120316 79376 126100 79404
rect 126256 79376 129004 79404
rect 120316 79364 120322 79376
rect 3970 79296 3976 79348
rect 4028 79336 4034 79348
rect 4028 79308 118694 79336
rect 4028 79296 4034 79308
rect 118666 79268 118694 79308
rect 125566 79308 125686 79336
rect 125566 79268 125594 79308
rect 118666 79240 125594 79268
rect 119338 79160 119344 79212
rect 119396 79200 119402 79212
rect 119396 79172 125594 79200
rect 119396 79160 119402 79172
rect 125566 78996 125594 79172
rect 125658 79064 125686 79308
rect 126072 79200 126100 79376
rect 128998 79364 129004 79376
rect 129056 79364 129062 79416
rect 129550 79364 129556 79416
rect 129608 79404 129614 79416
rect 130120 79404 130148 79648
rect 130626 79416 130654 79908
rect 131270 79824 131298 79908
rect 130884 79772 130890 79824
rect 130942 79772 130948 79824
rect 131252 79772 131258 79824
rect 131310 79772 131316 79824
rect 130746 79500 130752 79552
rect 130804 79540 130810 79552
rect 130902 79540 130930 79772
rect 131362 79688 131390 79908
rect 131298 79636 131304 79688
rect 131356 79648 131390 79688
rect 131356 79636 131362 79648
rect 131454 79620 131482 79908
rect 131390 79568 131396 79620
rect 131448 79580 131482 79620
rect 131448 79568 131454 79580
rect 130804 79512 130930 79540
rect 130804 79500 130810 79512
rect 131482 79500 131488 79552
rect 131540 79540 131546 79552
rect 132006 79540 132034 79908
rect 132080 79840 132086 79892
rect 132138 79840 132144 79892
rect 132356 79840 132362 79892
rect 132414 79840 132420 79892
rect 131540 79512 132034 79540
rect 132098 79552 132126 79840
rect 132264 79772 132270 79824
rect 132322 79772 132328 79824
rect 132282 79620 132310 79772
rect 132218 79568 132224 79620
rect 132276 79580 132310 79620
rect 132276 79568 132282 79580
rect 132374 79552 132402 79840
rect 132558 79824 132586 80056
rect 133478 79960 133506 80056
rect 134858 79988 135070 80016
rect 134858 79960 134886 79988
rect 132632 79908 132638 79960
rect 132690 79908 132696 79960
rect 132724 79908 132730 79960
rect 132782 79948 132788 79960
rect 132782 79908 132816 79948
rect 133184 79908 133190 79960
rect 133242 79908 133248 79960
rect 133460 79908 133466 79960
rect 133518 79908 133524 79960
rect 133552 79908 133558 79960
rect 133610 79908 133616 79960
rect 133736 79948 133742 79960
rect 133708 79908 133742 79948
rect 133794 79908 133800 79960
rect 133828 79908 133834 79960
rect 133886 79908 133892 79960
rect 133920 79908 133926 79960
rect 133978 79908 133984 79960
rect 134104 79908 134110 79960
rect 134162 79908 134168 79960
rect 134288 79908 134294 79960
rect 134346 79908 134352 79960
rect 134380 79908 134386 79960
rect 134438 79908 134444 79960
rect 134472 79908 134478 79960
rect 134530 79908 134536 79960
rect 134748 79948 134754 79960
rect 134628 79920 134754 79948
rect 132494 79772 132500 79824
rect 132552 79784 132586 79824
rect 132552 79772 132558 79784
rect 132650 79756 132678 79908
rect 132586 79704 132592 79756
rect 132644 79716 132678 79756
rect 132644 79704 132650 79716
rect 132788 79688 132816 79908
rect 133092 79880 133098 79892
rect 132880 79852 133098 79880
rect 132770 79636 132776 79688
rect 132828 79636 132834 79688
rect 132880 79552 132908 79852
rect 133092 79840 133098 79852
rect 133150 79840 133156 79892
rect 133000 79772 133006 79824
rect 133058 79772 133064 79824
rect 133018 79688 133046 79772
rect 133018 79648 133052 79688
rect 133046 79636 133052 79648
rect 133104 79636 133110 79688
rect 133202 79620 133230 79908
rect 133570 79744 133598 79908
rect 133708 79756 133736 79908
rect 133846 79880 133874 79908
rect 133800 79852 133874 79880
rect 133432 79716 133598 79744
rect 133432 79688 133460 79716
rect 133690 79704 133696 79756
rect 133748 79704 133754 79756
rect 133800 79744 133828 79852
rect 133938 79824 133966 79908
rect 134122 79880 134150 79908
rect 134076 79852 134150 79880
rect 134076 79824 134104 79852
rect 133874 79772 133880 79824
rect 133932 79784 133966 79824
rect 133932 79772 133938 79784
rect 134058 79772 134064 79824
rect 134116 79772 134122 79824
rect 134150 79772 134156 79824
rect 134208 79812 134214 79824
rect 134306 79812 134334 79908
rect 134208 79784 134334 79812
rect 134208 79772 134214 79784
rect 133966 79744 133972 79756
rect 133800 79716 133972 79744
rect 133966 79704 133972 79716
rect 134024 79704 134030 79756
rect 134242 79704 134248 79756
rect 134300 79744 134306 79756
rect 134398 79744 134426 79908
rect 134300 79716 134426 79744
rect 134300 79704 134306 79716
rect 133414 79636 133420 79688
rect 133472 79636 133478 79688
rect 133506 79636 133512 79688
rect 133564 79676 133570 79688
rect 134490 79676 134518 79908
rect 133564 79648 134518 79676
rect 133564 79636 133570 79648
rect 133138 79568 133144 79620
rect 133196 79580 133230 79620
rect 134628 79608 134656 79920
rect 134748 79908 134754 79920
rect 134806 79908 134812 79960
rect 134840 79908 134846 79960
rect 134898 79908 134904 79960
rect 134932 79908 134938 79960
rect 134990 79908 134996 79960
rect 134950 79880 134978 79908
rect 134260 79580 134656 79608
rect 134720 79852 134978 79880
rect 133196 79568 133202 79580
rect 132098 79512 132132 79552
rect 131540 79500 131546 79512
rect 132126 79500 132132 79512
rect 132184 79500 132190 79552
rect 132310 79500 132316 79552
rect 132368 79512 132402 79552
rect 132368 79500 132374 79512
rect 132862 79500 132868 79552
rect 132920 79500 132926 79552
rect 133782 79500 133788 79552
rect 133840 79540 133846 79552
rect 134260 79540 134288 79580
rect 134720 79552 134748 79852
rect 134794 79772 134800 79824
rect 134852 79812 134858 79824
rect 135042 79812 135070 79988
rect 140010 79988 140498 80016
rect 135392 79908 135398 79960
rect 135450 79908 135456 79960
rect 135576 79908 135582 79960
rect 135634 79908 135640 79960
rect 135760 79908 135766 79960
rect 135818 79908 135824 79960
rect 136128 79948 136134 79960
rect 135916 79920 136134 79948
rect 135410 79880 135438 79908
rect 134852 79784 135070 79812
rect 135318 79852 135438 79880
rect 134852 79772 134858 79784
rect 135318 79552 135346 79852
rect 135438 79772 135444 79824
rect 135496 79812 135502 79824
rect 135594 79812 135622 79908
rect 135496 79784 135622 79812
rect 135496 79772 135502 79784
rect 133840 79512 134288 79540
rect 133840 79500 133846 79512
rect 134702 79500 134708 79552
rect 134760 79500 134766 79552
rect 135254 79500 135260 79552
rect 135312 79512 135346 79552
rect 135312 79500 135318 79512
rect 135622 79500 135628 79552
rect 135680 79540 135686 79552
rect 135778 79540 135806 79908
rect 135916 79688 135944 79920
rect 136128 79908 136134 79920
rect 136186 79908 136192 79960
rect 136220 79908 136226 79960
rect 136278 79908 136284 79960
rect 137876 79908 137882 79960
rect 137934 79908 137940 79960
rect 138520 79908 138526 79960
rect 138578 79908 138584 79960
rect 138888 79908 138894 79960
rect 138946 79908 138952 79960
rect 138980 79908 138986 79960
rect 139038 79908 139044 79960
rect 139072 79908 139078 79960
rect 139130 79908 139136 79960
rect 139900 79948 139906 79960
rect 139596 79920 139906 79948
rect 136036 79840 136042 79892
rect 136094 79840 136100 79892
rect 136054 79744 136082 79840
rect 136054 79716 136128 79744
rect 135898 79636 135904 79688
rect 135956 79636 135962 79688
rect 136100 79620 136128 79716
rect 136238 79688 136266 79908
rect 137140 79880 137146 79892
rect 137112 79840 137146 79880
rect 137198 79840 137204 79892
rect 137416 79840 137422 79892
rect 137474 79840 137480 79892
rect 137600 79840 137606 79892
rect 137658 79840 137664 79892
rect 137112 79688 137140 79840
rect 136174 79636 136180 79688
rect 136232 79648 136266 79688
rect 136232 79636 136238 79648
rect 137094 79636 137100 79688
rect 137152 79636 137158 79688
rect 137434 79676 137462 79840
rect 137618 79744 137646 79840
rect 137894 79824 137922 79908
rect 138244 79880 138250 79892
rect 138216 79840 138250 79880
rect 138302 79840 138308 79892
rect 137894 79784 137928 79824
rect 137922 79772 137928 79784
rect 137980 79772 137986 79824
rect 138216 79756 138244 79840
rect 137618 79716 137968 79744
rect 137940 79688 137968 79716
rect 138198 79704 138204 79756
rect 138256 79704 138262 79756
rect 137554 79676 137560 79688
rect 137434 79648 137560 79676
rect 137554 79636 137560 79648
rect 137612 79636 137618 79688
rect 137922 79636 137928 79688
rect 137980 79636 137986 79688
rect 136082 79568 136088 79620
rect 136140 79568 136146 79620
rect 138538 79608 138566 79908
rect 138906 79824 138934 79908
rect 138704 79772 138710 79824
rect 138762 79772 138768 79824
rect 138842 79772 138848 79824
rect 138900 79784 138934 79824
rect 138900 79772 138906 79784
rect 138722 79688 138750 79772
rect 138998 79744 139026 79908
rect 139090 79880 139118 79908
rect 139090 79852 139348 79880
rect 138998 79716 139256 79744
rect 139228 79688 139256 79716
rect 138722 79648 138756 79688
rect 138750 79636 138756 79648
rect 138808 79636 138814 79688
rect 139210 79636 139216 79688
rect 139268 79636 139274 79688
rect 138658 79608 138664 79620
rect 138538 79580 138664 79608
rect 138658 79568 138664 79580
rect 138716 79568 138722 79620
rect 139026 79568 139032 79620
rect 139084 79608 139090 79620
rect 139320 79608 139348 79852
rect 139596 79688 139624 79920
rect 139900 79908 139906 79920
rect 139958 79908 139964 79960
rect 139716 79840 139722 79892
rect 139774 79880 139780 79892
rect 139774 79840 139808 79880
rect 139780 79688 139808 79840
rect 140010 79744 140038 79988
rect 140470 79960 140498 79988
rect 140884 79988 141694 80016
rect 140360 79908 140366 79960
rect 140418 79908 140424 79960
rect 140452 79908 140458 79960
rect 140510 79908 140516 79960
rect 140084 79840 140090 79892
rect 140142 79840 140148 79892
rect 140176 79840 140182 79892
rect 140234 79840 140240 79892
rect 140378 79880 140406 79908
rect 140378 79852 140452 79880
rect 139872 79716 140038 79744
rect 139578 79636 139584 79688
rect 139636 79636 139642 79688
rect 139762 79636 139768 79688
rect 139820 79636 139826 79688
rect 139084 79580 139348 79608
rect 139084 79568 139090 79580
rect 135680 79512 135806 79540
rect 135680 79500 135686 79512
rect 130838 79432 130844 79484
rect 130896 79472 130902 79484
rect 130896 79444 132494 79472
rect 130896 79432 130902 79444
rect 129608 79376 130148 79404
rect 129608 79364 129614 79376
rect 130562 79364 130568 79416
rect 130620 79376 130654 79416
rect 132466 79404 132494 79444
rect 133966 79432 133972 79484
rect 134024 79472 134030 79484
rect 135162 79472 135168 79484
rect 134024 79444 135168 79472
rect 134024 79432 134030 79444
rect 135162 79432 135168 79444
rect 135220 79432 135226 79484
rect 139872 79472 139900 79716
rect 139946 79636 139952 79688
rect 140004 79676 140010 79688
rect 140102 79676 140130 79840
rect 140004 79648 140130 79676
rect 140004 79636 140010 79648
rect 140194 79552 140222 79840
rect 140424 79824 140452 79852
rect 140544 79840 140550 79892
rect 140602 79840 140608 79892
rect 140636 79840 140642 79892
rect 140694 79840 140700 79892
rect 140406 79772 140412 79824
rect 140464 79772 140470 79824
rect 140562 79756 140590 79840
rect 140498 79704 140504 79756
rect 140556 79716 140590 79756
rect 140556 79704 140562 79716
rect 140654 79688 140682 79840
rect 140728 79772 140734 79824
rect 140786 79772 140792 79824
rect 140590 79636 140596 79688
rect 140648 79648 140682 79688
rect 140648 79636 140654 79648
rect 140314 79568 140320 79620
rect 140372 79608 140378 79620
rect 140746 79608 140774 79772
rect 140884 79688 140912 79988
rect 141666 79960 141694 79988
rect 145438 79988 145788 80016
rect 145438 79960 145466 79988
rect 141372 79908 141378 79960
rect 141430 79908 141436 79960
rect 141648 79908 141654 79960
rect 141706 79908 141712 79960
rect 141740 79908 141746 79960
rect 141798 79908 141804 79960
rect 141832 79908 141838 79960
rect 141890 79908 141896 79960
rect 142200 79908 142206 79960
rect 142258 79908 142264 79960
rect 142292 79908 142298 79960
rect 142350 79908 142356 79960
rect 142384 79908 142390 79960
rect 142442 79948 142448 79960
rect 142568 79948 142574 79960
rect 142442 79908 142476 79948
rect 141004 79840 141010 79892
rect 141062 79840 141068 79892
rect 141096 79840 141102 79892
rect 141154 79840 141160 79892
rect 140866 79636 140872 79688
rect 140924 79636 140930 79688
rect 141022 79620 141050 79840
rect 140372 79580 140774 79608
rect 140372 79568 140378 79580
rect 140958 79568 140964 79620
rect 141016 79580 141050 79620
rect 141016 79568 141022 79580
rect 140130 79500 140136 79552
rect 140188 79512 140222 79552
rect 140188 79500 140194 79512
rect 140314 79472 140320 79484
rect 139872 79444 140320 79472
rect 140314 79432 140320 79444
rect 140372 79432 140378 79484
rect 141114 79472 141142 79840
rect 141390 79688 141418 79908
rect 141556 79840 141562 79892
rect 141614 79880 141620 79892
rect 141614 79840 141648 79880
rect 141390 79648 141424 79688
rect 141418 79636 141424 79648
rect 141476 79636 141482 79688
rect 141620 79540 141648 79840
rect 141758 79608 141786 79908
rect 141850 79676 141878 79908
rect 142218 79812 142246 79908
rect 142080 79784 142246 79812
rect 141970 79676 141976 79688
rect 141850 79648 141976 79676
rect 141970 79636 141976 79648
rect 142028 79636 142034 79688
rect 142080 79608 142108 79784
rect 142310 79744 142338 79908
rect 142448 79824 142476 79908
rect 142540 79908 142574 79948
rect 142626 79908 142632 79960
rect 142660 79908 142666 79960
rect 142718 79908 142724 79960
rect 143120 79908 143126 79960
rect 143178 79908 143184 79960
rect 143212 79908 143218 79960
rect 143270 79908 143276 79960
rect 143672 79908 143678 79960
rect 143730 79908 143736 79960
rect 143856 79908 143862 79960
rect 143914 79908 143920 79960
rect 144224 79908 144230 79960
rect 144282 79908 144288 79960
rect 144408 79908 144414 79960
rect 144466 79908 144472 79960
rect 144684 79948 144690 79960
rect 144518 79920 144690 79948
rect 142540 79824 142568 79908
rect 142678 79824 142706 79908
rect 142430 79772 142436 79824
rect 142488 79772 142494 79824
rect 142522 79772 142528 79824
rect 142580 79772 142586 79824
rect 142614 79772 142620 79824
rect 142672 79784 142706 79824
rect 143138 79824 143166 79908
rect 143230 79880 143258 79908
rect 143230 79852 143304 79880
rect 143138 79784 143172 79824
rect 142672 79772 142678 79784
rect 143166 79772 143172 79784
rect 143224 79772 143230 79824
rect 142172 79716 142338 79744
rect 142172 79688 142200 79716
rect 142154 79636 142160 79688
rect 142212 79636 142218 79688
rect 142246 79608 142252 79620
rect 141758 79580 141924 79608
rect 142080 79580 142252 79608
rect 141694 79540 141700 79552
rect 141620 79512 141700 79540
rect 141694 79500 141700 79512
rect 141752 79500 141758 79552
rect 141786 79472 141792 79484
rect 141114 79444 141792 79472
rect 141786 79432 141792 79444
rect 141844 79432 141850 79484
rect 132678 79404 132684 79416
rect 132466 79376 132684 79404
rect 130620 79364 130626 79376
rect 132678 79364 132684 79376
rect 132736 79364 132742 79416
rect 139118 79404 139124 79416
rect 135226 79376 139124 79404
rect 135226 79336 135254 79376
rect 139118 79364 139124 79376
rect 139176 79364 139182 79416
rect 141142 79364 141148 79416
rect 141200 79404 141206 79416
rect 141896 79404 141924 79580
rect 142246 79568 142252 79580
rect 142304 79568 142310 79620
rect 142338 79568 142344 79620
rect 142396 79608 142402 79620
rect 143276 79608 143304 79852
rect 143690 79756 143718 79908
rect 143626 79704 143632 79756
rect 143684 79716 143718 79756
rect 143684 79704 143690 79716
rect 143718 79636 143724 79688
rect 143776 79676 143782 79688
rect 143874 79676 143902 79908
rect 144132 79880 144138 79892
rect 144104 79840 144138 79880
rect 144190 79840 144196 79892
rect 143948 79772 143954 79824
rect 144006 79812 144012 79824
rect 144006 79772 144040 79812
rect 144012 79688 144040 79772
rect 143776 79648 143902 79676
rect 143776 79636 143782 79648
rect 143994 79636 144000 79688
rect 144052 79636 144058 79688
rect 142396 79580 143304 79608
rect 144104 79608 144132 79840
rect 144242 79756 144270 79908
rect 144426 79756 144454 79908
rect 144178 79704 144184 79756
rect 144236 79716 144270 79756
rect 144236 79704 144242 79716
rect 144362 79704 144368 79756
rect 144420 79716 144454 79756
rect 144420 79704 144426 79716
rect 144518 79688 144546 79920
rect 144684 79908 144690 79920
rect 144742 79908 144748 79960
rect 145144 79908 145150 79960
rect 145202 79908 145208 79960
rect 145236 79908 145242 79960
rect 145294 79908 145300 79960
rect 145328 79908 145334 79960
rect 145386 79908 145392 79960
rect 145420 79908 145426 79960
rect 145478 79908 145484 79960
rect 145604 79908 145610 79960
rect 145662 79908 145668 79960
rect 144776 79880 144782 79892
rect 144748 79840 144782 79880
rect 144834 79840 144840 79892
rect 144592 79772 144598 79824
rect 144650 79772 144656 79824
rect 144454 79636 144460 79688
rect 144512 79648 144546 79688
rect 144610 79688 144638 79772
rect 144748 79756 144776 79840
rect 145162 79756 145190 79908
rect 145254 79824 145282 79908
rect 145346 79880 145374 79908
rect 145346 79852 145420 79880
rect 145254 79784 145288 79824
rect 145282 79772 145288 79784
rect 145340 79772 145346 79824
rect 144730 79704 144736 79756
rect 144788 79704 144794 79756
rect 145162 79716 145196 79756
rect 145190 79704 145196 79716
rect 145248 79704 145254 79756
rect 144610 79648 144644 79688
rect 144512 79636 144518 79648
rect 144638 79636 144644 79648
rect 144696 79636 144702 79688
rect 145098 79636 145104 79688
rect 145156 79676 145162 79688
rect 145392 79676 145420 79852
rect 145156 79648 145420 79676
rect 145156 79636 145162 79648
rect 144546 79608 144552 79620
rect 144104 79580 144552 79608
rect 142396 79568 142402 79580
rect 144546 79568 144552 79580
rect 144604 79568 144610 79620
rect 145374 79568 145380 79620
rect 145432 79608 145438 79620
rect 145622 79608 145650 79908
rect 145760 79620 145788 79988
rect 146156 79908 146162 79960
rect 146214 79908 146220 79960
rect 145972 79880 145978 79892
rect 145944 79840 145978 79880
rect 146030 79840 146036 79892
rect 145432 79580 145650 79608
rect 145432 79568 145438 79580
rect 145742 79568 145748 79620
rect 145800 79568 145806 79620
rect 145944 79552 145972 79840
rect 146174 79688 146202 79908
rect 146110 79636 146116 79688
rect 146168 79648 146202 79688
rect 146168 79636 146174 79648
rect 145926 79500 145932 79552
rect 145984 79500 145990 79552
rect 146404 79540 146432 80464
rect 148658 80124 151952 80152
rect 146634 79988 146938 80016
rect 146524 79908 146530 79960
rect 146582 79908 146588 79960
rect 146542 79756 146570 79908
rect 146478 79704 146484 79756
rect 146536 79716 146570 79756
rect 146536 79704 146542 79716
rect 146634 79620 146662 79988
rect 146910 79960 146938 79988
rect 147002 79988 147214 80016
rect 146800 79908 146806 79960
rect 146858 79908 146864 79960
rect 146892 79908 146898 79960
rect 146950 79908 146956 79960
rect 146818 79880 146846 79908
rect 147002 79880 147030 79988
rect 147076 79908 147082 79960
rect 147134 79908 147140 79960
rect 146818 79852 147030 79880
rect 147094 79812 147122 79908
rect 146956 79784 147122 79812
rect 146956 79688 146984 79784
rect 147186 79688 147214 79988
rect 148658 79960 148686 80124
rect 150774 79988 151814 80016
rect 150774 79960 150802 79988
rect 147812 79908 147818 79960
rect 147870 79908 147876 79960
rect 147996 79908 148002 79960
rect 148054 79908 148060 79960
rect 148548 79948 148554 79960
rect 148244 79920 148554 79948
rect 147536 79840 147542 79892
rect 147594 79840 147600 79892
rect 146938 79636 146944 79688
rect 146996 79636 147002 79688
rect 147122 79636 147128 79688
rect 147180 79648 147214 79688
rect 147554 79688 147582 79840
rect 147628 79772 147634 79824
rect 147686 79772 147692 79824
rect 147646 79744 147674 79772
rect 147646 79716 147720 79744
rect 147554 79648 147588 79688
rect 147180 79636 147186 79648
rect 147582 79636 147588 79648
rect 147640 79636 147646 79688
rect 146570 79568 146576 79620
rect 146628 79580 146662 79620
rect 146628 79568 146634 79580
rect 146846 79568 146852 79620
rect 146904 79608 146910 79620
rect 147692 79608 147720 79716
rect 146904 79580 147720 79608
rect 147830 79608 147858 79908
rect 148014 79688 148042 79908
rect 148244 79688 148272 79920
rect 148548 79908 148554 79920
rect 148606 79908 148612 79960
rect 148640 79908 148646 79960
rect 148698 79908 148704 79960
rect 149008 79908 149014 79960
rect 149066 79908 149072 79960
rect 149376 79948 149382 79960
rect 149164 79920 149382 79948
rect 148364 79840 148370 79892
rect 148422 79840 148428 79892
rect 148456 79840 148462 79892
rect 148514 79840 148520 79892
rect 148382 79744 148410 79840
rect 148336 79716 148410 79744
rect 147950 79636 147956 79688
rect 148008 79648 148042 79688
rect 148008 79636 148014 79648
rect 148226 79636 148232 79688
rect 148284 79636 148290 79688
rect 148042 79608 148048 79620
rect 147830 79580 148048 79608
rect 146904 79568 146910 79580
rect 148042 79568 148048 79580
rect 148100 79568 148106 79620
rect 147674 79540 147680 79552
rect 146404 79512 147680 79540
rect 147674 79500 147680 79512
rect 147732 79500 147738 79552
rect 148336 79540 148364 79716
rect 148474 79688 148502 79840
rect 148732 79772 148738 79824
rect 148790 79772 148796 79824
rect 148750 79688 148778 79772
rect 149026 79688 149054 79908
rect 149164 79688 149192 79920
rect 149376 79908 149382 79920
rect 149434 79908 149440 79960
rect 149652 79948 149658 79960
rect 149624 79908 149658 79948
rect 149710 79908 149716 79960
rect 149836 79908 149842 79960
rect 149894 79908 149900 79960
rect 150480 79908 150486 79960
rect 150538 79908 150544 79960
rect 150756 79908 150762 79960
rect 150814 79908 150820 79960
rect 150848 79908 150854 79960
rect 150906 79908 150912 79960
rect 150940 79908 150946 79960
rect 150998 79908 151004 79960
rect 151032 79908 151038 79960
rect 151090 79908 151096 79960
rect 151308 79948 151314 79960
rect 151280 79908 151314 79948
rect 151366 79908 151372 79960
rect 149284 79840 149290 79892
rect 149342 79840 149348 79892
rect 148410 79636 148416 79688
rect 148468 79648 148502 79688
rect 148468 79636 148474 79648
rect 148686 79636 148692 79688
rect 148744 79648 148778 79688
rect 148744 79636 148750 79648
rect 148962 79636 148968 79688
rect 149020 79648 149054 79688
rect 149020 79636 149026 79648
rect 149146 79636 149152 79688
rect 149204 79636 149210 79688
rect 149302 79676 149330 79840
rect 149624 79756 149652 79908
rect 149854 79880 149882 79908
rect 149716 79852 149882 79880
rect 149606 79704 149612 79756
rect 149664 79704 149670 79756
rect 149422 79676 149428 79688
rect 149302 79648 149428 79676
rect 149422 79636 149428 79648
rect 149480 79636 149486 79688
rect 149238 79568 149244 79620
rect 149296 79608 149302 79620
rect 149716 79608 149744 79852
rect 149928 79840 149934 79892
rect 149986 79840 149992 79892
rect 150296 79840 150302 79892
rect 150354 79840 150360 79892
rect 149946 79688 149974 79840
rect 150020 79772 150026 79824
rect 150078 79772 150084 79824
rect 149882 79636 149888 79688
rect 149940 79648 149974 79688
rect 149940 79636 149946 79648
rect 150038 79620 150066 79772
rect 150314 79688 150342 79840
rect 150250 79636 150256 79688
rect 150308 79648 150342 79688
rect 150308 79636 150314 79648
rect 149296 79580 149744 79608
rect 149296 79568 149302 79580
rect 149974 79568 149980 79620
rect 150032 79580 150066 79620
rect 150498 79620 150526 79908
rect 150866 79620 150894 79908
rect 150498 79580 150532 79620
rect 150032 79568 150038 79580
rect 150526 79568 150532 79580
rect 150584 79568 150590 79620
rect 150802 79568 150808 79620
rect 150860 79580 150894 79620
rect 150860 79568 150866 79580
rect 150958 79552 150986 79908
rect 151050 79620 151078 79908
rect 151280 79756 151308 79908
rect 151400 79880 151406 79892
rect 151372 79840 151406 79880
rect 151458 79840 151464 79892
rect 151372 79756 151400 79840
rect 151262 79704 151268 79756
rect 151320 79704 151326 79756
rect 151354 79704 151360 79756
rect 151412 79704 151418 79756
rect 151050 79580 151084 79620
rect 151078 79568 151084 79580
rect 151136 79568 151142 79620
rect 148594 79540 148600 79552
rect 148336 79512 148600 79540
rect 148594 79500 148600 79512
rect 148652 79500 148658 79552
rect 150958 79512 150992 79552
rect 150986 79500 150992 79512
rect 151044 79500 151050 79552
rect 151786 79540 151814 79988
rect 151924 79620 151952 80124
rect 152154 80124 153194 80152
rect 152154 79960 152182 80124
rect 153166 80084 153194 80124
rect 153166 80056 155862 80084
rect 152044 79908 152050 79960
rect 152102 79908 152108 79960
rect 152136 79908 152142 79960
rect 152194 79908 152200 79960
rect 152412 79908 152418 79960
rect 152470 79908 152476 79960
rect 152780 79908 152786 79960
rect 152838 79908 152844 79960
rect 152872 79908 152878 79960
rect 152930 79908 152936 79960
rect 152964 79908 152970 79960
rect 153022 79908 153028 79960
rect 153148 79908 153154 79960
rect 153206 79908 153212 79960
rect 153240 79908 153246 79960
rect 153298 79908 153304 79960
rect 153332 79908 153338 79960
rect 153390 79908 153396 79960
rect 153608 79908 153614 79960
rect 153666 79948 153672 79960
rect 154068 79948 154074 79960
rect 153666 79920 153838 79948
rect 153666 79908 153672 79920
rect 152062 79824 152090 79908
rect 152044 79772 152050 79824
rect 152102 79772 152108 79824
rect 152274 79636 152280 79688
rect 152332 79676 152338 79688
rect 152430 79676 152458 79908
rect 152504 79840 152510 79892
rect 152562 79840 152568 79892
rect 152688 79840 152694 79892
rect 152746 79840 152752 79892
rect 152522 79756 152550 79840
rect 152522 79716 152556 79756
rect 152550 79704 152556 79716
rect 152608 79704 152614 79756
rect 152332 79648 152458 79676
rect 152332 79636 152338 79648
rect 152706 79620 152734 79840
rect 152798 79688 152826 79908
rect 152890 79824 152918 79908
rect 152872 79772 152878 79824
rect 152930 79772 152936 79824
rect 152982 79744 153010 79908
rect 153056 79840 153062 79892
rect 153114 79840 153120 79892
rect 152936 79716 153010 79744
rect 152798 79648 152832 79688
rect 152826 79636 152832 79648
rect 152884 79636 152890 79688
rect 151906 79568 151912 79620
rect 151964 79568 151970 79620
rect 152642 79568 152648 79620
rect 152700 79580 152734 79620
rect 152936 79608 152964 79716
rect 153074 79688 153102 79840
rect 153010 79636 153016 79688
rect 153068 79648 153102 79688
rect 153068 79636 153074 79648
rect 152798 79580 152964 79608
rect 152700 79568 152706 79580
rect 152798 79552 152826 79580
rect 152458 79540 152464 79552
rect 151786 79512 152464 79540
rect 152458 79500 152464 79512
rect 152516 79500 152522 79552
rect 152734 79500 152740 79552
rect 152792 79512 152826 79552
rect 152792 79500 152798 79512
rect 152918 79500 152924 79552
rect 152976 79540 152982 79552
rect 153166 79540 153194 79908
rect 152976 79512 153194 79540
rect 153258 79540 153286 79908
rect 153350 79756 153378 79908
rect 153700 79772 153706 79824
rect 153758 79772 153764 79824
rect 153350 79716 153384 79756
rect 153378 79704 153384 79716
rect 153436 79704 153442 79756
rect 153718 79688 153746 79772
rect 153654 79636 153660 79688
rect 153712 79648 153746 79688
rect 153712 79636 153718 79648
rect 153810 79620 153838 79920
rect 154040 79908 154074 79948
rect 154126 79908 154132 79960
rect 154160 79908 154166 79960
rect 154218 79908 154224 79960
rect 154252 79908 154258 79960
rect 154310 79908 154316 79960
rect 154344 79908 154350 79960
rect 154402 79908 154408 79960
rect 154528 79908 154534 79960
rect 154586 79908 154592 79960
rect 154804 79908 154810 79960
rect 154862 79908 154868 79960
rect 154896 79908 154902 79960
rect 154954 79908 154960 79960
rect 155264 79948 155270 79960
rect 155236 79908 155270 79948
rect 155322 79908 155328 79960
rect 155448 79908 155454 79960
rect 155506 79908 155512 79960
rect 155540 79908 155546 79960
rect 155598 79908 155604 79960
rect 153884 79840 153890 79892
rect 153942 79840 153948 79892
rect 153902 79688 153930 79840
rect 154040 79756 154068 79908
rect 154178 79880 154206 79908
rect 154132 79852 154206 79880
rect 154022 79704 154028 79756
rect 154080 79704 154086 79756
rect 153902 79648 153936 79688
rect 153930 79636 153936 79648
rect 153988 79636 153994 79688
rect 153746 79568 153752 79620
rect 153804 79580 153838 79620
rect 153804 79568 153810 79580
rect 153838 79540 153844 79552
rect 153258 79512 153844 79540
rect 152976 79500 152982 79512
rect 153838 79500 153844 79512
rect 153896 79500 153902 79552
rect 154132 79540 154160 79852
rect 154270 79824 154298 79908
rect 154206 79772 154212 79824
rect 154264 79784 154298 79824
rect 154264 79772 154270 79784
rect 154362 79756 154390 79908
rect 154546 79824 154574 79908
rect 154546 79784 154580 79824
rect 154574 79772 154580 79784
rect 154632 79772 154638 79824
rect 154712 79772 154718 79824
rect 154770 79772 154776 79824
rect 154298 79704 154304 79756
rect 154356 79716 154390 79756
rect 154356 79704 154362 79716
rect 154482 79568 154488 79620
rect 154540 79608 154546 79620
rect 154730 79608 154758 79772
rect 154822 79756 154850 79908
rect 154914 79812 154942 79908
rect 155080 79880 155086 79892
rect 155052 79840 155086 79880
rect 155138 79840 155144 79892
rect 154914 79784 154988 79812
rect 154822 79716 154856 79756
rect 154850 79704 154856 79716
rect 154908 79704 154914 79756
rect 154960 79620 154988 79784
rect 155052 79756 155080 79840
rect 155236 79824 155264 79908
rect 155218 79772 155224 79824
rect 155276 79772 155282 79824
rect 155310 79772 155316 79824
rect 155368 79812 155374 79824
rect 155466 79812 155494 79908
rect 155368 79784 155494 79812
rect 155368 79772 155374 79784
rect 155034 79704 155040 79756
rect 155092 79704 155098 79756
rect 155126 79704 155132 79756
rect 155184 79744 155190 79756
rect 155184 79716 155448 79744
rect 155184 79704 155190 79716
rect 155420 79620 155448 79716
rect 155558 79688 155586 79908
rect 155724 79840 155730 79892
rect 155782 79840 155788 79892
rect 155742 79688 155770 79840
rect 155834 79824 155862 80056
rect 156386 80056 158300 80084
rect 155926 79988 156184 80016
rect 155926 79960 155954 79988
rect 155908 79908 155914 79960
rect 155966 79908 155972 79960
rect 156000 79908 156006 79960
rect 156058 79908 156064 79960
rect 155834 79784 155868 79824
rect 155862 79772 155868 79784
rect 155920 79772 155926 79824
rect 155494 79636 155500 79688
rect 155552 79648 155586 79688
rect 155552 79636 155558 79648
rect 155678 79636 155684 79688
rect 155736 79648 155770 79688
rect 155736 79636 155742 79648
rect 156018 79620 156046 79908
rect 154540 79580 154758 79608
rect 154540 79568 154546 79580
rect 154942 79568 154948 79620
rect 155000 79568 155006 79620
rect 155402 79568 155408 79620
rect 155460 79568 155466 79620
rect 155954 79568 155960 79620
rect 156012 79580 156046 79620
rect 156156 79608 156184 79988
rect 156386 79960 156414 80056
rect 156570 79988 156966 80016
rect 156368 79908 156374 79960
rect 156426 79908 156432 79960
rect 156460 79908 156466 79960
rect 156518 79908 156524 79960
rect 156478 79880 156506 79908
rect 156432 79852 156506 79880
rect 156322 79608 156328 79620
rect 156156 79580 156328 79608
rect 156012 79568 156018 79580
rect 156322 79568 156328 79580
rect 156380 79568 156386 79620
rect 155586 79540 155592 79552
rect 154132 79512 155592 79540
rect 155586 79500 155592 79512
rect 155644 79500 155650 79552
rect 156432 79540 156460 79852
rect 156570 79812 156598 79988
rect 156644 79908 156650 79960
rect 156702 79908 156708 79960
rect 156736 79908 156742 79960
rect 156794 79908 156800 79960
rect 156828 79908 156834 79960
rect 156886 79908 156892 79960
rect 156524 79784 156598 79812
rect 156524 79608 156552 79784
rect 156662 79756 156690 79908
rect 156598 79704 156604 79756
rect 156656 79716 156690 79756
rect 156656 79704 156662 79716
rect 156754 79676 156782 79908
rect 156846 79744 156874 79908
rect 156938 79892 156966 79988
rect 157196 79908 157202 79960
rect 157254 79908 157260 79960
rect 157472 79908 157478 79960
rect 157530 79948 157536 79960
rect 157530 79908 157564 79948
rect 157656 79908 157662 79960
rect 157714 79908 157720 79960
rect 157748 79908 157754 79960
rect 157806 79908 157812 79960
rect 157932 79908 157938 79960
rect 157990 79908 157996 79960
rect 156920 79840 156926 79892
rect 156978 79840 156984 79892
rect 157012 79840 157018 79892
rect 157070 79840 157076 79892
rect 157030 79812 157058 79840
rect 157030 79784 157104 79812
rect 156846 79716 157012 79744
rect 156874 79676 156880 79688
rect 156754 79648 156880 79676
rect 156874 79636 156880 79648
rect 156932 79636 156938 79688
rect 156524 79580 156736 79608
rect 156506 79540 156512 79552
rect 156432 79512 156512 79540
rect 156506 79500 156512 79512
rect 156564 79500 156570 79552
rect 156708 79540 156736 79580
rect 156782 79568 156788 79620
rect 156840 79608 156846 79620
rect 156984 79608 157012 79716
rect 157076 79620 157104 79784
rect 157214 79688 157242 79908
rect 157288 79840 157294 79892
rect 157346 79880 157352 79892
rect 157346 79852 157472 79880
rect 157346 79840 157352 79852
rect 157444 79824 157472 79852
rect 157426 79772 157432 79824
rect 157484 79772 157490 79824
rect 157150 79636 157156 79688
rect 157208 79648 157242 79688
rect 157208 79636 157214 79648
rect 157536 79620 157564 79908
rect 157674 79880 157702 79908
rect 157628 79852 157702 79880
rect 156840 79580 157012 79608
rect 156840 79568 156846 79580
rect 157058 79568 157064 79620
rect 157116 79568 157122 79620
rect 157518 79568 157524 79620
rect 157576 79568 157582 79620
rect 156966 79540 156972 79552
rect 156708 79512 156972 79540
rect 156966 79500 156972 79512
rect 157024 79500 157030 79552
rect 157628 79540 157656 79852
rect 157766 79824 157794 79908
rect 157840 79840 157846 79892
rect 157898 79840 157904 79892
rect 157702 79772 157708 79824
rect 157760 79784 157794 79824
rect 157760 79772 157766 79784
rect 157858 79744 157886 79840
rect 157812 79716 157886 79744
rect 157812 79608 157840 79716
rect 157950 79688 157978 79908
rect 158024 79840 158030 79892
rect 158082 79840 158088 79892
rect 158272 79880 158300 80056
rect 158778 79892 158806 80600
rect 174446 80588 174452 80640
rect 174504 80588 174510 80640
rect 174538 80588 174544 80640
rect 174596 80628 174602 80640
rect 176626 80628 176654 80668
rect 580718 80656 580724 80668
rect 580776 80656 580782 80708
rect 174596 80600 176654 80628
rect 174596 80588 174602 80600
rect 178034 80588 178040 80640
rect 178092 80628 178098 80640
rect 580626 80628 580632 80640
rect 178092 80600 580632 80628
rect 178092 80588 178098 80600
rect 580626 80588 580632 80600
rect 580684 80588 580690 80640
rect 174722 80560 174728 80572
rect 168346 80532 174728 80560
rect 168346 80220 168374 80532
rect 174722 80520 174728 80532
rect 174780 80520 174786 80572
rect 174832 80532 178034 80560
rect 174630 80424 174636 80436
rect 161262 80192 168374 80220
rect 168898 80396 174636 80424
rect 158870 79988 160186 80016
rect 158272 79852 158438 79880
rect 158042 79812 158070 79840
rect 158042 79784 158162 79812
rect 158134 79688 158162 79784
rect 158208 79772 158214 79824
rect 158266 79812 158272 79824
rect 158266 79784 158346 79812
rect 158266 79772 158272 79784
rect 157886 79636 157892 79688
rect 157944 79648 157978 79688
rect 157944 79636 157950 79648
rect 158116 79636 158122 79688
rect 158174 79636 158180 79688
rect 157978 79608 157984 79620
rect 157812 79580 157984 79608
rect 157978 79568 157984 79580
rect 158036 79568 158042 79620
rect 158318 79552 158346 79784
rect 158410 79688 158438 79852
rect 158760 79840 158766 79892
rect 158818 79840 158824 79892
rect 158484 79772 158490 79824
rect 158542 79812 158548 79824
rect 158542 79772 158576 79812
rect 158548 79688 158576 79772
rect 158714 79704 158720 79756
rect 158772 79744 158778 79756
rect 158870 79744 158898 79988
rect 159036 79908 159042 79960
rect 159094 79908 159100 79960
rect 159680 79908 159686 79960
rect 159738 79908 159744 79960
rect 158772 79716 158898 79744
rect 158772 79704 158778 79716
rect 158410 79648 158444 79688
rect 158438 79636 158444 79648
rect 158496 79636 158502 79688
rect 158530 79636 158536 79688
rect 158588 79636 158594 79688
rect 158070 79540 158076 79552
rect 157628 79512 158076 79540
rect 158070 79500 158076 79512
rect 158128 79500 158134 79552
rect 158254 79500 158260 79552
rect 158312 79512 158346 79552
rect 159054 79540 159082 79908
rect 159404 79840 159410 79892
rect 159462 79840 159468 79892
rect 159496 79840 159502 79892
rect 159554 79840 159560 79892
rect 159588 79840 159594 79892
rect 159646 79840 159652 79892
rect 159422 79744 159450 79840
rect 159284 79716 159450 79744
rect 159284 79608 159312 79716
rect 159358 79636 159364 79688
rect 159416 79676 159422 79688
rect 159514 79676 159542 79840
rect 159416 79648 159542 79676
rect 159416 79636 159422 79648
rect 159606 79620 159634 79840
rect 159450 79608 159456 79620
rect 159284 79580 159456 79608
rect 159450 79568 159456 79580
rect 159508 79568 159514 79620
rect 159542 79568 159548 79620
rect 159600 79580 159634 79620
rect 159600 79568 159606 79580
rect 159358 79540 159364 79552
rect 159054 79512 159364 79540
rect 158312 79500 158318 79512
rect 159358 79500 159364 79512
rect 159416 79500 159422 79552
rect 159698 79540 159726 79908
rect 160158 79892 160186 79988
rect 160802 79988 161014 80016
rect 160692 79948 160698 79960
rect 160572 79920 160698 79948
rect 160048 79840 160054 79892
rect 160106 79840 160112 79892
rect 160140 79840 160146 79892
rect 160198 79840 160204 79892
rect 160416 79840 160422 79892
rect 160474 79880 160480 79892
rect 160474 79840 160508 79880
rect 159864 79772 159870 79824
rect 159922 79772 159928 79824
rect 159882 79744 159910 79772
rect 159836 79716 159910 79744
rect 159836 79688 159864 79716
rect 159818 79636 159824 79688
rect 159876 79636 159882 79688
rect 159910 79636 159916 79688
rect 159968 79676 159974 79688
rect 160066 79676 160094 79840
rect 160480 79756 160508 79840
rect 160462 79704 160468 79756
rect 160520 79704 160526 79756
rect 159968 79648 160094 79676
rect 159968 79636 159974 79648
rect 160572 79620 160600 79920
rect 160692 79908 160698 79920
rect 160750 79908 160756 79960
rect 160802 79620 160830 79988
rect 160986 79960 161014 79988
rect 160876 79908 160882 79960
rect 160934 79908 160940 79960
rect 160968 79908 160974 79960
rect 161026 79908 161032 79960
rect 160894 79880 160922 79908
rect 161152 79880 161158 79892
rect 160894 79852 160968 79880
rect 160940 79676 160968 79852
rect 161124 79840 161158 79880
rect 161210 79840 161216 79892
rect 161124 79756 161152 79840
rect 161262 79756 161290 80192
rect 168898 80152 168926 80396
rect 174630 80384 174636 80396
rect 174688 80384 174694 80436
rect 174832 80288 174860 80532
rect 178006 80424 178034 80532
rect 178006 80396 180794 80424
rect 180766 80356 180794 80396
rect 554774 80356 554780 80368
rect 180766 80328 554780 80356
rect 554774 80316 554780 80328
rect 554832 80316 554838 80368
rect 164298 80124 168926 80152
rect 168990 80260 174860 80288
rect 161354 79988 161612 80016
rect 161354 79960 161382 79988
rect 161336 79908 161342 79960
rect 161394 79908 161400 79960
rect 161428 79908 161434 79960
rect 161486 79908 161492 79960
rect 161106 79704 161112 79756
rect 161164 79704 161170 79756
rect 161198 79704 161204 79756
rect 161256 79716 161290 79756
rect 161256 79704 161262 79716
rect 161014 79676 161020 79688
rect 160940 79648 161020 79676
rect 161014 79636 161020 79648
rect 161072 79636 161078 79688
rect 160554 79568 160560 79620
rect 160612 79568 160618 79620
rect 160738 79568 160744 79620
rect 160796 79580 160830 79620
rect 160796 79568 160802 79580
rect 161446 79552 161474 79908
rect 161584 79688 161612 79988
rect 162734 79988 163406 80016
rect 161796 79908 161802 79960
rect 161854 79908 161860 79960
rect 162164 79948 162170 79960
rect 161998 79920 162170 79948
rect 161814 79744 161842 79908
rect 161888 79772 161894 79824
rect 161946 79772 161952 79824
rect 161676 79716 161842 79744
rect 161566 79636 161572 79688
rect 161624 79636 161630 79688
rect 160646 79540 160652 79552
rect 159698 79512 160652 79540
rect 160646 79500 160652 79512
rect 160704 79500 160710 79552
rect 161382 79500 161388 79552
rect 161440 79512 161474 79552
rect 161440 79500 161446 79512
rect 161676 79484 161704 79716
rect 161906 79688 161934 79772
rect 161842 79636 161848 79688
rect 161900 79648 161934 79688
rect 161900 79636 161906 79648
rect 161998 79608 162026 79920
rect 162164 79908 162170 79920
rect 162222 79908 162228 79960
rect 162624 79908 162630 79960
rect 162682 79908 162688 79960
rect 162072 79840 162078 79892
rect 162130 79840 162136 79892
rect 162256 79840 162262 79892
rect 162314 79840 162320 79892
rect 161860 79580 162026 79608
rect 144086 79432 144092 79484
rect 144144 79472 144150 79484
rect 161566 79472 161572 79484
rect 144144 79444 161572 79472
rect 144144 79432 144150 79444
rect 161566 79432 161572 79444
rect 161624 79432 161630 79484
rect 161658 79432 161664 79484
rect 161716 79432 161722 79484
rect 161860 79472 161888 79580
rect 161934 79500 161940 79552
rect 161992 79540 161998 79552
rect 162090 79540 162118 79840
rect 161992 79512 162118 79540
rect 161992 79500 161998 79512
rect 162118 79472 162124 79484
rect 161860 79444 162124 79472
rect 162118 79432 162124 79444
rect 162176 79432 162182 79484
rect 162274 79472 162302 79840
rect 162440 79812 162446 79824
rect 162412 79772 162446 79812
rect 162498 79772 162504 79824
rect 162412 79620 162440 79772
rect 162642 79688 162670 79908
rect 162734 79744 162762 79988
rect 163378 79960 163406 79988
rect 164298 79960 164326 80124
rect 168990 80016 169018 80260
rect 174906 80248 174912 80300
rect 174964 80288 174970 80300
rect 252554 80288 252560 80300
rect 174964 80260 252560 80288
rect 174964 80248 174970 80260
rect 252554 80248 252560 80260
rect 252612 80248 252618 80300
rect 174722 80180 174728 80232
rect 174780 80220 174786 80232
rect 320174 80220 320180 80232
rect 174780 80192 320180 80220
rect 174780 80180 174786 80192
rect 320174 80180 320180 80192
rect 320232 80180 320238 80232
rect 171566 80124 174078 80152
rect 165678 79988 167546 80016
rect 165678 79960 165706 79988
rect 163360 79908 163366 79960
rect 163418 79908 163424 79960
rect 163636 79908 163642 79960
rect 163694 79908 163700 79960
rect 163728 79908 163734 79960
rect 163786 79908 163792 79960
rect 164280 79908 164286 79960
rect 164338 79908 164344 79960
rect 164556 79908 164562 79960
rect 164614 79908 164620 79960
rect 164740 79908 164746 79960
rect 164798 79908 164804 79960
rect 165384 79948 165390 79960
rect 165034 79920 165390 79948
rect 163176 79880 163182 79892
rect 163148 79840 163182 79880
rect 163234 79840 163240 79892
rect 162734 79716 162808 79744
rect 162780 79688 162808 79716
rect 162642 79648 162676 79688
rect 162670 79636 162676 79648
rect 162728 79636 162734 79688
rect 162762 79636 162768 79688
rect 162820 79636 162826 79688
rect 162394 79568 162400 79620
rect 162452 79568 162458 79620
rect 163148 79608 163176 79840
rect 163268 79812 163274 79824
rect 163240 79772 163274 79812
rect 163326 79772 163332 79824
rect 163544 79772 163550 79824
rect 163602 79772 163608 79824
rect 163240 79688 163268 79772
rect 163222 79636 163228 79688
rect 163280 79636 163286 79688
rect 163314 79636 163320 79688
rect 163372 79676 163378 79688
rect 163562 79676 163590 79772
rect 163372 79648 163590 79676
rect 163654 79676 163682 79908
rect 163746 79756 163774 79908
rect 163820 79840 163826 79892
rect 163878 79880 163884 79892
rect 163878 79840 163912 79880
rect 164188 79840 164194 79892
rect 164246 79840 164252 79892
rect 163746 79716 163780 79756
rect 163774 79704 163780 79716
rect 163832 79704 163838 79756
rect 163884 79688 163912 79840
rect 163654 79648 163820 79676
rect 163372 79636 163378 79648
rect 163590 79608 163596 79620
rect 163148 79580 163596 79608
rect 163590 79568 163596 79580
rect 163648 79568 163654 79620
rect 163792 79608 163820 79648
rect 163866 79636 163872 79688
rect 163924 79636 163930 79688
rect 164206 79676 164234 79840
rect 164418 79676 164424 79688
rect 164206 79648 164424 79676
rect 164418 79636 164424 79648
rect 164476 79636 164482 79688
rect 164142 79608 164148 79620
rect 163792 79580 164148 79608
rect 164142 79568 164148 79580
rect 164200 79568 164206 79620
rect 164574 79608 164602 79908
rect 164758 79756 164786 79908
rect 164924 79772 164930 79824
rect 164982 79772 164988 79824
rect 164694 79704 164700 79756
rect 164752 79716 164786 79756
rect 164752 79704 164758 79716
rect 164942 79688 164970 79772
rect 164878 79636 164884 79688
rect 164936 79648 164970 79688
rect 164936 79636 164942 79648
rect 165034 79620 165062 79920
rect 165384 79908 165390 79920
rect 165442 79908 165448 79960
rect 165476 79908 165482 79960
rect 165534 79908 165540 79960
rect 165660 79908 165666 79960
rect 165718 79908 165724 79960
rect 165844 79908 165850 79960
rect 165902 79908 165908 79960
rect 166028 79908 166034 79960
rect 166086 79908 166092 79960
rect 167408 79908 167414 79960
rect 167466 79908 167472 79960
rect 165108 79840 165114 79892
rect 165166 79840 165172 79892
rect 165292 79840 165298 79892
rect 165350 79840 165356 79892
rect 164252 79580 164602 79608
rect 164050 79500 164056 79552
rect 164108 79540 164114 79552
rect 164252 79540 164280 79580
rect 164970 79568 164976 79620
rect 165028 79580 165062 79620
rect 165126 79620 165154 79840
rect 165200 79772 165206 79824
rect 165258 79772 165264 79824
rect 165218 79688 165246 79772
rect 165310 79744 165338 79840
rect 165494 79824 165522 79908
rect 165476 79772 165482 79824
rect 165534 79772 165540 79824
rect 165706 79772 165712 79824
rect 165764 79812 165770 79824
rect 165862 79812 165890 79908
rect 165764 79784 165890 79812
rect 165764 79772 165770 79784
rect 166046 79744 166074 79908
rect 166856 79880 166862 79892
rect 166828 79840 166862 79880
rect 166914 79840 166920 79892
rect 166120 79772 166126 79824
rect 166178 79772 166184 79824
rect 166304 79772 166310 79824
rect 166362 79772 166368 79824
rect 165310 79716 165476 79744
rect 165218 79648 165252 79688
rect 165246 79636 165252 79648
rect 165304 79636 165310 79688
rect 165448 79620 165476 79716
rect 165540 79716 166074 79744
rect 165540 79688 165568 79716
rect 165522 79636 165528 79688
rect 165580 79636 165586 79688
rect 165890 79636 165896 79688
rect 165948 79676 165954 79688
rect 166138 79676 166166 79772
rect 165948 79648 166166 79676
rect 166322 79676 166350 79772
rect 166534 79676 166540 79688
rect 166322 79648 166540 79676
rect 165948 79636 165954 79648
rect 166534 79636 166540 79648
rect 166592 79636 166598 79688
rect 166828 79620 166856 79840
rect 167224 79772 167230 79824
rect 167282 79772 167288 79824
rect 167242 79688 167270 79772
rect 167242 79648 167276 79688
rect 167270 79636 167276 79648
rect 167328 79636 167334 79688
rect 167426 79620 167454 79908
rect 167518 79676 167546 79988
rect 168760 79988 169018 80016
rect 169082 79988 171502 80016
rect 168760 79960 168788 79988
rect 168236 79908 168242 79960
rect 168294 79908 168300 79960
rect 168696 79908 168702 79960
rect 168754 79920 168788 79960
rect 168754 79908 168760 79920
rect 168880 79908 168886 79960
rect 168938 79948 168944 79960
rect 168938 79920 169018 79948
rect 168938 79908 168944 79920
rect 167592 79840 167598 79892
rect 167650 79880 167656 79892
rect 168254 79880 168282 79908
rect 167650 79852 168144 79880
rect 167650 79840 167656 79852
rect 167868 79772 167874 79824
rect 167926 79772 167932 79824
rect 167886 79688 167914 79772
rect 167518 79648 167776 79676
rect 165126 79580 165160 79620
rect 165028 79568 165034 79580
rect 165154 79568 165160 79580
rect 165212 79568 165218 79620
rect 165430 79568 165436 79620
rect 165488 79568 165494 79620
rect 166810 79568 166816 79620
rect 166868 79568 166874 79620
rect 167426 79580 167460 79620
rect 167454 79568 167460 79580
rect 167512 79568 167518 79620
rect 167748 79608 167776 79648
rect 167822 79636 167828 79688
rect 167880 79648 167914 79688
rect 168116 79676 168144 79852
rect 168208 79852 168282 79880
rect 168208 79824 168236 79852
rect 168190 79772 168196 79824
rect 168248 79772 168254 79824
rect 168990 79744 169018 79920
rect 168392 79716 169018 79744
rect 168392 79688 168420 79716
rect 168282 79676 168288 79688
rect 168116 79648 168288 79676
rect 167880 79636 167886 79648
rect 168282 79636 168288 79648
rect 168340 79636 168346 79688
rect 168374 79636 168380 79688
rect 168432 79636 168438 79688
rect 169082 79676 169110 79988
rect 169984 79908 169990 79960
rect 170042 79908 170048 79960
rect 170076 79908 170082 79960
rect 170134 79908 170140 79960
rect 170168 79908 170174 79960
rect 170226 79908 170232 79960
rect 170352 79908 170358 79960
rect 170410 79908 170416 79960
rect 170904 79948 170910 79960
rect 170462 79920 170910 79948
rect 169156 79840 169162 79892
rect 169214 79840 169220 79892
rect 169524 79840 169530 79892
rect 169582 79840 169588 79892
rect 169616 79840 169622 79892
rect 169674 79840 169680 79892
rect 170002 79880 170030 79908
rect 169956 79852 170030 79880
rect 169036 79648 169110 79676
rect 169036 79608 169064 79648
rect 169174 79620 169202 79840
rect 169340 79812 169346 79824
rect 169312 79772 169346 79812
rect 169398 79772 169404 79824
rect 169432 79772 169438 79824
rect 169490 79772 169496 79824
rect 169312 79620 169340 79772
rect 169450 79744 169478 79772
rect 169404 79716 169478 79744
rect 169404 79688 169432 79716
rect 169542 79688 169570 79840
rect 169386 79636 169392 79688
rect 169444 79636 169450 79688
rect 169478 79636 169484 79688
rect 169536 79648 169570 79688
rect 169634 79688 169662 79840
rect 169634 79648 169668 79688
rect 169536 79636 169542 79648
rect 169662 79636 169668 79648
rect 169720 79636 169726 79688
rect 169956 79676 169984 79852
rect 170094 79756 170122 79908
rect 170186 79812 170214 79908
rect 170186 79784 170260 79812
rect 170094 79716 170128 79756
rect 170122 79704 170128 79716
rect 170180 79704 170186 79756
rect 170232 79688 170260 79784
rect 170370 79688 170398 79908
rect 170030 79676 170036 79688
rect 169956 79648 170036 79676
rect 170030 79636 170036 79648
rect 170088 79636 170094 79688
rect 170214 79636 170220 79688
rect 170272 79636 170278 79688
rect 170306 79636 170312 79688
rect 170364 79648 170398 79688
rect 170364 79636 170370 79648
rect 167748 79580 169064 79608
rect 169110 79568 169116 79620
rect 169168 79580 169202 79620
rect 169168 79568 169174 79580
rect 169294 79568 169300 79620
rect 169352 79568 169358 79620
rect 169570 79568 169576 79620
rect 169628 79608 169634 79620
rect 169628 79580 170168 79608
rect 169628 79568 169634 79580
rect 164108 79512 164280 79540
rect 164108 79500 164114 79512
rect 164418 79500 164424 79552
rect 164476 79540 164482 79552
rect 164476 79512 170076 79540
rect 164476 79500 164482 79512
rect 162486 79472 162492 79484
rect 162274 79444 162492 79472
rect 162486 79432 162492 79444
rect 162544 79432 162550 79484
rect 169570 79432 169576 79484
rect 169628 79432 169634 79484
rect 141200 79376 141924 79404
rect 141200 79364 141206 79376
rect 143534 79364 143540 79416
rect 143592 79404 143598 79416
rect 159082 79404 159088 79416
rect 143592 79376 159088 79404
rect 143592 79364 143598 79376
rect 159082 79364 159088 79376
rect 159140 79364 159146 79416
rect 160250 79376 160508 79404
rect 126532 79308 135254 79336
rect 126532 79200 126560 79308
rect 137278 79296 137284 79348
rect 137336 79336 137342 79348
rect 137336 79308 142844 79336
rect 137336 79296 137342 79308
rect 126974 79228 126980 79280
rect 127032 79268 127038 79280
rect 140774 79268 140780 79280
rect 127032 79240 140780 79268
rect 127032 79228 127038 79240
rect 140774 79228 140780 79240
rect 140832 79228 140838 79280
rect 142816 79268 142844 79308
rect 142890 79296 142896 79348
rect 142948 79336 142954 79348
rect 160250 79336 160278 79376
rect 142948 79308 160278 79336
rect 160480 79336 160508 79376
rect 161290 79364 161296 79416
rect 161348 79404 161354 79416
rect 169588 79404 169616 79432
rect 161348 79376 169616 79404
rect 161348 79364 161354 79376
rect 169938 79336 169944 79348
rect 160480 79308 169944 79336
rect 142948 79296 142954 79308
rect 169938 79296 169944 79308
rect 169996 79296 170002 79348
rect 170048 79336 170076 79512
rect 170140 79404 170168 79580
rect 170462 79472 170490 79920
rect 170904 79908 170910 79920
rect 170962 79908 170968 79960
rect 170536 79840 170542 79892
rect 170594 79840 170600 79892
rect 170720 79840 170726 79892
rect 170778 79880 170784 79892
rect 170778 79852 171226 79880
rect 170778 79840 170784 79852
rect 170554 79688 170582 79840
rect 170996 79772 171002 79824
rect 171054 79772 171060 79824
rect 171014 79688 171042 79772
rect 170554 79648 170588 79688
rect 170582 79636 170588 79648
rect 170640 79636 170646 79688
rect 171014 79648 171048 79688
rect 171042 79636 171048 79648
rect 171100 79636 171106 79688
rect 171198 79676 171226 79852
rect 171364 79840 171370 79892
rect 171422 79840 171428 79892
rect 171474 79880 171502 79988
rect 171566 79960 171594 80124
rect 174050 80084 174078 80124
rect 174446 80112 174452 80164
rect 174504 80152 174510 80164
rect 426434 80152 426440 80164
rect 174504 80124 426440 80152
rect 174504 80112 174510 80124
rect 426434 80112 426440 80124
rect 426492 80112 426498 80164
rect 177390 80084 177396 80096
rect 172164 80056 173710 80084
rect 174050 80056 177396 80084
rect 171548 79908 171554 79960
rect 171606 79908 171612 79960
rect 172164 79880 172192 80056
rect 171474 79852 172192 79880
rect 172256 79988 172882 80016
rect 171382 79812 171410 79840
rect 172100 79812 172106 79824
rect 171382 79784 171548 79812
rect 171410 79676 171416 79688
rect 171198 79648 171416 79676
rect 171410 79636 171416 79648
rect 171468 79636 171474 79688
rect 171226 79568 171232 79620
rect 171284 79608 171290 79620
rect 171520 79608 171548 79784
rect 171284 79580 171548 79608
rect 171612 79784 172106 79812
rect 171612 79608 171640 79784
rect 172100 79772 172106 79784
rect 172158 79772 172164 79824
rect 171686 79636 171692 79688
rect 171744 79676 171750 79688
rect 172256 79676 172284 79988
rect 172854 79960 172882 79988
rect 172744 79908 172750 79960
rect 172802 79908 172808 79960
rect 172836 79908 172842 79960
rect 172894 79908 172900 79960
rect 173296 79908 173302 79960
rect 173354 79908 173360 79960
rect 173388 79908 173394 79960
rect 173446 79908 173452 79960
rect 173572 79908 173578 79960
rect 173630 79908 173636 79960
rect 171744 79648 172284 79676
rect 171744 79636 171750 79648
rect 172054 79608 172060 79620
rect 171612 79580 172060 79608
rect 171284 79568 171290 79580
rect 172054 79568 172060 79580
rect 172112 79568 172118 79620
rect 172606 79568 172612 79620
rect 172664 79608 172670 79620
rect 172762 79608 172790 79908
rect 172928 79880 172934 79892
rect 172854 79852 172934 79880
rect 172854 79744 172882 79852
rect 172928 79840 172934 79852
rect 172986 79840 172992 79892
rect 173020 79840 173026 79892
rect 173078 79880 173084 79892
rect 173078 79852 173204 79880
rect 173078 79840 173084 79852
rect 172974 79744 172980 79756
rect 172854 79716 172980 79744
rect 172974 79704 172980 79716
rect 173032 79704 173038 79756
rect 172664 79580 172790 79608
rect 172664 79568 172670 79580
rect 172882 79568 172888 79620
rect 172940 79608 172946 79620
rect 173176 79608 173204 79852
rect 173314 79756 173342 79908
rect 173296 79704 173302 79756
rect 173354 79704 173360 79756
rect 173406 79676 173434 79908
rect 173480 79840 173486 79892
rect 173538 79840 173544 79892
rect 173360 79648 173434 79676
rect 173360 79620 173388 79648
rect 173498 79620 173526 79840
rect 173590 79744 173618 79908
rect 173682 79880 173710 80056
rect 177390 80044 177396 80056
rect 177448 80044 177454 80096
rect 182174 80044 182180 80096
rect 182232 80084 182238 80096
rect 184198 80084 184204 80096
rect 182232 80056 184204 80084
rect 182232 80044 182238 80056
rect 184198 80044 184204 80056
rect 184256 80044 184262 80096
rect 174124 79908 174130 79960
rect 174182 79948 174188 79960
rect 174354 79948 174360 79960
rect 174182 79920 174360 79948
rect 174182 79908 174188 79920
rect 174354 79908 174360 79920
rect 174412 79908 174418 79960
rect 174630 79908 174636 79960
rect 174688 79948 174694 79960
rect 174688 79920 181576 79948
rect 174688 79908 174694 79920
rect 181548 79880 181576 79920
rect 498194 79880 498200 79892
rect 173682 79852 180794 79880
rect 181548 79852 498200 79880
rect 173848 79772 173854 79824
rect 173906 79812 173912 79824
rect 174446 79812 174452 79824
rect 173906 79784 174452 79812
rect 173906 79772 173912 79784
rect 174446 79772 174452 79784
rect 174504 79772 174510 79824
rect 180766 79812 180794 79852
rect 498194 79840 498200 79852
rect 498252 79840 498258 79892
rect 514754 79812 514760 79824
rect 180766 79784 514760 79812
rect 514754 79772 514760 79784
rect 514812 79772 514818 79824
rect 173756 79744 173762 79756
rect 173590 79716 173762 79744
rect 173756 79704 173762 79716
rect 173814 79704 173820 79756
rect 180150 79676 180156 79688
rect 172940 79580 173204 79608
rect 172940 79568 172946 79580
rect 173342 79568 173348 79620
rect 173400 79568 173406 79620
rect 173434 79568 173440 79620
rect 173492 79580 173526 79620
rect 173728 79648 180156 79676
rect 173492 79568 173498 79580
rect 170766 79500 170772 79552
rect 170824 79540 170830 79552
rect 173618 79540 173624 79552
rect 170824 79512 173624 79540
rect 170824 79500 170830 79512
rect 173618 79500 173624 79512
rect 173676 79500 173682 79552
rect 170858 79472 170864 79484
rect 170462 79444 170864 79472
rect 170858 79432 170864 79444
rect 170916 79432 170922 79484
rect 171134 79432 171140 79484
rect 171192 79472 171198 79484
rect 173728 79472 173756 79648
rect 180150 79636 180156 79648
rect 180208 79636 180214 79688
rect 171192 79444 173756 79472
rect 171192 79432 171198 79444
rect 170140 79376 171088 79404
rect 170766 79336 170772 79348
rect 170048 79308 170772 79336
rect 170766 79296 170772 79308
rect 170824 79296 170830 79348
rect 171060 79336 171088 79376
rect 171778 79364 171784 79416
rect 171836 79404 171842 79416
rect 181438 79404 181444 79416
rect 171836 79376 181444 79404
rect 171836 79364 171842 79376
rect 181438 79364 181444 79376
rect 181496 79364 181502 79416
rect 184934 79364 184940 79416
rect 184992 79404 184998 79416
rect 580350 79404 580356 79416
rect 184992 79376 580356 79404
rect 184992 79364 184998 79376
rect 580350 79364 580356 79376
rect 580408 79364 580414 79416
rect 174354 79336 174360 79348
rect 171060 79308 174360 79336
rect 174354 79296 174360 79308
rect 174412 79296 174418 79348
rect 177390 79296 177396 79348
rect 177448 79336 177454 79348
rect 580902 79336 580908 79348
rect 177448 79308 580908 79336
rect 177448 79296 177454 79308
rect 580902 79296 580908 79308
rect 580960 79296 580966 79348
rect 146662 79268 146668 79280
rect 142816 79240 146668 79268
rect 146662 79228 146668 79240
rect 146720 79228 146726 79280
rect 147674 79228 147680 79280
rect 147732 79268 147738 79280
rect 157794 79268 157800 79280
rect 147732 79240 157800 79268
rect 147732 79228 147738 79240
rect 157794 79228 157800 79240
rect 157852 79228 157858 79280
rect 161566 79228 161572 79280
rect 161624 79268 161630 79280
rect 164418 79268 164424 79280
rect 161624 79240 164424 79268
rect 161624 79228 161630 79240
rect 164418 79228 164424 79240
rect 164476 79228 164482 79280
rect 164694 79228 164700 79280
rect 164752 79268 164758 79280
rect 164752 79240 171180 79268
rect 164752 79228 164758 79240
rect 126072 79172 126560 79200
rect 128630 79160 128636 79212
rect 128688 79200 128694 79212
rect 128906 79200 128912 79212
rect 128688 79172 128912 79200
rect 128688 79160 128694 79172
rect 128906 79160 128912 79172
rect 128964 79160 128970 79212
rect 128998 79160 129004 79212
rect 129056 79200 129062 79212
rect 130838 79200 130844 79212
rect 129056 79172 130844 79200
rect 129056 79160 129062 79172
rect 130838 79160 130844 79172
rect 130896 79160 130902 79212
rect 131022 79160 131028 79212
rect 131080 79200 131086 79212
rect 134334 79200 134340 79212
rect 131080 79172 134340 79200
rect 131080 79160 131086 79172
rect 134334 79160 134340 79172
rect 134392 79160 134398 79212
rect 135162 79160 135168 79212
rect 135220 79200 135226 79212
rect 170398 79200 170404 79212
rect 135220 79172 170404 79200
rect 135220 79160 135226 79172
rect 170398 79160 170404 79172
rect 170456 79160 170462 79212
rect 171152 79200 171180 79240
rect 171226 79228 171232 79280
rect 171284 79268 171290 79280
rect 174078 79268 174084 79280
rect 171284 79240 174084 79268
rect 171284 79228 171290 79240
rect 174078 79228 174084 79240
rect 174136 79228 174142 79280
rect 174262 79228 174268 79280
rect 174320 79268 174326 79280
rect 288434 79268 288440 79280
rect 174320 79240 288440 79268
rect 174320 79228 174326 79240
rect 288434 79228 288440 79240
rect 288492 79228 288498 79280
rect 173986 79200 173992 79212
rect 171152 79172 173992 79200
rect 173986 79160 173992 79172
rect 174044 79160 174050 79212
rect 125962 79092 125968 79144
rect 126020 79132 126026 79144
rect 126238 79132 126244 79144
rect 126020 79104 126244 79132
rect 126020 79092 126026 79104
rect 126238 79092 126244 79104
rect 126296 79092 126302 79144
rect 127250 79092 127256 79144
rect 127308 79132 127314 79144
rect 137278 79132 137284 79144
rect 127308 79104 137284 79132
rect 127308 79092 127314 79104
rect 137278 79092 137284 79104
rect 137336 79092 137342 79144
rect 140774 79092 140780 79144
rect 140832 79132 140838 79144
rect 142890 79132 142896 79144
rect 140832 79104 142896 79132
rect 140832 79092 140838 79104
rect 142890 79092 142896 79104
rect 142948 79092 142954 79144
rect 146662 79092 146668 79144
rect 146720 79132 146726 79144
rect 146720 79104 157334 79132
rect 146720 79092 146726 79104
rect 126974 79064 126980 79076
rect 125658 79036 126980 79064
rect 126974 79024 126980 79036
rect 127032 79024 127038 79076
rect 139118 79024 139124 79076
rect 139176 79064 139182 79076
rect 143534 79064 143540 79076
rect 139176 79036 143540 79064
rect 139176 79024 139182 79036
rect 143534 79024 143540 79036
rect 143592 79024 143598 79076
rect 157306 79064 157334 79104
rect 158346 79092 158352 79144
rect 158404 79132 158410 79144
rect 161198 79132 161204 79144
rect 158404 79104 161204 79132
rect 158404 79092 158410 79104
rect 161198 79092 161204 79104
rect 161256 79092 161262 79144
rect 161566 79092 161572 79144
rect 161624 79132 161630 79144
rect 161934 79132 161940 79144
rect 161624 79104 161940 79132
rect 161624 79092 161630 79104
rect 161934 79092 161940 79104
rect 161992 79092 161998 79144
rect 162210 79092 162216 79144
rect 162268 79132 162274 79144
rect 324314 79132 324320 79144
rect 162268 79104 324320 79132
rect 162268 79092 162274 79104
rect 324314 79092 324320 79104
rect 324372 79092 324378 79144
rect 158806 79064 158812 79076
rect 157306 79036 158812 79064
rect 158806 79024 158812 79036
rect 158864 79024 158870 79076
rect 159358 79024 159364 79076
rect 159416 79064 159422 79076
rect 164694 79064 164700 79076
rect 159416 79036 164700 79064
rect 159416 79024 159422 79036
rect 164694 79024 164700 79036
rect 164752 79024 164758 79076
rect 172422 79064 172428 79076
rect 166966 79036 172428 79064
rect 135162 78996 135168 79008
rect 125566 78968 135168 78996
rect 135162 78956 135168 78968
rect 135220 78956 135226 79008
rect 144086 78996 144092 79008
rect 137296 78968 144092 78996
rect 125594 78888 125600 78940
rect 125652 78928 125658 78940
rect 127250 78928 127256 78940
rect 125652 78900 127256 78928
rect 125652 78888 125658 78900
rect 127250 78888 127256 78900
rect 127308 78888 127314 78940
rect 132678 78888 132684 78940
rect 132736 78928 132742 78940
rect 132736 78900 133368 78928
rect 132736 78888 132742 78900
rect 133340 78860 133368 78900
rect 137296 78860 137324 78968
rect 144086 78956 144092 78968
rect 144144 78956 144150 79008
rect 150434 78956 150440 79008
rect 150492 78996 150498 79008
rect 150894 78996 150900 79008
rect 150492 78968 150900 78996
rect 150492 78956 150498 78968
rect 150894 78956 150900 78968
rect 150952 78956 150958 79008
rect 157794 78956 157800 79008
rect 157852 78996 157858 79008
rect 166258 78996 166264 79008
rect 157852 78968 166264 78996
rect 157852 78956 157858 78968
rect 166258 78956 166264 78968
rect 166316 78956 166322 79008
rect 150986 78888 150992 78940
rect 151044 78888 151050 78940
rect 158806 78888 158812 78940
rect 158864 78928 158870 78940
rect 159358 78928 159364 78940
rect 158864 78900 159364 78928
rect 158864 78888 158870 78900
rect 159358 78888 159364 78900
rect 159416 78888 159422 78940
rect 166966 78928 166994 79036
rect 172422 79024 172428 79036
rect 172480 79024 172486 79076
rect 172698 79024 172704 79076
rect 172756 79064 172762 79076
rect 293954 79064 293960 79076
rect 172756 79036 293960 79064
rect 172756 79024 172762 79036
rect 293954 79024 293960 79036
rect 294012 79024 294018 79076
rect 167362 78956 167368 79008
rect 167420 78996 167426 79008
rect 167730 78996 167736 79008
rect 167420 78968 167736 78996
rect 167420 78956 167426 78968
rect 167730 78956 167736 78968
rect 167788 78956 167794 79008
rect 169294 78956 169300 79008
rect 169352 78996 169358 79008
rect 169662 78996 169668 79008
rect 169352 78968 169668 78996
rect 169352 78956 169358 78968
rect 169662 78956 169668 78968
rect 169720 78956 169726 79008
rect 172514 78956 172520 79008
rect 172572 78996 172578 79008
rect 367738 78996 367744 79008
rect 172572 78968 367744 78996
rect 172572 78956 172578 78968
rect 367738 78956 367744 78968
rect 367796 78956 367802 79008
rect 172790 78928 172796 78940
rect 159468 78900 166994 78928
rect 167058 78900 172796 78928
rect 133340 78832 137324 78860
rect 133598 78752 133604 78804
rect 133656 78752 133662 78804
rect 138014 78752 138020 78804
rect 138072 78752 138078 78804
rect 138106 78752 138112 78804
rect 138164 78792 138170 78804
rect 138382 78792 138388 78804
rect 138164 78764 138388 78792
rect 138164 78752 138170 78764
rect 138382 78752 138388 78764
rect 138440 78752 138446 78804
rect 140314 78752 140320 78804
rect 140372 78792 140378 78804
rect 140774 78792 140780 78804
rect 140372 78764 140780 78792
rect 140372 78752 140378 78764
rect 140774 78752 140780 78764
rect 140832 78752 140838 78804
rect 132678 78684 132684 78736
rect 132736 78724 132742 78736
rect 132954 78724 132960 78736
rect 132736 78696 132960 78724
rect 132736 78684 132742 78696
rect 132954 78684 132960 78696
rect 133012 78684 133018 78736
rect 133414 78656 133420 78668
rect 125566 78628 133420 78656
rect 125042 78548 125048 78600
rect 125100 78588 125106 78600
rect 125566 78588 125594 78628
rect 133414 78616 133420 78628
rect 133472 78616 133478 78668
rect 125100 78560 125594 78588
rect 125100 78548 125106 78560
rect 125410 78412 125416 78464
rect 125468 78452 125474 78464
rect 133046 78452 133052 78464
rect 125468 78424 133052 78452
rect 125468 78412 125474 78424
rect 133046 78412 133052 78424
rect 133104 78412 133110 78464
rect 133506 78412 133512 78464
rect 133564 78452 133570 78464
rect 133616 78452 133644 78752
rect 138032 78656 138060 78752
rect 146662 78684 146668 78736
rect 146720 78724 146726 78736
rect 147030 78724 147036 78736
rect 146720 78696 147036 78724
rect 146720 78684 146726 78696
rect 147030 78684 147036 78696
rect 147088 78684 147094 78736
rect 138382 78656 138388 78668
rect 138032 78628 138388 78656
rect 138382 78616 138388 78628
rect 138440 78616 138446 78668
rect 139946 78616 139952 78668
rect 140004 78656 140010 78668
rect 140314 78656 140320 78668
rect 140004 78628 140320 78656
rect 140004 78616 140010 78628
rect 140314 78616 140320 78628
rect 140372 78616 140378 78668
rect 146478 78616 146484 78668
rect 146536 78656 146542 78668
rect 147214 78656 147220 78668
rect 146536 78628 147220 78656
rect 146536 78616 146542 78628
rect 147214 78616 147220 78628
rect 147272 78616 147278 78668
rect 147674 78616 147680 78668
rect 147732 78656 147738 78668
rect 147858 78656 147864 78668
rect 147732 78628 147864 78656
rect 147732 78616 147738 78628
rect 147858 78616 147864 78628
rect 147916 78616 147922 78668
rect 151004 78656 151032 78888
rect 155862 78820 155868 78872
rect 155920 78860 155926 78872
rect 159468 78860 159496 78900
rect 155920 78832 159496 78860
rect 155920 78820 155926 78832
rect 160830 78820 160836 78872
rect 160888 78860 160894 78872
rect 161198 78860 161204 78872
rect 160888 78832 161204 78860
rect 160888 78820 160894 78832
rect 161198 78820 161204 78832
rect 161256 78820 161262 78872
rect 165982 78820 165988 78872
rect 166040 78860 166046 78872
rect 167058 78860 167086 78900
rect 172790 78888 172796 78900
rect 172848 78888 172854 78940
rect 172882 78888 172888 78940
rect 172940 78928 172946 78940
rect 173894 78928 173900 78940
rect 172940 78900 173900 78928
rect 172940 78888 172946 78900
rect 173894 78888 173900 78900
rect 173952 78888 173958 78940
rect 174078 78888 174084 78940
rect 174136 78928 174142 78940
rect 393958 78928 393964 78940
rect 174136 78900 393964 78928
rect 174136 78888 174142 78900
rect 393958 78888 393964 78900
rect 394016 78888 394022 78940
rect 430574 78860 430580 78872
rect 166040 78832 167086 78860
rect 168944 78832 430580 78860
rect 166040 78820 166046 78832
rect 159450 78752 159456 78804
rect 159508 78792 159514 78804
rect 168944 78792 168972 78832
rect 430574 78820 430580 78832
rect 430632 78820 430638 78872
rect 159508 78764 168972 78792
rect 159508 78752 159514 78764
rect 169938 78752 169944 78804
rect 169996 78792 170002 78804
rect 173342 78792 173348 78804
rect 169996 78764 173348 78792
rect 169996 78752 170002 78764
rect 173342 78752 173348 78764
rect 173400 78752 173406 78804
rect 151906 78684 151912 78736
rect 151964 78724 151970 78736
rect 153102 78724 153108 78736
rect 151964 78696 153108 78724
rect 151964 78684 151970 78696
rect 153102 78684 153108 78696
rect 153160 78684 153166 78736
rect 154850 78684 154856 78736
rect 154908 78724 154914 78736
rect 162394 78724 162400 78736
rect 154908 78696 162400 78724
rect 154908 78684 154914 78696
rect 162394 78684 162400 78696
rect 162452 78684 162458 78736
rect 174262 78724 174268 78736
rect 167288 78696 174268 78724
rect 151078 78656 151084 78668
rect 151004 78628 151084 78656
rect 151078 78616 151084 78628
rect 151136 78616 151142 78668
rect 158806 78616 158812 78668
rect 158864 78656 158870 78668
rect 158990 78656 158996 78668
rect 158864 78628 158996 78656
rect 158864 78616 158870 78628
rect 158990 78616 158996 78628
rect 159048 78616 159054 78668
rect 159082 78616 159088 78668
rect 159140 78656 159146 78668
rect 161290 78656 161296 78668
rect 159140 78628 161296 78656
rect 159140 78616 159146 78628
rect 161290 78616 161296 78628
rect 161348 78616 161354 78668
rect 166258 78656 166264 78668
rect 162044 78628 166264 78656
rect 136542 78548 136548 78600
rect 136600 78588 136606 78600
rect 144454 78588 144460 78600
rect 136600 78560 144460 78588
rect 136600 78548 136606 78560
rect 144454 78548 144460 78560
rect 144512 78548 144518 78600
rect 145282 78548 145288 78600
rect 145340 78588 145346 78600
rect 162044 78588 162072 78628
rect 166258 78616 166264 78628
rect 166316 78616 166322 78668
rect 145340 78560 162072 78588
rect 145340 78548 145346 78560
rect 164970 78548 164976 78600
rect 165028 78588 165034 78600
rect 165246 78588 165252 78600
rect 165028 78560 165252 78588
rect 165028 78548 165034 78560
rect 165246 78548 165252 78560
rect 165304 78548 165310 78600
rect 166994 78548 167000 78600
rect 167052 78588 167058 78600
rect 167288 78588 167316 78696
rect 174262 78684 174268 78696
rect 174320 78684 174326 78736
rect 168834 78616 168840 78668
rect 168892 78656 168898 78668
rect 170766 78656 170772 78668
rect 168892 78628 170772 78656
rect 168892 78616 168898 78628
rect 170766 78616 170772 78628
rect 170824 78616 170830 78668
rect 171870 78616 171876 78668
rect 171928 78656 171934 78668
rect 178034 78656 178040 78668
rect 171928 78628 178040 78656
rect 171928 78616 171934 78628
rect 178034 78616 178040 78628
rect 178092 78616 178098 78668
rect 167052 78560 167316 78588
rect 167052 78548 167058 78560
rect 171594 78548 171600 78600
rect 171652 78588 171658 78600
rect 396810 78588 396816 78600
rect 171652 78560 396816 78588
rect 171652 78548 171658 78560
rect 396810 78548 396816 78560
rect 396868 78548 396874 78600
rect 139486 78480 139492 78532
rect 139544 78520 139550 78532
rect 171778 78520 171784 78532
rect 139544 78492 171784 78520
rect 139544 78480 139550 78492
rect 171778 78480 171784 78492
rect 171836 78480 171842 78532
rect 172054 78480 172060 78532
rect 172112 78520 172118 78532
rect 178954 78520 178960 78532
rect 172112 78492 178960 78520
rect 172112 78480 172118 78492
rect 178954 78480 178960 78492
rect 179012 78480 179018 78532
rect 133564 78424 133644 78452
rect 133564 78412 133570 78424
rect 140682 78412 140688 78464
rect 140740 78452 140746 78464
rect 195974 78452 195980 78464
rect 140740 78424 195980 78452
rect 140740 78412 140746 78424
rect 195974 78412 195980 78424
rect 196032 78412 196038 78464
rect 133690 78344 133696 78396
rect 133748 78344 133754 78396
rect 140774 78344 140780 78396
rect 140832 78384 140838 78396
rect 141326 78384 141332 78396
rect 140832 78356 141332 78384
rect 140832 78344 140838 78356
rect 141326 78344 141332 78356
rect 141384 78344 141390 78396
rect 145190 78344 145196 78396
rect 145248 78384 145254 78396
rect 147306 78384 147312 78396
rect 145248 78356 147312 78384
rect 145248 78344 145254 78356
rect 147306 78344 147312 78356
rect 147364 78344 147370 78396
rect 150710 78344 150716 78396
rect 150768 78384 150774 78396
rect 150894 78384 150900 78396
rect 150768 78356 150900 78384
rect 150768 78344 150774 78356
rect 150894 78344 150900 78356
rect 150952 78344 150958 78396
rect 159542 78344 159548 78396
rect 159600 78384 159606 78396
rect 160002 78384 160008 78396
rect 159600 78356 160008 78384
rect 159600 78344 159606 78356
rect 160002 78344 160008 78356
rect 160060 78344 160066 78396
rect 160830 78344 160836 78396
rect 160888 78384 160894 78396
rect 161014 78384 161020 78396
rect 160888 78356 161020 78384
rect 160888 78344 160894 78356
rect 161014 78344 161020 78356
rect 161072 78344 161078 78396
rect 161106 78344 161112 78396
rect 161164 78384 161170 78396
rect 255958 78384 255964 78396
rect 161164 78356 255964 78384
rect 161164 78344 161170 78356
rect 255958 78344 255964 78356
rect 256016 78344 256022 78396
rect 132954 78276 132960 78328
rect 133012 78316 133018 78328
rect 133708 78316 133736 78344
rect 133012 78288 133736 78316
rect 133012 78276 133018 78288
rect 145834 78276 145840 78328
rect 145892 78316 145898 78328
rect 150802 78316 150808 78328
rect 145892 78288 150808 78316
rect 145892 78276 145898 78288
rect 150802 78276 150808 78288
rect 150860 78276 150866 78328
rect 153654 78276 153660 78328
rect 153712 78316 153718 78328
rect 157242 78316 157248 78328
rect 153712 78288 157248 78316
rect 153712 78276 153718 78288
rect 157242 78276 157248 78288
rect 157300 78276 157306 78328
rect 158622 78276 158628 78328
rect 158680 78316 158686 78328
rect 158990 78316 158996 78328
rect 158680 78288 158996 78316
rect 158680 78276 158686 78288
rect 158990 78276 158996 78288
rect 159048 78276 159054 78328
rect 162578 78276 162584 78328
rect 162636 78316 162642 78328
rect 315298 78316 315304 78328
rect 162636 78288 315304 78316
rect 162636 78276 162642 78288
rect 315298 78276 315304 78288
rect 315356 78276 315362 78328
rect 106918 78208 106924 78260
rect 106976 78248 106982 78260
rect 127434 78248 127440 78260
rect 106976 78220 127440 78248
rect 106976 78208 106982 78220
rect 127434 78208 127440 78220
rect 127492 78208 127498 78260
rect 133690 78208 133696 78260
rect 133748 78248 133754 78260
rect 137002 78248 137008 78260
rect 133748 78220 137008 78248
rect 133748 78208 133754 78220
rect 137002 78208 137008 78220
rect 137060 78208 137066 78260
rect 140866 78208 140872 78260
rect 140924 78248 140930 78260
rect 141326 78248 141332 78260
rect 140924 78220 141332 78248
rect 140924 78208 140930 78220
rect 141326 78208 141332 78220
rect 141384 78208 141390 78260
rect 156414 78208 156420 78260
rect 156472 78248 156478 78260
rect 161014 78248 161020 78260
rect 156472 78220 161020 78248
rect 156472 78208 156478 78220
rect 161014 78208 161020 78220
rect 161072 78208 161078 78260
rect 164786 78208 164792 78260
rect 164844 78248 164850 78260
rect 341518 78248 341524 78260
rect 164844 78220 341524 78248
rect 164844 78208 164850 78220
rect 341518 78208 341524 78220
rect 341576 78208 341582 78260
rect 110414 78140 110420 78192
rect 110472 78180 110478 78192
rect 123110 78180 123116 78192
rect 110472 78152 123116 78180
rect 110472 78140 110478 78152
rect 123110 78140 123116 78152
rect 123168 78140 123174 78192
rect 141050 78140 141056 78192
rect 141108 78180 141114 78192
rect 141108 78152 148916 78180
rect 141108 78140 141114 78152
rect 89714 78072 89720 78124
rect 89772 78112 89778 78124
rect 132494 78112 132500 78124
rect 89772 78084 132500 78112
rect 89772 78072 89778 78084
rect 132494 78072 132500 78084
rect 132552 78072 132558 78124
rect 140406 78072 140412 78124
rect 140464 78112 140470 78124
rect 148778 78112 148784 78124
rect 140464 78084 148784 78112
rect 140464 78072 140470 78084
rect 148778 78072 148784 78084
rect 148836 78072 148842 78124
rect 71774 78004 71780 78056
rect 71832 78044 71838 78056
rect 126146 78044 126152 78056
rect 71832 78016 126152 78044
rect 71832 78004 71838 78016
rect 126146 78004 126152 78016
rect 126204 78004 126210 78056
rect 132770 78004 132776 78056
rect 132828 78044 132834 78056
rect 133322 78044 133328 78056
rect 132828 78016 133328 78044
rect 132828 78004 132834 78016
rect 133322 78004 133328 78016
rect 133380 78004 133386 78056
rect 148888 78044 148916 78152
rect 149054 78140 149060 78192
rect 149112 78180 149118 78192
rect 151538 78180 151544 78192
rect 149112 78152 151544 78180
rect 149112 78140 149118 78152
rect 151538 78140 151544 78152
rect 151596 78140 151602 78192
rect 152458 78140 152464 78192
rect 152516 78140 152522 78192
rect 154850 78140 154856 78192
rect 154908 78180 154914 78192
rect 155310 78180 155316 78192
rect 154908 78152 155316 78180
rect 154908 78140 154914 78152
rect 155310 78140 155316 78152
rect 155368 78140 155374 78192
rect 157334 78140 157340 78192
rect 157392 78180 157398 78192
rect 157702 78180 157708 78192
rect 157392 78152 157708 78180
rect 157392 78140 157398 78152
rect 157702 78140 157708 78152
rect 157760 78140 157766 78192
rect 163682 78140 163688 78192
rect 163740 78180 163746 78192
rect 480254 78180 480260 78192
rect 163740 78152 480260 78180
rect 163740 78140 163746 78152
rect 480254 78140 480260 78152
rect 480312 78140 480318 78192
rect 152476 78112 152504 78140
rect 162210 78112 162216 78124
rect 152476 78084 162216 78112
rect 162210 78072 162216 78084
rect 162268 78072 162274 78124
rect 163130 78072 163136 78124
rect 163188 78112 163194 78124
rect 163498 78112 163504 78124
rect 163188 78084 163504 78112
rect 163188 78072 163194 78084
rect 163498 78072 163504 78084
rect 163556 78072 163562 78124
rect 167178 78072 167184 78124
rect 167236 78112 167242 78124
rect 532694 78112 532700 78124
rect 167236 78084 532700 78112
rect 167236 78072 167242 78084
rect 532694 78072 532700 78084
rect 532752 78072 532758 78124
rect 152458 78044 152464 78056
rect 148888 78016 152464 78044
rect 152458 78004 152464 78016
rect 152516 78004 152522 78056
rect 153470 78004 153476 78056
rect 153528 78044 153534 78056
rect 153654 78044 153660 78056
rect 153528 78016 153660 78044
rect 153528 78004 153534 78016
rect 153654 78004 153660 78016
rect 153712 78004 153718 78056
rect 154482 78004 154488 78056
rect 154540 78044 154546 78056
rect 155126 78044 155132 78056
rect 154540 78016 155132 78044
rect 154540 78004 154546 78016
rect 155126 78004 155132 78016
rect 155184 78004 155190 78056
rect 156506 78004 156512 78056
rect 156564 78044 156570 78056
rect 156564 78016 164234 78044
rect 156564 78004 156570 78016
rect 53834 77936 53840 77988
rect 53892 77976 53898 77988
rect 129734 77976 129740 77988
rect 53892 77948 129740 77976
rect 53892 77936 53898 77948
rect 129734 77936 129740 77948
rect 129792 77936 129798 77988
rect 134702 77976 134708 77988
rect 131040 77948 134708 77976
rect 123662 77868 123668 77920
rect 123720 77908 123726 77920
rect 131040 77908 131068 77948
rect 134702 77936 134708 77948
rect 134760 77936 134766 77988
rect 139762 77936 139768 77988
rect 139820 77976 139826 77988
rect 139820 77948 147674 77976
rect 139820 77936 139826 77948
rect 123720 77880 131068 77908
rect 123720 77868 123726 77880
rect 132862 77868 132868 77920
rect 132920 77908 132926 77920
rect 133322 77908 133328 77920
rect 132920 77880 133328 77908
rect 132920 77868 132926 77880
rect 133322 77868 133328 77880
rect 133380 77868 133386 77920
rect 137646 77868 137652 77920
rect 137704 77908 137710 77920
rect 140406 77908 140412 77920
rect 137704 77880 140412 77908
rect 137704 77868 137710 77880
rect 140406 77868 140412 77880
rect 140464 77868 140470 77920
rect 147646 77908 147674 77948
rect 154574 77936 154580 77988
rect 154632 77976 154638 77988
rect 155034 77976 155040 77988
rect 154632 77948 155040 77976
rect 154632 77936 154638 77948
rect 155034 77936 155040 77948
rect 155092 77936 155098 77988
rect 156046 77936 156052 77988
rect 156104 77976 156110 77988
rect 156598 77976 156604 77988
rect 156104 77948 156604 77976
rect 156104 77936 156110 77948
rect 156598 77936 156604 77948
rect 156656 77936 156662 77988
rect 157702 77936 157708 77988
rect 157760 77976 157766 77988
rect 157978 77976 157984 77988
rect 157760 77948 157984 77976
rect 157760 77936 157766 77948
rect 157978 77936 157984 77948
rect 158036 77936 158042 77988
rect 164206 77976 164234 78016
rect 165982 78004 165988 78056
rect 166040 78044 166046 78056
rect 166040 78016 167086 78044
rect 166040 78004 166046 78016
rect 167058 77976 167086 78016
rect 170674 78004 170680 78056
rect 170732 78044 170738 78056
rect 538858 78044 538864 78056
rect 170732 78016 538864 78044
rect 170732 78004 170738 78016
rect 538858 78004 538864 78016
rect 538916 78004 538922 78056
rect 174446 77976 174452 77988
rect 164206 77948 166994 77976
rect 167058 77948 174452 77976
rect 147646 77880 160692 77908
rect 131114 77800 131120 77852
rect 131172 77840 131178 77852
rect 133874 77840 133880 77852
rect 131172 77812 133880 77840
rect 131172 77800 131178 77812
rect 133874 77800 133880 77812
rect 133932 77800 133938 77852
rect 140958 77800 140964 77852
rect 141016 77840 141022 77852
rect 141694 77840 141700 77852
rect 141016 77812 141700 77840
rect 141016 77800 141022 77812
rect 141694 77800 141700 77812
rect 141752 77800 141758 77852
rect 143534 77800 143540 77852
rect 143592 77840 143598 77852
rect 144362 77840 144368 77852
rect 143592 77812 144368 77840
rect 143592 77800 143598 77812
rect 144362 77800 144368 77812
rect 144420 77800 144426 77852
rect 149146 77800 149152 77852
rect 149204 77840 149210 77852
rect 149882 77840 149888 77852
rect 149204 77812 149888 77840
rect 149204 77800 149210 77812
rect 149882 77800 149888 77812
rect 149940 77800 149946 77852
rect 153286 77800 153292 77852
rect 153344 77840 153350 77852
rect 153746 77840 153752 77852
rect 153344 77812 153752 77840
rect 153344 77800 153350 77812
rect 153746 77800 153752 77812
rect 153804 77800 153810 77852
rect 155034 77732 155040 77784
rect 155092 77772 155098 77784
rect 155402 77772 155408 77784
rect 155092 77744 155408 77772
rect 155092 77732 155098 77744
rect 155402 77732 155408 77744
rect 155460 77732 155466 77784
rect 157610 77732 157616 77784
rect 157668 77772 157674 77784
rect 160664 77772 160692 77880
rect 166966 77840 166994 77948
rect 174446 77936 174452 77948
rect 174504 77936 174510 77988
rect 580994 77976 581000 77988
rect 176626 77948 581000 77976
rect 171410 77868 171416 77920
rect 171468 77908 171474 77920
rect 176626 77908 176654 77948
rect 580994 77936 581000 77948
rect 581052 77936 581058 77988
rect 171468 77880 176654 77908
rect 171468 77868 171474 77880
rect 171962 77840 171968 77852
rect 166966 77812 171968 77840
rect 171962 77800 171968 77812
rect 172020 77800 172026 77852
rect 171870 77772 171876 77784
rect 157668 77744 160600 77772
rect 160664 77744 171876 77772
rect 157668 77732 157674 77744
rect 125134 77664 125140 77716
rect 125192 77704 125198 77716
rect 134058 77704 134064 77716
rect 125192 77676 134064 77704
rect 125192 77664 125198 77676
rect 134058 77664 134064 77676
rect 134116 77664 134122 77716
rect 134518 77664 134524 77716
rect 134576 77704 134582 77716
rect 135346 77704 135352 77716
rect 134576 77676 135352 77704
rect 134576 77664 134582 77676
rect 135346 77664 135352 77676
rect 135404 77664 135410 77716
rect 149422 77664 149428 77716
rect 149480 77704 149486 77716
rect 149882 77704 149888 77716
rect 149480 77676 149888 77704
rect 149480 77664 149486 77676
rect 149882 77664 149888 77676
rect 149940 77664 149946 77716
rect 160572 77704 160600 77744
rect 171870 77732 171876 77744
rect 171928 77732 171934 77784
rect 171410 77704 171416 77716
rect 160572 77676 171416 77704
rect 171410 77664 171416 77676
rect 171468 77664 171474 77716
rect 136634 77596 136640 77648
rect 136692 77636 136698 77648
rect 139118 77636 139124 77648
rect 136692 77608 139124 77636
rect 136692 77596 136698 77608
rect 139118 77596 139124 77608
rect 139176 77596 139182 77648
rect 144914 77596 144920 77648
rect 144972 77636 144978 77648
rect 157058 77636 157064 77648
rect 144972 77608 157064 77636
rect 144972 77596 144978 77608
rect 157058 77596 157064 77608
rect 157116 77596 157122 77648
rect 160094 77596 160100 77648
rect 160152 77636 160158 77648
rect 171686 77636 171692 77648
rect 160152 77608 171692 77636
rect 160152 77596 160158 77608
rect 171686 77596 171692 77608
rect 171744 77596 171750 77648
rect 123110 77528 123116 77580
rect 123168 77568 123174 77580
rect 131022 77568 131028 77580
rect 123168 77540 131028 77568
rect 123168 77528 123174 77540
rect 131022 77528 131028 77540
rect 131080 77528 131086 77580
rect 141786 77528 141792 77580
rect 141844 77568 141850 77580
rect 172238 77568 172244 77580
rect 141844 77540 172244 77568
rect 141844 77528 141850 77540
rect 172238 77528 172244 77540
rect 172296 77528 172302 77580
rect 172790 77528 172796 77580
rect 172848 77568 172854 77580
rect 396718 77568 396724 77580
rect 172848 77540 396724 77568
rect 172848 77528 172854 77540
rect 396718 77528 396724 77540
rect 396776 77528 396782 77580
rect 147950 77460 147956 77512
rect 148008 77500 148014 77512
rect 166994 77500 167000 77512
rect 148008 77472 167000 77500
rect 148008 77460 148014 77472
rect 166994 77460 167000 77472
rect 167052 77460 167058 77512
rect 169018 77500 169024 77512
rect 167104 77472 169024 77500
rect 122926 77392 122932 77444
rect 122984 77432 122990 77444
rect 130102 77432 130108 77444
rect 122984 77404 130108 77432
rect 122984 77392 122990 77404
rect 130102 77392 130108 77404
rect 130160 77392 130166 77444
rect 133874 77392 133880 77444
rect 133932 77432 133938 77444
rect 135990 77432 135996 77444
rect 133932 77404 135996 77432
rect 133932 77392 133938 77404
rect 135990 77392 135996 77404
rect 136048 77392 136054 77444
rect 150526 77392 150532 77444
rect 150584 77432 150590 77444
rect 158346 77432 158352 77444
rect 150584 77404 158352 77432
rect 150584 77392 150590 77404
rect 158346 77392 158352 77404
rect 158404 77392 158410 77444
rect 164418 77392 164424 77444
rect 164476 77432 164482 77444
rect 167104 77432 167132 77472
rect 169018 77460 169024 77472
rect 169076 77460 169082 77512
rect 171778 77460 171784 77512
rect 171836 77500 171842 77512
rect 178034 77500 178040 77512
rect 171836 77472 178040 77500
rect 171836 77460 171842 77472
rect 178034 77460 178040 77472
rect 178092 77460 178098 77512
rect 164476 77404 167132 77432
rect 164476 77392 164482 77404
rect 145006 77324 145012 77376
rect 145064 77364 145070 77376
rect 145742 77364 145748 77376
rect 145064 77336 145748 77364
rect 145064 77324 145070 77336
rect 145742 77324 145748 77336
rect 145800 77324 145806 77376
rect 155862 77324 155868 77376
rect 155920 77364 155926 77376
rect 156598 77364 156604 77376
rect 155920 77336 156604 77364
rect 155920 77324 155926 77336
rect 156598 77324 156604 77336
rect 156656 77324 156662 77376
rect 161106 77324 161112 77376
rect 161164 77364 161170 77376
rect 172146 77364 172152 77376
rect 161164 77336 172152 77364
rect 161164 77324 161170 77336
rect 172146 77324 172152 77336
rect 172204 77324 172210 77376
rect 128998 77256 129004 77308
rect 129056 77296 129062 77308
rect 131666 77296 131672 77308
rect 129056 77268 131672 77296
rect 129056 77256 129062 77268
rect 131666 77256 131672 77268
rect 131724 77256 131730 77308
rect 135714 77256 135720 77308
rect 135772 77296 135778 77308
rect 135990 77296 135996 77308
rect 135772 77268 135996 77296
rect 135772 77256 135778 77268
rect 135990 77256 135996 77268
rect 136048 77256 136054 77308
rect 139946 77256 139952 77308
rect 140004 77296 140010 77308
rect 140222 77296 140228 77308
rect 140004 77268 140228 77296
rect 140004 77256 140010 77268
rect 140222 77256 140228 77268
rect 140280 77256 140286 77308
rect 151906 77256 151912 77308
rect 151964 77296 151970 77308
rect 152182 77296 152188 77308
rect 151964 77268 152188 77296
rect 151964 77256 151970 77268
rect 152182 77256 152188 77268
rect 152240 77256 152246 77308
rect 154206 77256 154212 77308
rect 154264 77296 154270 77308
rect 157978 77296 157984 77308
rect 154264 77268 157984 77296
rect 154264 77256 154270 77268
rect 157978 77256 157984 77268
rect 158036 77256 158042 77308
rect 160646 77256 160652 77308
rect 160704 77296 160710 77308
rect 166902 77296 166908 77308
rect 160704 77268 166908 77296
rect 160704 77256 160710 77268
rect 166902 77256 166908 77268
rect 166960 77256 166966 77308
rect 169018 77256 169024 77308
rect 169076 77296 169082 77308
rect 171686 77296 171692 77308
rect 169076 77268 171692 77296
rect 169076 77256 169082 77268
rect 171686 77256 171692 77268
rect 171744 77256 171750 77308
rect 121822 77188 121828 77240
rect 121880 77228 121886 77240
rect 123938 77228 123944 77240
rect 121880 77200 123944 77228
rect 121880 77188 121886 77200
rect 123938 77188 123944 77200
rect 123996 77188 124002 77240
rect 131390 77188 131396 77240
rect 131448 77228 131454 77240
rect 131942 77228 131948 77240
rect 131448 77200 131948 77228
rect 131448 77188 131454 77200
rect 131942 77188 131948 77200
rect 132000 77188 132006 77240
rect 139486 77188 139492 77240
rect 139544 77228 139550 77240
rect 140130 77228 140136 77240
rect 139544 77200 140136 77228
rect 139544 77188 139550 77200
rect 140130 77188 140136 77200
rect 140188 77188 140194 77240
rect 153470 77188 153476 77240
rect 153528 77228 153534 77240
rect 154022 77228 154028 77240
rect 153528 77200 154028 77228
rect 153528 77188 153534 77200
rect 154022 77188 154028 77200
rect 154080 77188 154086 77240
rect 162210 77188 162216 77240
rect 162268 77228 162274 77240
rect 197354 77228 197360 77240
rect 162268 77200 197360 77228
rect 162268 77188 162274 77200
rect 197354 77188 197360 77200
rect 197412 77188 197418 77240
rect 139302 77120 139308 77172
rect 139360 77160 139366 77172
rect 140590 77160 140596 77172
rect 139360 77132 140596 77160
rect 139360 77120 139366 77132
rect 140590 77120 140596 77132
rect 140648 77120 140654 77172
rect 142246 77120 142252 77172
rect 142304 77160 142310 77172
rect 213914 77160 213920 77172
rect 142304 77132 213920 77160
rect 142304 77120 142310 77132
rect 213914 77120 213920 77132
rect 213972 77120 213978 77172
rect 126974 77052 126980 77104
rect 127032 77092 127038 77104
rect 129182 77092 129188 77104
rect 127032 77064 129188 77092
rect 127032 77052 127038 77064
rect 129182 77052 129188 77064
rect 129240 77052 129246 77104
rect 131298 77052 131304 77104
rect 131356 77092 131362 77104
rect 132126 77092 132132 77104
rect 131356 77064 132132 77092
rect 131356 77052 131362 77064
rect 132126 77052 132132 77064
rect 132184 77052 132190 77104
rect 143166 77052 143172 77104
rect 143224 77092 143230 77104
rect 226334 77092 226340 77104
rect 143224 77064 226340 77092
rect 143224 77052 143230 77064
rect 226334 77052 226340 77064
rect 226392 77052 226398 77104
rect 143442 76984 143448 77036
rect 143500 77024 143506 77036
rect 231854 77024 231860 77036
rect 143500 76996 231860 77024
rect 143500 76984 143506 76996
rect 231854 76984 231860 76996
rect 231912 76984 231918 77036
rect 129182 76916 129188 76968
rect 129240 76956 129246 76968
rect 129918 76956 129924 76968
rect 129240 76928 129924 76956
rect 129240 76916 129246 76928
rect 129918 76916 129924 76928
rect 129976 76916 129982 76968
rect 144178 76916 144184 76968
rect 144236 76956 144242 76968
rect 240134 76956 240140 76968
rect 144236 76928 240140 76956
rect 144236 76916 144242 76928
rect 240134 76916 240140 76928
rect 240192 76916 240198 76968
rect 122098 76848 122104 76900
rect 122156 76888 122162 76900
rect 134794 76888 134800 76900
rect 122156 76860 134800 76888
rect 122156 76848 122162 76860
rect 134794 76848 134800 76860
rect 134852 76848 134858 76900
rect 138290 76848 138296 76900
rect 138348 76888 138354 76900
rect 138566 76888 138572 76900
rect 138348 76860 138572 76888
rect 138348 76848 138354 76860
rect 138566 76848 138572 76860
rect 138624 76848 138630 76900
rect 150802 76848 150808 76900
rect 150860 76888 150866 76900
rect 260834 76888 260840 76900
rect 150860 76860 260840 76888
rect 150860 76848 150866 76860
rect 260834 76848 260840 76860
rect 260892 76848 260898 76900
rect 129918 76780 129924 76832
rect 129976 76820 129982 76832
rect 130194 76820 130200 76832
rect 129976 76792 130200 76820
rect 129976 76780 129982 76792
rect 130194 76780 130200 76792
rect 130252 76780 130258 76832
rect 146294 76780 146300 76832
rect 146352 76820 146358 76832
rect 267734 76820 267740 76832
rect 146352 76792 267740 76820
rect 146352 76780 146358 76792
rect 267734 76780 267740 76792
rect 267792 76780 267798 76832
rect 102134 76712 102140 76764
rect 102192 76752 102198 76764
rect 132402 76752 132408 76764
rect 102192 76724 132408 76752
rect 102192 76712 102198 76724
rect 132402 76712 132408 76724
rect 132460 76712 132466 76764
rect 142246 76712 142252 76764
rect 142304 76752 142310 76764
rect 142706 76752 142712 76764
rect 142304 76724 142712 76752
rect 142304 76712 142310 76724
rect 142706 76712 142712 76724
rect 142764 76712 142770 76764
rect 147766 76712 147772 76764
rect 147824 76752 147830 76764
rect 284294 76752 284300 76764
rect 147824 76724 284300 76752
rect 147824 76712 147830 76724
rect 284294 76712 284300 76724
rect 284352 76712 284358 76764
rect 86954 76644 86960 76696
rect 87012 76684 87018 76696
rect 132310 76684 132316 76696
rect 87012 76656 132316 76684
rect 87012 76644 87018 76656
rect 132310 76644 132316 76656
rect 132368 76644 132374 76696
rect 145098 76644 145104 76696
rect 145156 76684 145162 76696
rect 145374 76684 145380 76696
rect 145156 76656 145380 76684
rect 145156 76644 145162 76656
rect 145374 76644 145380 76656
rect 145432 76644 145438 76696
rect 152550 76644 152556 76696
rect 152608 76684 152614 76696
rect 153102 76684 153108 76696
rect 152608 76656 153108 76684
rect 152608 76644 152614 76656
rect 153102 76644 153108 76656
rect 153160 76644 153166 76696
rect 156138 76644 156144 76696
rect 156196 76684 156202 76696
rect 156874 76684 156880 76696
rect 156196 76656 156880 76684
rect 156196 76644 156202 76656
rect 156874 76644 156880 76656
rect 156932 76644 156938 76696
rect 157518 76644 157524 76696
rect 157576 76684 157582 76696
rect 296714 76684 296720 76696
rect 157576 76656 296720 76684
rect 157576 76644 157582 76656
rect 296714 76644 296720 76656
rect 296772 76644 296778 76696
rect 44174 76576 44180 76628
rect 44232 76616 44238 76628
rect 120902 76616 120908 76628
rect 44232 76588 120908 76616
rect 44232 76576 44238 76588
rect 120902 76576 120908 76588
rect 120960 76576 120966 76628
rect 130194 76576 130200 76628
rect 130252 76616 130258 76628
rect 130562 76616 130568 76628
rect 130252 76588 130568 76616
rect 130252 76576 130258 76588
rect 130562 76576 130568 76588
rect 130620 76576 130626 76628
rect 142338 76576 142344 76628
rect 142396 76616 142402 76628
rect 142798 76616 142804 76628
rect 142396 76588 142804 76616
rect 142396 76576 142402 76588
rect 142798 76576 142804 76588
rect 142856 76576 142862 76628
rect 146018 76576 146024 76628
rect 146076 76616 146082 76628
rect 146754 76616 146760 76628
rect 146076 76588 146760 76616
rect 146076 76576 146082 76588
rect 146754 76576 146760 76588
rect 146812 76576 146818 76628
rect 147950 76576 147956 76628
rect 148008 76616 148014 76628
rect 148410 76616 148416 76628
rect 148008 76588 148416 76616
rect 148008 76576 148014 76588
rect 148410 76576 148416 76588
rect 148468 76576 148474 76628
rect 151538 76576 151544 76628
rect 151596 76616 151602 76628
rect 151596 76588 154574 76616
rect 151596 76576 151602 76588
rect 30374 76508 30380 76560
rect 30432 76548 30438 76560
rect 30432 76520 120074 76548
rect 30432 76508 30438 76520
rect 120046 76480 120074 76520
rect 137554 76508 137560 76560
rect 137612 76548 137618 76560
rect 144454 76548 144460 76560
rect 137612 76520 144460 76548
rect 137612 76508 137618 76520
rect 144454 76508 144460 76520
rect 144512 76508 144518 76560
rect 154546 76548 154574 76588
rect 156322 76576 156328 76628
rect 156380 76616 156386 76628
rect 156506 76616 156512 76628
rect 156380 76588 156512 76616
rect 156380 76576 156386 76588
rect 156506 76576 156512 76588
rect 156564 76576 156570 76628
rect 157426 76576 157432 76628
rect 157484 76616 157490 76628
rect 158162 76616 158168 76628
rect 157484 76588 158168 76616
rect 157484 76576 157490 76588
rect 158162 76576 158168 76588
rect 158220 76576 158226 76628
rect 302234 76616 302240 76628
rect 162412 76588 302240 76616
rect 162412 76548 162440 76588
rect 302234 76576 302240 76588
rect 302292 76576 302298 76628
rect 154546 76520 162440 76548
rect 171226 76508 171232 76560
rect 171284 76548 171290 76560
rect 373994 76548 374000 76560
rect 171284 76520 374000 76548
rect 171284 76508 171290 76520
rect 373994 76508 374000 76520
rect 374052 76508 374058 76560
rect 126330 76480 126336 76492
rect 120046 76452 126336 76480
rect 126330 76440 126336 76452
rect 126388 76440 126394 76492
rect 130102 76440 130108 76492
rect 130160 76480 130166 76492
rect 130654 76480 130660 76492
rect 130160 76452 130660 76480
rect 130160 76440 130166 76452
rect 130654 76440 130660 76452
rect 130712 76440 130718 76492
rect 141142 76440 141148 76492
rect 141200 76480 141206 76492
rect 141510 76480 141516 76492
rect 141200 76452 141516 76480
rect 141200 76440 141206 76452
rect 141510 76440 141516 76452
rect 141568 76440 141574 76492
rect 142154 76440 142160 76492
rect 142212 76480 142218 76492
rect 142614 76480 142620 76492
rect 142212 76452 142620 76480
rect 142212 76440 142218 76452
rect 142614 76440 142620 76452
rect 142672 76440 142678 76492
rect 147766 76440 147772 76492
rect 147824 76480 147830 76492
rect 148594 76480 148600 76492
rect 147824 76452 148600 76480
rect 147824 76440 147830 76452
rect 148594 76440 148600 76452
rect 148652 76440 148658 76492
rect 152458 76440 152464 76492
rect 152516 76480 152522 76492
rect 162210 76480 162216 76492
rect 152516 76452 162216 76480
rect 152516 76440 152522 76452
rect 162210 76440 162216 76452
rect 162268 76440 162274 76492
rect 153194 76372 153200 76424
rect 153252 76412 153258 76424
rect 157518 76412 157524 76424
rect 153252 76384 157524 76412
rect 153252 76372 153258 76384
rect 157518 76372 157524 76384
rect 157576 76372 157582 76424
rect 145374 76304 145380 76356
rect 145432 76344 145438 76356
rect 145650 76344 145656 76356
rect 145432 76316 145656 76344
rect 145432 76304 145438 76316
rect 145650 76304 145656 76316
rect 145708 76304 145714 76356
rect 162486 76304 162492 76356
rect 162544 76344 162550 76356
rect 173250 76344 173256 76356
rect 162544 76316 173256 76344
rect 162544 76304 162550 76316
rect 173250 76304 173256 76316
rect 173308 76304 173314 76356
rect 153194 76236 153200 76288
rect 153252 76276 153258 76288
rect 153930 76276 153936 76288
rect 153252 76248 153936 76276
rect 153252 76236 153258 76248
rect 153930 76236 153936 76248
rect 153988 76236 153994 76288
rect 157518 76236 157524 76288
rect 157576 76276 157582 76288
rect 158254 76276 158260 76288
rect 157576 76248 158260 76276
rect 157576 76236 157582 76248
rect 158254 76236 158260 76248
rect 158312 76236 158318 76288
rect 161934 76236 161940 76288
rect 161992 76276 161998 76288
rect 162118 76276 162124 76288
rect 161992 76248 162124 76276
rect 161992 76236 161998 76248
rect 162118 76236 162124 76248
rect 162176 76236 162182 76288
rect 159082 76168 159088 76220
rect 159140 76208 159146 76220
rect 159266 76208 159272 76220
rect 159140 76180 159272 76208
rect 159140 76168 159146 76180
rect 159266 76168 159272 76180
rect 159324 76168 159330 76220
rect 120902 76100 120908 76152
rect 120960 76140 120966 76152
rect 128262 76140 128268 76152
rect 120960 76112 128268 76140
rect 120960 76100 120966 76112
rect 128262 76100 128268 76112
rect 128320 76100 128326 76152
rect 161750 76100 161756 76152
rect 161808 76140 161814 76152
rect 162118 76140 162124 76152
rect 161808 76112 162124 76140
rect 161808 76100 161814 76112
rect 162118 76100 162124 76112
rect 162176 76100 162182 76152
rect 122282 76032 122288 76084
rect 122340 76072 122346 76084
rect 127342 76072 127348 76084
rect 122340 76044 127348 76072
rect 122340 76032 122346 76044
rect 127342 76032 127348 76044
rect 127400 76032 127406 76084
rect 145098 76032 145104 76084
rect 145156 76072 145162 76084
rect 145926 76072 145932 76084
rect 145156 76044 145932 76072
rect 145156 76032 145162 76044
rect 145926 76032 145932 76044
rect 145984 76032 145990 76084
rect 161566 76032 161572 76084
rect 161624 76072 161630 76084
rect 161624 76044 161796 76072
rect 161624 76032 161630 76044
rect 161768 76016 161796 76044
rect 167454 76032 167460 76084
rect 167512 76072 167518 76084
rect 167914 76072 167920 76084
rect 167512 76044 167920 76072
rect 167512 76032 167518 76044
rect 167914 76032 167920 76044
rect 167972 76032 167978 76084
rect 155770 75964 155776 76016
rect 155828 76004 155834 76016
rect 156966 76004 156972 76016
rect 155828 75976 156972 76004
rect 155828 75964 155834 75976
rect 156966 75964 156972 75976
rect 157024 75964 157030 76016
rect 161750 75964 161756 76016
rect 161808 75964 161814 76016
rect 163130 75964 163136 76016
rect 163188 76004 163194 76016
rect 163866 76004 163872 76016
rect 163188 75976 163872 76004
rect 163188 75964 163194 75976
rect 163866 75964 163872 75976
rect 163924 75964 163930 76016
rect 125870 75896 125876 75948
rect 125928 75936 125934 75948
rect 126054 75936 126060 75948
rect 125928 75908 126060 75936
rect 125928 75896 125934 75908
rect 126054 75896 126060 75908
rect 126112 75896 126118 75948
rect 127250 75896 127256 75948
rect 127308 75936 127314 75948
rect 127710 75936 127716 75948
rect 127308 75908 127716 75936
rect 127308 75896 127314 75908
rect 127710 75896 127716 75908
rect 127768 75896 127774 75948
rect 127894 75896 127900 75948
rect 127952 75936 127958 75948
rect 128262 75936 128268 75948
rect 127952 75908 128268 75936
rect 127952 75896 127958 75908
rect 128262 75896 128268 75908
rect 128320 75896 128326 75948
rect 128906 75896 128912 75948
rect 128964 75936 128970 75948
rect 129274 75936 129280 75948
rect 128964 75908 129280 75936
rect 128964 75896 128970 75908
rect 129274 75896 129280 75908
rect 129332 75896 129338 75948
rect 160094 75896 160100 75948
rect 160152 75936 160158 75948
rect 160370 75936 160376 75948
rect 160152 75908 160376 75936
rect 160152 75896 160158 75908
rect 160370 75896 160376 75908
rect 160428 75896 160434 75948
rect 160462 75896 160468 75948
rect 160520 75936 160526 75948
rect 160646 75936 160652 75948
rect 160520 75908 160652 75936
rect 160520 75896 160526 75908
rect 160646 75896 160652 75908
rect 160704 75896 160710 75948
rect 165798 75896 165804 75948
rect 165856 75936 165862 75948
rect 166626 75936 166632 75948
rect 165856 75908 166632 75936
rect 165856 75896 165862 75908
rect 166626 75896 166632 75908
rect 166684 75896 166690 75948
rect 44910 75828 44916 75880
rect 44968 75868 44974 75880
rect 173066 75868 173072 75880
rect 44968 75840 173072 75868
rect 44968 75828 44974 75840
rect 173066 75828 173072 75840
rect 173124 75828 173130 75880
rect 125042 75760 125048 75812
rect 125100 75800 125106 75812
rect 125502 75800 125508 75812
rect 125100 75772 125508 75800
rect 125100 75760 125106 75772
rect 125502 75760 125508 75772
rect 125560 75760 125566 75812
rect 125594 75760 125600 75812
rect 125652 75800 125658 75812
rect 172606 75800 172612 75812
rect 125652 75772 172612 75800
rect 125652 75760 125658 75772
rect 172606 75760 172612 75772
rect 172664 75760 172670 75812
rect 123938 75692 123944 75744
rect 123996 75732 124002 75744
rect 171502 75732 171508 75744
rect 123996 75704 171508 75732
rect 123996 75692 124002 75704
rect 171502 75692 171508 75704
rect 171560 75692 171566 75744
rect 125870 75624 125876 75676
rect 125928 75664 125934 75676
rect 126882 75664 126888 75676
rect 125928 75636 126888 75664
rect 125928 75624 125934 75636
rect 126882 75624 126888 75636
rect 126940 75624 126946 75676
rect 127342 75624 127348 75676
rect 127400 75664 127406 75676
rect 127802 75664 127808 75676
rect 127400 75636 127808 75664
rect 127400 75624 127406 75636
rect 127802 75624 127808 75636
rect 127860 75624 127866 75676
rect 133782 75664 133788 75676
rect 128326 75636 133788 75664
rect 120718 75488 120724 75540
rect 120776 75528 120782 75540
rect 128326 75528 128354 75636
rect 133782 75624 133788 75636
rect 133840 75624 133846 75676
rect 135438 75624 135444 75676
rect 135496 75664 135502 75676
rect 136266 75664 136272 75676
rect 135496 75636 136272 75664
rect 135496 75624 135502 75636
rect 136266 75624 136272 75636
rect 136324 75624 136330 75676
rect 164694 75624 164700 75676
rect 164752 75664 164758 75676
rect 165246 75664 165252 75676
rect 164752 75636 165252 75664
rect 164752 75624 164758 75636
rect 165246 75624 165252 75636
rect 165304 75624 165310 75676
rect 129734 75556 129740 75608
rect 129792 75596 129798 75608
rect 135530 75596 135536 75608
rect 129792 75568 135536 75596
rect 129792 75556 129798 75568
rect 135530 75556 135536 75568
rect 135588 75556 135594 75608
rect 163038 75556 163044 75608
rect 163096 75596 163102 75608
rect 163406 75596 163412 75608
rect 163096 75568 163412 75596
rect 163096 75556 163102 75568
rect 163406 75556 163412 75568
rect 163464 75556 163470 75608
rect 131114 75528 131120 75540
rect 120776 75500 128354 75528
rect 128648 75500 131120 75528
rect 120776 75488 120782 75500
rect 107654 75420 107660 75472
rect 107712 75460 107718 75472
rect 128648 75460 128676 75500
rect 131114 75488 131120 75500
rect 131172 75488 131178 75540
rect 150986 75488 150992 75540
rect 151044 75528 151050 75540
rect 322934 75528 322940 75540
rect 151044 75500 322940 75528
rect 151044 75488 151050 75500
rect 322934 75488 322940 75500
rect 322992 75488 322998 75540
rect 107712 75432 128676 75460
rect 107712 75420 107718 75432
rect 135530 75420 135536 75472
rect 135588 75460 135594 75472
rect 136174 75460 136180 75472
rect 135588 75432 136180 75460
rect 135588 75420 135594 75432
rect 136174 75420 136180 75432
rect 136232 75420 136238 75472
rect 157242 75420 157248 75472
rect 157300 75460 157306 75472
rect 361574 75460 361580 75472
rect 157300 75432 361580 75460
rect 157300 75420 157306 75432
rect 361574 75420 361580 75432
rect 361632 75420 361638 75472
rect 70394 75352 70400 75404
rect 70452 75392 70458 75404
rect 130930 75392 130936 75404
rect 70452 75364 130936 75392
rect 70452 75352 70458 75364
rect 130930 75352 130936 75364
rect 130988 75352 130994 75404
rect 162946 75352 162952 75404
rect 163004 75392 163010 75404
rect 163958 75392 163964 75404
rect 163004 75364 163964 75392
rect 163004 75352 163010 75364
rect 163958 75352 163964 75364
rect 164016 75352 164022 75404
rect 164142 75352 164148 75404
rect 164200 75392 164206 75404
rect 164200 75364 166856 75392
rect 164200 75352 164206 75364
rect 60734 75284 60740 75336
rect 60792 75324 60798 75336
rect 124950 75324 124956 75336
rect 60792 75296 124956 75324
rect 60792 75284 60798 75296
rect 124950 75284 124956 75296
rect 125008 75284 125014 75336
rect 137094 75284 137100 75336
rect 137152 75324 137158 75336
rect 137278 75324 137284 75336
rect 137152 75296 137284 75324
rect 137152 75284 137158 75296
rect 137278 75284 137284 75296
rect 137336 75284 137342 75336
rect 138014 75284 138020 75336
rect 138072 75324 138078 75336
rect 138474 75324 138480 75336
rect 138072 75296 138480 75324
rect 138072 75284 138078 75296
rect 138474 75284 138480 75296
rect 138532 75284 138538 75336
rect 160278 75284 160284 75336
rect 160336 75324 160342 75336
rect 160830 75324 160836 75336
rect 160336 75296 160836 75324
rect 160336 75284 160342 75296
rect 160830 75284 160836 75296
rect 160888 75284 160894 75336
rect 164326 75284 164332 75336
rect 164384 75324 164390 75336
rect 164694 75324 164700 75336
rect 164384 75296 164700 75324
rect 164384 75284 164390 75296
rect 164694 75284 164700 75296
rect 164752 75284 164758 75336
rect 166074 75284 166080 75336
rect 166132 75324 166138 75336
rect 166718 75324 166724 75336
rect 166132 75296 166724 75324
rect 166132 75284 166138 75296
rect 166718 75284 166724 75296
rect 166776 75284 166782 75336
rect 166828 75324 166856 75364
rect 166902 75352 166908 75404
rect 166960 75392 166966 75404
rect 438854 75392 438860 75404
rect 166960 75364 438860 75392
rect 166960 75352 166966 75364
rect 438854 75352 438860 75364
rect 438912 75352 438918 75404
rect 490006 75324 490012 75336
rect 166828 75296 490012 75324
rect 490006 75284 490012 75296
rect 490064 75284 490070 75336
rect 35894 75216 35900 75268
rect 35952 75256 35958 75268
rect 35952 75228 120074 75256
rect 35952 75216 35958 75228
rect 6914 75148 6920 75200
rect 6972 75188 6978 75200
rect 120046 75188 120074 75228
rect 121086 75216 121092 75268
rect 121144 75256 121150 75268
rect 125594 75256 125600 75268
rect 121144 75228 125600 75256
rect 121144 75216 121150 75228
rect 125594 75216 125600 75228
rect 125652 75216 125658 75268
rect 135806 75216 135812 75268
rect 135864 75256 135870 75268
rect 136450 75256 136456 75268
rect 135864 75228 136456 75256
rect 135864 75216 135870 75228
rect 136450 75216 136456 75228
rect 136508 75216 136514 75268
rect 136818 75216 136824 75268
rect 136876 75256 136882 75268
rect 137002 75256 137008 75268
rect 136876 75228 137008 75256
rect 136876 75216 136882 75228
rect 137002 75216 137008 75228
rect 137060 75216 137066 75268
rect 139394 75216 139400 75268
rect 139452 75256 139458 75268
rect 139762 75256 139768 75268
rect 139452 75228 139768 75256
rect 139452 75216 139458 75228
rect 139762 75216 139768 75228
rect 139820 75216 139826 75268
rect 143626 75216 143632 75268
rect 143684 75256 143690 75268
rect 144178 75256 144184 75268
rect 143684 75228 144184 75256
rect 143684 75216 143690 75228
rect 144178 75216 144184 75228
rect 144236 75216 144242 75268
rect 149238 75216 149244 75268
rect 149296 75256 149302 75268
rect 149422 75256 149428 75268
rect 149296 75228 149428 75256
rect 149296 75216 149302 75228
rect 149422 75216 149428 75228
rect 149480 75216 149486 75268
rect 149514 75216 149520 75268
rect 149572 75256 149578 75268
rect 149790 75256 149796 75268
rect 149572 75228 149796 75256
rect 149572 75216 149578 75228
rect 149790 75216 149796 75228
rect 149848 75216 149854 75268
rect 150802 75216 150808 75268
rect 150860 75256 150866 75268
rect 151262 75256 151268 75268
rect 150860 75228 151268 75256
rect 150860 75216 150866 75228
rect 151262 75216 151268 75228
rect 151320 75216 151326 75268
rect 159174 75216 159180 75268
rect 159232 75256 159238 75268
rect 159818 75256 159824 75268
rect 159232 75228 159824 75256
rect 159232 75216 159238 75228
rect 159818 75216 159824 75228
rect 159876 75216 159882 75268
rect 160370 75216 160376 75268
rect 160428 75256 160434 75268
rect 160922 75256 160928 75268
rect 160428 75228 160928 75256
rect 160428 75216 160434 75228
rect 160922 75216 160928 75228
rect 160980 75216 160986 75268
rect 163038 75216 163044 75268
rect 163096 75256 163102 75268
rect 163590 75256 163596 75268
rect 163096 75228 163596 75256
rect 163096 75216 163102 75228
rect 163590 75216 163596 75228
rect 163648 75216 163654 75268
rect 166258 75216 166264 75268
rect 166316 75256 166322 75268
rect 166442 75256 166448 75268
rect 166316 75228 166448 75256
rect 166316 75216 166322 75228
rect 166442 75216 166448 75228
rect 166500 75216 166506 75268
rect 168466 75216 168472 75268
rect 168524 75256 168530 75268
rect 168834 75256 168840 75268
rect 168524 75228 168840 75256
rect 168524 75216 168530 75228
rect 168834 75216 168840 75228
rect 168892 75216 168898 75268
rect 169938 75216 169944 75268
rect 169996 75256 170002 75268
rect 170214 75256 170220 75268
rect 169996 75228 170220 75256
rect 169996 75216 170002 75228
rect 170214 75216 170220 75228
rect 170272 75216 170278 75268
rect 178678 75216 178684 75268
rect 178736 75256 178742 75268
rect 506474 75256 506480 75268
rect 178736 75228 506480 75256
rect 178736 75216 178742 75228
rect 506474 75216 506480 75228
rect 506532 75216 506538 75268
rect 128354 75188 128360 75200
rect 6972 75160 118694 75188
rect 120046 75160 128360 75188
rect 6972 75148 6978 75160
rect 118666 75052 118694 75160
rect 128354 75148 128360 75160
rect 128412 75148 128418 75200
rect 135714 75148 135720 75200
rect 135772 75188 135778 75200
rect 136358 75188 136364 75200
rect 135772 75160 136364 75188
rect 135772 75148 135778 75160
rect 136358 75148 136364 75160
rect 136416 75148 136422 75200
rect 136726 75148 136732 75200
rect 136784 75188 136790 75200
rect 137094 75188 137100 75200
rect 136784 75160 137100 75188
rect 136784 75148 136790 75160
rect 137094 75148 137100 75160
rect 137152 75148 137158 75200
rect 138014 75148 138020 75200
rect 138072 75188 138078 75200
rect 138658 75188 138664 75200
rect 138072 75160 138664 75188
rect 138072 75148 138078 75160
rect 138658 75148 138664 75160
rect 138716 75148 138722 75200
rect 150526 75148 150532 75200
rect 150584 75188 150590 75200
rect 151170 75188 151176 75200
rect 150584 75160 151176 75188
rect 150584 75148 150590 75160
rect 151170 75148 151176 75160
rect 151228 75148 151234 75200
rect 164418 75148 164424 75200
rect 164476 75188 164482 75200
rect 164970 75188 164976 75200
rect 164476 75160 164976 75188
rect 164476 75148 164482 75160
rect 164970 75148 164976 75160
rect 165028 75148 165034 75200
rect 165798 75148 165804 75200
rect 165856 75188 165862 75200
rect 166534 75188 166540 75200
rect 165856 75160 166540 75188
rect 165856 75148 165862 75160
rect 166534 75148 166540 75160
rect 166592 75148 166598 75200
rect 169386 75148 169392 75200
rect 169444 75188 169450 75200
rect 564434 75188 564440 75200
rect 169444 75160 178816 75188
rect 169444 75148 169450 75160
rect 136818 75080 136824 75132
rect 136876 75120 136882 75132
rect 137462 75120 137468 75132
rect 136876 75092 137468 75120
rect 136876 75080 136882 75092
rect 137462 75080 137468 75092
rect 137520 75080 137526 75132
rect 138198 75080 138204 75132
rect 138256 75120 138262 75132
rect 138566 75120 138572 75132
rect 138256 75092 138572 75120
rect 138256 75080 138262 75092
rect 138566 75080 138572 75092
rect 138624 75080 138630 75132
rect 139394 75080 139400 75132
rect 139452 75120 139458 75132
rect 140314 75120 140320 75132
rect 139452 75092 140320 75120
rect 139452 75080 139458 75092
rect 140314 75080 140320 75092
rect 140372 75080 140378 75132
rect 149238 75080 149244 75132
rect 149296 75120 149302 75132
rect 149606 75120 149612 75132
rect 149296 75092 149612 75120
rect 149296 75080 149302 75092
rect 149606 75080 149612 75092
rect 149664 75080 149670 75132
rect 153010 75080 153016 75132
rect 153068 75120 153074 75132
rect 154022 75120 154028 75132
rect 153068 75092 154028 75120
rect 153068 75080 153074 75092
rect 154022 75080 154028 75092
rect 154080 75080 154086 75132
rect 156322 75080 156328 75132
rect 156380 75120 156386 75132
rect 156782 75120 156788 75132
rect 156380 75092 156788 75120
rect 156380 75080 156386 75092
rect 156782 75080 156788 75092
rect 156840 75080 156846 75132
rect 164326 75080 164332 75132
rect 164384 75120 164390 75132
rect 164878 75120 164884 75132
rect 164384 75092 164884 75120
rect 164384 75080 164390 75092
rect 164878 75080 164884 75092
rect 164936 75080 164942 75132
rect 165154 75080 165160 75132
rect 165212 75120 165218 75132
rect 178678 75120 178684 75132
rect 165212 75092 178684 75120
rect 165212 75080 165218 75092
rect 178678 75080 178684 75092
rect 178736 75080 178742 75132
rect 178788 75120 178816 75160
rect 183526 75160 564440 75188
rect 183526 75120 183554 75160
rect 564434 75148 564440 75160
rect 564492 75148 564498 75200
rect 178788 75092 183554 75120
rect 123018 75052 123024 75064
rect 118666 75024 123024 75052
rect 123018 75012 123024 75024
rect 123076 75012 123082 75064
rect 136726 75012 136732 75064
rect 136784 75052 136790 75064
rect 137738 75052 137744 75064
rect 136784 75024 137744 75052
rect 136784 75012 136790 75024
rect 137738 75012 137744 75024
rect 137796 75012 137802 75064
rect 167086 75012 167092 75064
rect 167144 75052 167150 75064
rect 167546 75052 167552 75064
rect 167144 75024 167552 75052
rect 167144 75012 167150 75024
rect 167546 75012 167552 75024
rect 167604 75012 167610 75064
rect 168466 75012 168472 75064
rect 168524 75052 168530 75064
rect 169110 75052 169116 75064
rect 168524 75024 169116 75052
rect 168524 75012 168530 75024
rect 169110 75012 169116 75024
rect 169168 75012 169174 75064
rect 169754 75012 169760 75064
rect 169812 75052 169818 75064
rect 170214 75052 170220 75064
rect 169812 75024 170220 75052
rect 169812 75012 169818 75024
rect 170214 75012 170220 75024
rect 170272 75012 170278 75064
rect 120810 74944 120816 74996
rect 120868 74984 120874 74996
rect 128538 74984 128544 74996
rect 120868 74956 128544 74984
rect 120868 74944 120874 74956
rect 128538 74944 128544 74956
rect 128596 74944 128602 74996
rect 138198 74944 138204 74996
rect 138256 74984 138262 74996
rect 138750 74984 138756 74996
rect 138256 74956 138756 74984
rect 138256 74944 138262 74956
rect 138750 74944 138756 74956
rect 138808 74944 138814 74996
rect 149606 74944 149612 74996
rect 149664 74984 149670 74996
rect 149974 74984 149980 74996
rect 149664 74956 149980 74984
rect 149664 74944 149670 74956
rect 149974 74944 149980 74956
rect 150032 74944 150038 74996
rect 167086 74876 167092 74928
rect 167144 74916 167150 74928
rect 167822 74916 167828 74928
rect 167144 74888 167828 74916
rect 167144 74876 167150 74888
rect 167822 74876 167828 74888
rect 167880 74876 167886 74928
rect 169754 74876 169760 74928
rect 169812 74916 169818 74928
rect 170490 74916 170496 74928
rect 169812 74888 170496 74916
rect 169812 74876 169818 74888
rect 170490 74876 170496 74888
rect 170548 74876 170554 74928
rect 154666 74672 154672 74724
rect 154724 74712 154730 74724
rect 155494 74712 155500 74724
rect 154724 74684 155500 74712
rect 154724 74672 154730 74684
rect 155494 74672 155500 74684
rect 155552 74672 155558 74724
rect 134610 74468 134616 74520
rect 134668 74508 134674 74520
rect 135346 74508 135352 74520
rect 134668 74480 135352 74508
rect 134668 74468 134674 74480
rect 135346 74468 135352 74480
rect 135404 74468 135410 74520
rect 126238 74264 126244 74316
rect 126296 74304 126302 74316
rect 129550 74304 129556 74316
rect 126296 74276 129556 74304
rect 126296 74264 126302 74276
rect 129550 74264 129556 74276
rect 129608 74264 129614 74316
rect 137922 74264 137928 74316
rect 137980 74304 137986 74316
rect 142890 74304 142896 74316
rect 137980 74276 142896 74304
rect 137980 74264 137986 74276
rect 142890 74264 142896 74276
rect 142948 74264 142954 74316
rect 164050 74128 164056 74180
rect 164108 74168 164114 74180
rect 173434 74168 173440 74180
rect 164108 74140 173440 74168
rect 164108 74128 164114 74140
rect 173434 74128 173440 74140
rect 173492 74128 173498 74180
rect 139210 74060 139216 74112
rect 139268 74100 139274 74112
rect 173894 74100 173900 74112
rect 139268 74072 173900 74100
rect 139268 74060 139274 74072
rect 173894 74060 173900 74072
rect 173952 74060 173958 74112
rect 122834 73992 122840 74044
rect 122892 74032 122898 74044
rect 135070 74032 135076 74044
rect 122892 74004 135076 74032
rect 122892 73992 122898 74004
rect 135070 73992 135076 74004
rect 135128 73992 135134 74044
rect 141970 73992 141976 74044
rect 142028 74032 142034 74044
rect 209774 74032 209780 74044
rect 142028 74004 209780 74032
rect 142028 73992 142034 74004
rect 209774 73992 209780 74004
rect 209832 73992 209838 74044
rect 93946 73924 93952 73976
rect 94004 73964 94010 73976
rect 133230 73964 133236 73976
rect 94004 73936 133236 73964
rect 94004 73924 94010 73936
rect 133230 73924 133236 73936
rect 133288 73924 133294 73976
rect 142982 73924 142988 73976
rect 143040 73964 143046 73976
rect 223574 73964 223580 73976
rect 143040 73936 223580 73964
rect 143040 73924 143046 73936
rect 223574 73924 223580 73936
rect 223632 73924 223638 73976
rect 51074 73856 51080 73908
rect 51132 73896 51138 73908
rect 129458 73896 129464 73908
rect 51132 73868 129464 73896
rect 51132 73856 51138 73868
rect 129458 73856 129464 73868
rect 129516 73856 129522 73908
rect 147306 73856 147312 73908
rect 147364 73896 147370 73908
rect 251174 73896 251180 73908
rect 147364 73868 251180 73896
rect 147364 73856 147370 73868
rect 251174 73856 251180 73868
rect 251232 73856 251238 73908
rect 4798 73788 4804 73840
rect 4856 73828 4862 73840
rect 125226 73828 125232 73840
rect 4856 73800 125232 73828
rect 4856 73788 4862 73800
rect 125226 73788 125232 73800
rect 125284 73788 125290 73840
rect 155310 73788 155316 73840
rect 155368 73828 155374 73840
rect 357434 73828 357440 73840
rect 155368 73800 357440 73828
rect 155368 73788 155374 73800
rect 357434 73788 357440 73800
rect 357492 73788 357498 73840
rect 124766 73652 124772 73704
rect 124824 73692 124830 73704
rect 125226 73692 125232 73704
rect 124824 73664 125232 73692
rect 124824 73652 124830 73664
rect 125226 73652 125232 73664
rect 125284 73652 125290 73704
rect 161474 73380 161480 73432
rect 161532 73420 161538 73432
rect 161842 73420 161848 73432
rect 161532 73392 161848 73420
rect 161532 73380 161538 73392
rect 161842 73380 161848 73392
rect 161900 73380 161906 73432
rect 125042 73312 125048 73364
rect 125100 73352 125106 73364
rect 127986 73352 127992 73364
rect 125100 73324 127992 73352
rect 125100 73312 125106 73324
rect 127986 73312 127992 73324
rect 128044 73312 128050 73364
rect 161842 73244 161848 73296
rect 161900 73284 161906 73296
rect 162302 73284 162308 73296
rect 161900 73256 162308 73284
rect 161900 73244 161906 73256
rect 162302 73244 162308 73256
rect 162360 73244 162366 73296
rect 171134 73108 171140 73160
rect 171192 73148 171198 73160
rect 580166 73148 580172 73160
rect 171192 73120 580172 73148
rect 171192 73108 171198 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 126146 73040 126152 73092
rect 126204 73080 126210 73092
rect 126698 73080 126704 73092
rect 126204 73052 126704 73080
rect 126204 73040 126210 73052
rect 126698 73040 126704 73052
rect 126756 73040 126762 73092
rect 163774 72904 163780 72956
rect 163832 72944 163838 72956
rect 173526 72944 173532 72956
rect 163832 72916 173532 72944
rect 163832 72904 163838 72916
rect 173526 72904 173532 72916
rect 173584 72904 173590 72956
rect 162026 72836 162032 72888
rect 162084 72876 162090 72888
rect 181438 72876 181444 72888
rect 162084 72848 181444 72876
rect 162084 72836 162090 72848
rect 181438 72836 181444 72848
rect 181496 72836 181502 72888
rect 114554 72768 114560 72820
rect 114612 72808 114618 72820
rect 133414 72808 133420 72820
rect 114612 72780 133420 72808
rect 114612 72768 114618 72780
rect 133414 72768 133420 72780
rect 133472 72768 133478 72820
rect 151078 72768 151084 72820
rect 151136 72808 151142 72820
rect 325694 72808 325700 72820
rect 151136 72780 325700 72808
rect 151136 72768 151142 72780
rect 325694 72768 325700 72780
rect 325752 72768 325758 72820
rect 103514 72700 103520 72752
rect 103572 72740 103578 72752
rect 133598 72740 133604 72752
rect 103572 72712 133604 72740
rect 103572 72700 103578 72712
rect 133598 72700 133604 72712
rect 133656 72700 133662 72752
rect 151446 72700 151452 72752
rect 151504 72740 151510 72752
rect 332594 72740 332600 72752
rect 151504 72712 332600 72740
rect 151504 72700 151510 72712
rect 332594 72700 332600 72712
rect 332652 72700 332658 72752
rect 69014 72632 69020 72684
rect 69072 72672 69078 72684
rect 130654 72672 130660 72684
rect 69072 72644 130660 72672
rect 69072 72632 69078 72644
rect 130654 72632 130660 72644
rect 130712 72632 130718 72684
rect 151998 72632 152004 72684
rect 152056 72672 152062 72684
rect 340874 72672 340880 72684
rect 152056 72644 340880 72672
rect 152056 72632 152062 72644
rect 340874 72632 340880 72644
rect 340932 72632 340938 72684
rect 341518 72632 341524 72684
rect 341576 72672 341582 72684
rect 465074 72672 465080 72684
rect 341576 72644 465080 72672
rect 341576 72632 341582 72644
rect 465074 72632 465080 72644
rect 465132 72632 465138 72684
rect 26234 72564 26240 72616
rect 26292 72604 26298 72616
rect 127434 72604 127440 72616
rect 26292 72576 127440 72604
rect 26292 72564 26298 72576
rect 127434 72564 127440 72576
rect 127492 72564 127498 72616
rect 152734 72564 152740 72616
rect 152792 72604 152798 72616
rect 347774 72604 347780 72616
rect 152792 72576 347780 72604
rect 152792 72564 152798 72576
rect 347774 72564 347780 72576
rect 347832 72564 347838 72616
rect 13814 72496 13820 72548
rect 13872 72536 13878 72548
rect 123202 72536 123208 72548
rect 13872 72508 123208 72536
rect 13872 72496 13878 72508
rect 123202 72496 123208 72508
rect 123260 72496 123266 72548
rect 157978 72496 157984 72548
rect 158036 72536 158042 72548
rect 368474 72536 368480 72548
rect 158036 72508 368480 72536
rect 158036 72496 158042 72508
rect 368474 72496 368480 72508
rect 368532 72496 368538 72548
rect 11054 72428 11060 72480
rect 11112 72468 11118 72480
rect 126606 72468 126612 72480
rect 11112 72440 126612 72468
rect 11112 72428 11118 72440
rect 126606 72428 126612 72440
rect 126664 72428 126670 72480
rect 127434 72428 127440 72480
rect 127492 72468 127498 72480
rect 128078 72468 128084 72480
rect 127492 72440 128084 72468
rect 127492 72428 127498 72440
rect 128078 72428 128084 72440
rect 128136 72428 128142 72480
rect 159450 72428 159456 72480
rect 159508 72468 159514 72480
rect 382274 72468 382280 72480
rect 159508 72440 382280 72468
rect 159508 72428 159514 72440
rect 382274 72428 382280 72440
rect 382332 72428 382338 72480
rect 124950 72224 124956 72276
rect 125008 72264 125014 72276
rect 125686 72264 125692 72276
rect 125008 72236 125692 72264
rect 125008 72224 125014 72236
rect 125686 72224 125692 72236
rect 125744 72224 125750 72276
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 97258 71720 97264 71732
rect 3476 71692 97264 71720
rect 3476 71680 3482 71692
rect 97258 71680 97264 71692
rect 97316 71680 97322 71732
rect 132678 71680 132684 71732
rect 132736 71720 132742 71732
rect 135990 71720 135996 71732
rect 132736 71692 135996 71720
rect 132736 71680 132742 71692
rect 135990 71680 135996 71692
rect 136048 71680 136054 71732
rect 140590 71340 140596 71392
rect 140648 71380 140654 71392
rect 176746 71380 176752 71392
rect 140648 71352 176752 71380
rect 140648 71340 140654 71352
rect 176746 71340 176752 71352
rect 176804 71340 176810 71392
rect 121454 71272 121460 71324
rect 121512 71312 121518 71324
rect 134886 71312 134892 71324
rect 121512 71284 134892 71312
rect 121512 71272 121518 71284
rect 134886 71272 134892 71284
rect 134944 71272 134950 71324
rect 155586 71272 155592 71324
rect 155644 71312 155650 71324
rect 367094 71312 367100 71324
rect 155644 71284 367100 71312
rect 155644 71272 155650 71284
rect 367094 71272 367100 71284
rect 367152 71272 367158 71324
rect 100754 71204 100760 71256
rect 100812 71244 100818 71256
rect 133506 71244 133512 71256
rect 100812 71216 133512 71244
rect 100812 71204 100818 71216
rect 133506 71204 133512 71216
rect 133564 71204 133570 71256
rect 155218 71204 155224 71256
rect 155276 71244 155282 71256
rect 382366 71244 382372 71256
rect 155276 71216 382372 71244
rect 155276 71204 155282 71216
rect 382366 71204 382372 71216
rect 382424 71204 382430 71256
rect 96614 71136 96620 71188
rect 96672 71176 96678 71188
rect 133322 71176 133328 71188
rect 96672 71148 133328 71176
rect 96672 71136 96678 71148
rect 133322 71136 133328 71148
rect 133380 71136 133386 71188
rect 165246 71136 165252 71188
rect 165304 71176 165310 71188
rect 505094 71176 505100 71188
rect 165304 71148 505100 71176
rect 165304 71136 165310 71148
rect 505094 71136 505100 71148
rect 505152 71136 505158 71188
rect 49694 71068 49700 71120
rect 49752 71108 49758 71120
rect 126974 71108 126980 71120
rect 49752 71080 126980 71108
rect 49752 71068 49758 71080
rect 126974 71068 126980 71080
rect 127032 71068 127038 71120
rect 166626 71068 166632 71120
rect 166684 71108 166690 71120
rect 518894 71108 518900 71120
rect 166684 71080 518900 71108
rect 166684 71068 166690 71080
rect 518894 71068 518900 71080
rect 518952 71068 518958 71120
rect 28994 71000 29000 71052
rect 29052 71040 29058 71052
rect 128262 71040 128268 71052
rect 29052 71012 128268 71040
rect 29052 71000 29058 71012
rect 128262 71000 128268 71012
rect 128320 71000 128326 71052
rect 168282 71000 168288 71052
rect 168340 71040 168346 71052
rect 539594 71040 539600 71052
rect 168340 71012 539600 71040
rect 168340 71000 168346 71012
rect 539594 71000 539600 71012
rect 539652 71000 539658 71052
rect 137278 70388 137284 70440
rect 137336 70428 137342 70440
rect 138750 70428 138756 70440
rect 137336 70400 138756 70428
rect 137336 70388 137342 70400
rect 138750 70388 138756 70400
rect 138808 70388 138814 70440
rect 140038 70184 140044 70236
rect 140096 70224 140102 70236
rect 184934 70224 184940 70236
rect 140096 70196 184940 70224
rect 140096 70184 140102 70196
rect 184934 70184 184940 70196
rect 184992 70184 184998 70236
rect 141510 70116 141516 70168
rect 141568 70156 141574 70168
rect 209866 70156 209872 70168
rect 141568 70128 209872 70156
rect 141568 70116 141574 70128
rect 209866 70116 209872 70128
rect 209924 70116 209930 70168
rect 3418 70048 3424 70100
rect 3476 70088 3482 70100
rect 174538 70088 174544 70100
rect 3476 70060 174544 70088
rect 3476 70048 3482 70060
rect 174538 70048 174544 70060
rect 174596 70048 174602 70100
rect 162394 69980 162400 70032
rect 162452 70020 162458 70032
rect 375374 70020 375380 70032
rect 162452 69992 375380 70020
rect 162452 69980 162458 69992
rect 375374 69980 375380 69992
rect 375432 69980 375438 70032
rect 159358 69912 159364 69964
rect 159416 69952 159422 69964
rect 437474 69952 437480 69964
rect 159416 69924 437480 69952
rect 159416 69912 159422 69924
rect 437474 69912 437480 69924
rect 437532 69912 437538 69964
rect 82814 69844 82820 69896
rect 82872 69884 82878 69896
rect 131482 69884 131488 69896
rect 82872 69856 131488 69884
rect 82872 69844 82878 69856
rect 131482 69844 131488 69856
rect 131540 69844 131546 69896
rect 166350 69844 166356 69896
rect 166408 69884 166414 69896
rect 523034 69884 523040 69896
rect 166408 69856 523040 69884
rect 166408 69844 166414 69856
rect 523034 69844 523040 69856
rect 523092 69844 523098 69896
rect 78674 69776 78680 69828
rect 78732 69816 78738 69828
rect 131206 69816 131212 69828
rect 78732 69788 131212 69816
rect 78732 69776 78738 69788
rect 131206 69776 131212 69788
rect 131264 69776 131270 69828
rect 167730 69776 167736 69828
rect 167788 69816 167794 69828
rect 536834 69816 536840 69828
rect 167788 69788 536840 69816
rect 167788 69776 167794 69788
rect 536834 69776 536840 69788
rect 536892 69776 536898 69828
rect 52454 69708 52460 69760
rect 52512 69748 52518 69760
rect 128814 69748 128820 69760
rect 52512 69720 128820 69748
rect 52512 69708 52518 69720
rect 128814 69708 128820 69720
rect 128872 69708 128878 69760
rect 170766 69708 170772 69760
rect 170824 69748 170830 69760
rect 558914 69748 558920 69760
rect 170824 69720 558920 69748
rect 170824 69708 170830 69720
rect 558914 69708 558920 69720
rect 558972 69708 558978 69760
rect 33134 69640 33140 69692
rect 33192 69680 33198 69692
rect 127434 69680 127440 69692
rect 33192 69652 127440 69680
rect 33192 69640 33198 69652
rect 127434 69640 127440 69652
rect 127492 69640 127498 69692
rect 169478 69640 169484 69692
rect 169536 69680 169542 69692
rect 564526 69680 564532 69692
rect 169536 69652 564532 69680
rect 169536 69640 169542 69652
rect 564526 69640 564532 69652
rect 564584 69640 564590 69692
rect 137186 68960 137192 69012
rect 137244 69000 137250 69012
rect 138842 69000 138848 69012
rect 137244 68972 138848 69000
rect 137244 68960 137250 68972
rect 138842 68960 138848 68972
rect 138900 68960 138906 69012
rect 138658 68824 138664 68876
rect 138716 68864 138722 68876
rect 171134 68864 171140 68876
rect 138716 68836 171140 68864
rect 138716 68824 138722 68836
rect 171134 68824 171140 68836
rect 171192 68824 171198 68876
rect 141418 68756 141424 68808
rect 141476 68796 141482 68808
rect 202874 68796 202880 68808
rect 141476 68768 202880 68796
rect 141476 68756 141482 68768
rect 202874 68756 202880 68768
rect 202932 68756 202938 68808
rect 157058 68688 157064 68740
rect 157116 68728 157122 68740
rect 249794 68728 249800 68740
rect 157116 68700 249800 68728
rect 157116 68688 157122 68700
rect 249794 68688 249800 68700
rect 249852 68688 249858 68740
rect 18598 68620 18604 68672
rect 18656 68660 18662 68672
rect 183002 68660 183008 68672
rect 18656 68632 183008 68660
rect 18656 68620 18662 68632
rect 183002 68620 183008 68632
rect 183060 68620 183066 68672
rect 150986 68552 150992 68604
rect 151044 68592 151050 68604
rect 332686 68592 332692 68604
rect 151044 68564 332692 68592
rect 151044 68552 151050 68564
rect 332686 68552 332692 68564
rect 332744 68552 332750 68604
rect 159266 68484 159272 68536
rect 159324 68524 159330 68536
rect 431954 68524 431960 68536
rect 159324 68496 431960 68524
rect 159324 68484 159330 68496
rect 431954 68484 431960 68496
rect 432012 68484 432018 68536
rect 115934 68416 115940 68468
rect 115992 68456 115998 68468
rect 134242 68456 134248 68468
rect 115992 68428 134248 68456
rect 115992 68416 115998 68428
rect 134242 68416 134248 68428
rect 134300 68416 134306 68468
rect 163498 68416 163504 68468
rect 163556 68456 163562 68468
rect 481634 68456 481640 68468
rect 163556 68428 481640 68456
rect 163556 68416 163562 68428
rect 481634 68416 481640 68428
rect 481692 68416 481698 68468
rect 85574 68348 85580 68400
rect 85632 68388 85638 68400
rect 132126 68388 132132 68400
rect 85632 68360 132132 68388
rect 85632 68348 85638 68360
rect 132126 68348 132132 68360
rect 132184 68348 132190 68400
rect 167638 68348 167644 68400
rect 167696 68388 167702 68400
rect 543734 68388 543740 68400
rect 167696 68360 543740 68388
rect 167696 68348 167702 68360
rect 543734 68348 543740 68360
rect 543792 68348 543798 68400
rect 59354 68280 59360 68332
rect 59412 68320 59418 68332
rect 129826 68320 129832 68332
rect 59412 68292 129832 68320
rect 59412 68280 59418 68292
rect 129826 68280 129832 68292
rect 129884 68280 129890 68332
rect 170582 68280 170588 68332
rect 170640 68320 170646 68332
rect 550634 68320 550640 68332
rect 170640 68292 550640 68320
rect 170640 68280 170646 68292
rect 550634 68280 550640 68292
rect 550692 68280 550698 68332
rect 139946 67124 139952 67176
rect 140004 67164 140010 67176
rect 189074 67164 189080 67176
rect 140004 67136 189080 67164
rect 140004 67124 140010 67136
rect 189074 67124 189080 67136
rect 189132 67124 189138 67176
rect 141326 67056 141332 67108
rect 141384 67096 141390 67108
rect 207014 67096 207020 67108
rect 141384 67068 207020 67096
rect 141384 67056 141390 67068
rect 207014 67056 207020 67068
rect 207072 67056 207078 67108
rect 153746 66988 153752 67040
rect 153804 67028 153810 67040
rect 356054 67028 356060 67040
rect 153804 67000 356060 67028
rect 153804 66988 153810 67000
rect 356054 66988 356060 67000
rect 356112 66988 356118 67040
rect 64874 66920 64880 66972
rect 64932 66960 64938 66972
rect 130194 66960 130200 66972
rect 64932 66932 130200 66960
rect 64932 66920 64938 66932
rect 130194 66920 130200 66932
rect 130252 66920 130258 66972
rect 155126 66920 155132 66972
rect 155184 66960 155190 66972
rect 374086 66960 374092 66972
rect 155184 66932 374092 66960
rect 155184 66920 155190 66932
rect 374086 66920 374092 66932
rect 374144 66920 374150 66972
rect 16574 66852 16580 66904
rect 16632 66892 16638 66904
rect 126146 66892 126152 66904
rect 16632 66864 126152 66892
rect 16632 66852 16638 66864
rect 126146 66852 126152 66864
rect 126204 66852 126210 66904
rect 166258 66852 166264 66904
rect 166316 66892 166322 66904
rect 525794 66892 525800 66904
rect 166316 66864 525800 66892
rect 166316 66852 166322 66864
rect 525794 66852 525800 66864
rect 525852 66852 525858 66904
rect 138566 66172 138572 66224
rect 138624 66212 138630 66224
rect 140130 66212 140136 66224
rect 138624 66184 140136 66212
rect 138624 66172 138630 66184
rect 140130 66172 140136 66184
rect 140188 66172 140194 66224
rect 148318 65696 148324 65748
rect 148376 65736 148382 65748
rect 292574 65736 292580 65748
rect 148376 65708 292580 65736
rect 148376 65696 148382 65708
rect 292574 65696 292580 65708
rect 292632 65696 292638 65748
rect 156598 65628 156604 65680
rect 156656 65668 156662 65680
rect 390554 65668 390560 65680
rect 156656 65640 390560 65668
rect 156656 65628 156662 65640
rect 390554 65628 390560 65640
rect 390612 65628 390618 65680
rect 158346 65560 158352 65612
rect 158404 65600 158410 65612
rect 396074 65600 396080 65612
rect 158404 65572 396080 65600
rect 158404 65560 158410 65572
rect 396074 65560 396080 65572
rect 396132 65560 396138 65612
rect 170214 65492 170220 65544
rect 170272 65532 170278 65544
rect 568574 65532 568580 65544
rect 170272 65504 568580 65532
rect 170272 65492 170278 65504
rect 568574 65492 568580 65504
rect 568632 65492 568638 65544
rect 120074 64880 120080 64932
rect 120132 64920 120138 64932
rect 123662 64920 123668 64932
rect 120132 64892 123668 64920
rect 120132 64880 120138 64892
rect 123662 64880 123668 64892
rect 123720 64880 123726 64932
rect 145558 64336 145564 64388
rect 145616 64376 145622 64388
rect 256694 64376 256700 64388
rect 145616 64348 256700 64376
rect 145616 64336 145622 64348
rect 256694 64336 256700 64348
rect 256752 64336 256758 64388
rect 157978 64268 157984 64320
rect 158036 64308 158042 64320
rect 412634 64308 412640 64320
rect 158036 64280 412640 64308
rect 158036 64268 158042 64280
rect 412634 64268 412640 64280
rect 412692 64268 412698 64320
rect 160830 64200 160836 64252
rect 160888 64240 160894 64252
rect 444374 64240 444380 64252
rect 160888 64212 444380 64240
rect 160888 64200 160894 64212
rect 444374 64200 444380 64212
rect 444432 64200 444438 64252
rect 169018 64132 169024 64184
rect 169076 64172 169082 64184
rect 561674 64172 561680 64184
rect 169076 64144 561680 64172
rect 169076 64132 169082 64144
rect 561674 64132 561680 64144
rect 561732 64132 561738 64184
rect 148686 62908 148692 62960
rect 148744 62948 148750 62960
rect 190454 62948 190460 62960
rect 148744 62920 190460 62948
rect 148744 62908 148750 62920
rect 190454 62908 190460 62920
rect 190512 62908 190518 62960
rect 157886 62840 157892 62892
rect 157944 62880 157950 62892
rect 408494 62880 408500 62892
rect 157944 62852 408500 62880
rect 157944 62840 157950 62852
rect 408494 62840 408500 62852
rect 408552 62840 408558 62892
rect 159174 62772 159180 62824
rect 159232 62812 159238 62824
rect 440234 62812 440240 62824
rect 159232 62784 440240 62812
rect 159232 62772 159238 62784
rect 440234 62772 440240 62784
rect 440292 62772 440298 62824
rect 145466 61548 145472 61600
rect 145524 61588 145530 61600
rect 259454 61588 259460 61600
rect 145524 61560 259460 61588
rect 145524 61548 145530 61560
rect 259454 61548 259460 61560
rect 259512 61548 259518 61600
rect 155034 61480 155040 61532
rect 155092 61520 155098 61532
rect 380894 61520 380900 61532
rect 155092 61492 380900 61520
rect 155092 61480 155098 61492
rect 380894 61480 380900 61492
rect 380952 61480 380958 61532
rect 163406 61412 163412 61464
rect 163464 61452 163470 61464
rect 481726 61452 481732 61464
rect 163464 61424 481732 61452
rect 163464 61412 163470 61424
rect 481726 61412 481732 61424
rect 481784 61412 481790 61464
rect 118326 61344 118332 61396
rect 118384 61384 118390 61396
rect 580258 61384 580264 61396
rect 118384 61356 580264 61384
rect 118384 61344 118390 61356
rect 580258 61344 580264 61356
rect 580316 61344 580322 61396
rect 138474 60664 138480 60716
rect 138532 60704 138538 60716
rect 144270 60704 144276 60716
rect 138532 60676 144276 60704
rect 138532 60664 138538 60676
rect 144270 60664 144276 60676
rect 144328 60664 144334 60716
rect 182818 60664 182824 60716
rect 182876 60704 182882 60716
rect 580166 60704 580172 60716
rect 182876 60676 580172 60704
rect 182876 60664 182882 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 139762 60256 139768 60308
rect 139820 60296 139826 60308
rect 179506 60296 179512 60308
rect 139820 60268 179512 60296
rect 139820 60256 139826 60268
rect 179506 60256 179512 60268
rect 179564 60256 179570 60308
rect 139854 60188 139860 60240
rect 139912 60228 139918 60240
rect 183554 60228 183560 60240
rect 139912 60200 183560 60228
rect 139912 60188 139918 60200
rect 183554 60188 183560 60200
rect 183612 60188 183618 60240
rect 148226 60120 148232 60172
rect 148284 60160 148290 60172
rect 295334 60160 295340 60172
rect 148284 60132 295340 60160
rect 148284 60120 148290 60132
rect 295334 60120 295340 60132
rect 295392 60120 295398 60172
rect 154942 60052 154948 60104
rect 155000 60092 155006 60104
rect 376754 60092 376760 60104
rect 155000 60064 376760 60092
rect 155000 60052 155006 60064
rect 376754 60052 376760 60064
rect 376812 60052 376818 60104
rect 102226 59984 102232 60036
rect 102284 60024 102290 60036
rect 125410 60024 125416 60036
rect 102284 59996 125416 60024
rect 102284 59984 102290 59996
rect 125410 59984 125416 59996
rect 125468 59984 125474 60036
rect 161106 59984 161112 60036
rect 161164 60024 161170 60036
rect 390646 60024 390652 60036
rect 161164 59996 390652 60024
rect 161164 59984 161170 59996
rect 390646 59984 390652 59996
rect 390704 59984 390710 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 18598 59344 18604 59356
rect 3108 59316 18604 59344
rect 3108 59304 3114 59316
rect 18598 59304 18604 59316
rect 18656 59304 18662 59356
rect 137094 59304 137100 59356
rect 137152 59344 137158 59356
rect 140222 59344 140228 59356
rect 137152 59316 140228 59344
rect 137152 59304 137158 59316
rect 140222 59304 140228 59316
rect 140280 59304 140286 59356
rect 139670 58964 139676 59016
rect 139728 59004 139734 59016
rect 180794 59004 180800 59016
rect 139728 58976 180800 59004
rect 139728 58964 139734 58976
rect 180794 58964 180800 58976
rect 180852 58964 180858 59016
rect 150894 58896 150900 58948
rect 150952 58936 150958 58948
rect 327074 58936 327080 58948
rect 150952 58908 327080 58936
rect 150952 58896 150958 58908
rect 327074 58896 327080 58908
rect 327132 58896 327138 58948
rect 153654 58828 153660 58880
rect 153712 58868 153718 58880
rect 358814 58868 358820 58880
rect 153712 58840 358820 58868
rect 153712 58828 153718 58840
rect 358814 58828 358820 58840
rect 358872 58828 358878 58880
rect 159082 58760 159088 58812
rect 159140 58800 159146 58812
rect 433334 58800 433340 58812
rect 159140 58772 433340 58800
rect 159140 58760 159146 58772
rect 433334 58760 433340 58772
rect 433392 58760 433398 58812
rect 164786 58692 164792 58744
rect 164844 58732 164850 58744
rect 507854 58732 507860 58744
rect 164844 58704 507860 58732
rect 164844 58692 164850 58704
rect 507854 58692 507860 58704
rect 507912 58692 507918 58744
rect 170122 58624 170128 58676
rect 170180 58664 170186 58676
rect 572714 58664 572720 58676
rect 170180 58636 572720 58664
rect 170180 58624 170186 58636
rect 572714 58624 572720 58636
rect 572772 58624 572778 58676
rect 141234 57264 141240 57316
rect 141292 57304 141298 57316
rect 201494 57304 201500 57316
rect 141292 57276 201500 57304
rect 141292 57264 141298 57276
rect 201494 57264 201500 57276
rect 201552 57264 201558 57316
rect 156506 57196 156512 57248
rect 156564 57236 156570 57248
rect 394694 57236 394700 57248
rect 156564 57208 394700 57236
rect 156564 57196 156570 57208
rect 394694 57196 394700 57208
rect 394752 57196 394758 57248
rect 150802 55904 150808 55956
rect 150860 55944 150866 55956
rect 331214 55944 331220 55956
rect 150860 55916 331220 55944
rect 150860 55904 150866 55916
rect 331214 55904 331220 55916
rect 331272 55904 331278 55956
rect 95234 55836 95240 55888
rect 95292 55876 95298 55888
rect 125318 55876 125324 55888
rect 95292 55848 125324 55876
rect 95292 55836 95298 55848
rect 125318 55836 125324 55848
rect 125376 55836 125382 55888
rect 154850 55836 154856 55888
rect 154908 55876 154914 55888
rect 383654 55876 383660 55888
rect 154908 55848 383660 55876
rect 154908 55836 154914 55848
rect 383654 55836 383660 55848
rect 383712 55836 383718 55888
rect 142706 54680 142712 54732
rect 142764 54720 142770 54732
rect 219434 54720 219440 54732
rect 142764 54692 219440 54720
rect 142764 54680 142770 54692
rect 219434 54680 219440 54692
rect 219492 54680 219498 54732
rect 152366 54612 152372 54664
rect 152424 54652 152430 54664
rect 349154 54652 349160 54664
rect 152424 54624 349160 54652
rect 152424 54612 152430 54624
rect 349154 54612 349160 54624
rect 349212 54612 349218 54664
rect 153562 54544 153568 54596
rect 153620 54584 153626 54596
rect 362954 54584 362960 54596
rect 153620 54556 362960 54584
rect 153620 54544 153626 54556
rect 362954 54544 362960 54556
rect 363012 54544 363018 54596
rect 156414 54476 156420 54528
rect 156472 54516 156478 54528
rect 398834 54516 398840 54528
rect 156472 54488 398840 54516
rect 156472 54476 156478 54488
rect 398834 54476 398840 54488
rect 398892 54476 398898 54528
rect 139578 53252 139584 53304
rect 139636 53292 139642 53304
rect 185026 53292 185032 53304
rect 139636 53264 185032 53292
rect 139636 53252 139642 53264
rect 185026 53252 185032 53264
rect 185084 53252 185090 53304
rect 160738 53184 160744 53236
rect 160796 53224 160802 53236
rect 455414 53224 455420 53236
rect 160796 53196 455420 53224
rect 160796 53184 160802 53196
rect 455414 53184 455420 53196
rect 455472 53184 455478 53236
rect 163314 53116 163320 53168
rect 163372 53156 163378 53168
rect 488534 53156 488540 53168
rect 163372 53128 488540 53156
rect 163372 53116 163378 53128
rect 488534 53116 488540 53128
rect 488592 53116 488598 53168
rect 166166 53048 166172 53100
rect 166224 53088 166230 53100
rect 516134 53088 516140 53100
rect 166224 53060 516140 53088
rect 166224 53048 166230 53060
rect 516134 53048 516140 53060
rect 516192 53048 516198 53100
rect 135806 52980 135812 53032
rect 135864 53020 135870 53032
rect 140314 53020 140320 53032
rect 135864 52992 140320 53020
rect 135864 52980 135870 52992
rect 140314 52980 140320 52992
rect 140372 52980 140378 53032
rect 141142 51824 141148 51876
rect 141200 51864 141206 51876
rect 204254 51864 204260 51876
rect 141200 51836 204260 51864
rect 141200 51824 141206 51836
rect 204254 51824 204260 51836
rect 204312 51824 204318 51876
rect 153470 51756 153476 51808
rect 153528 51796 153534 51808
rect 365714 51796 365720 51808
rect 153528 51768 365720 51796
rect 153528 51756 153534 51768
rect 365714 51756 365720 51768
rect 365772 51756 365778 51808
rect 157794 51688 157800 51740
rect 157852 51728 157858 51740
rect 415394 51728 415400 51740
rect 157852 51700 415400 51728
rect 157852 51688 157858 51700
rect 415394 51688 415400 51700
rect 415452 51688 415458 51740
rect 154022 50668 154028 50720
rect 154080 50708 154086 50720
rect 353294 50708 353300 50720
rect 154080 50680 353300 50708
rect 154080 50668 154086 50680
rect 353294 50668 353300 50680
rect 353352 50668 353358 50720
rect 156322 50600 156328 50652
rect 156380 50640 156386 50652
rect 401594 50640 401600 50652
rect 156380 50612 401600 50640
rect 156380 50600 156386 50612
rect 401594 50600 401600 50612
rect 401652 50600 401658 50652
rect 160646 50532 160652 50584
rect 160704 50572 160710 50584
rect 448514 50572 448520 50584
rect 160704 50544 448520 50572
rect 160704 50532 160710 50544
rect 448514 50532 448520 50544
rect 448572 50532 448578 50584
rect 167546 50464 167552 50516
rect 167604 50504 167610 50516
rect 534074 50504 534080 50516
rect 167604 50476 534080 50504
rect 167604 50464 167610 50476
rect 534074 50464 534080 50476
rect 534132 50464 534138 50516
rect 167454 50396 167460 50448
rect 167512 50436 167518 50448
rect 542354 50436 542360 50448
rect 167512 50408 542360 50436
rect 167512 50396 167518 50408
rect 542354 50396 542360 50408
rect 542412 50396 542418 50448
rect 168926 50328 168932 50380
rect 168984 50368 168990 50380
rect 557534 50368 557540 50380
rect 168984 50340 557540 50368
rect 168984 50328 168990 50340
rect 557534 50328 557540 50340
rect 557592 50328 557598 50380
rect 145374 49240 145380 49292
rect 145432 49280 145438 49292
rect 259546 49280 259552 49292
rect 145432 49252 259552 49280
rect 145432 49240 145438 49252
rect 259546 49240 259552 49252
rect 259604 49240 259610 49292
rect 156966 49172 156972 49224
rect 157024 49212 157030 49224
rect 389174 49212 389180 49224
rect 157024 49184 389180 49212
rect 157024 49172 157030 49184
rect 389174 49172 389180 49184
rect 389232 49172 389238 49224
rect 171686 49104 171692 49156
rect 171744 49144 171750 49156
rect 425054 49144 425060 49156
rect 171744 49116 425060 49144
rect 171744 49104 171750 49116
rect 425054 49104 425060 49116
rect 425112 49104 425118 49156
rect 164694 49036 164700 49088
rect 164752 49076 164758 49088
rect 498286 49076 498292 49088
rect 164752 49048 498292 49076
rect 164752 49036 164758 49048
rect 498286 49036 498292 49048
rect 498344 49036 498350 49088
rect 168834 48968 168840 49020
rect 168892 49008 168898 49020
rect 552014 49008 552020 49020
rect 168892 48980 552020 49008
rect 168892 48968 168898 48980
rect 552014 48968 552020 48980
rect 552072 48968 552078 49020
rect 142614 47812 142620 47864
rect 142672 47852 142678 47864
rect 215294 47852 215300 47864
rect 142672 47824 215300 47852
rect 142672 47812 142678 47824
rect 215294 47812 215300 47824
rect 215352 47812 215358 47864
rect 158990 47744 158996 47796
rect 159048 47784 159054 47796
rect 436094 47784 436100 47796
rect 159048 47756 436100 47784
rect 159048 47744 159054 47756
rect 436094 47744 436100 47756
rect 436152 47744 436158 47796
rect 160554 47676 160560 47728
rect 160612 47716 160618 47728
rect 451274 47716 451280 47728
rect 160612 47688 451280 47716
rect 160612 47676 160618 47688
rect 451274 47676 451280 47688
rect 451332 47676 451338 47728
rect 163222 47608 163228 47660
rect 163280 47648 163286 47660
rect 484394 47648 484400 47660
rect 163280 47620 484400 47648
rect 163280 47608 163286 47620
rect 484394 47608 484400 47620
rect 484452 47608 484458 47660
rect 45554 47540 45560 47592
rect 45612 47580 45618 47592
rect 120902 47580 120908 47592
rect 45612 47552 120908 47580
rect 45612 47540 45618 47552
rect 120902 47540 120908 47552
rect 120960 47540 120966 47592
rect 138382 47540 138388 47592
rect 138440 47580 138446 47592
rect 153838 47580 153844 47592
rect 138440 47552 153844 47580
rect 138440 47540 138446 47552
rect 153838 47540 153844 47552
rect 153896 47540 153902 47592
rect 170030 47540 170036 47592
rect 170088 47580 170094 47592
rect 571334 47580 571340 47592
rect 170088 47552 571340 47580
rect 170088 47540 170094 47552
rect 571334 47540 571340 47552
rect 571392 47540 571398 47592
rect 118418 46860 118424 46912
rect 118476 46900 118482 46912
rect 580166 46900 580172 46912
rect 118476 46872 580172 46900
rect 118476 46860 118482 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 137002 46792 137008 46844
rect 137060 46832 137066 46844
rect 138658 46832 138664 46844
rect 137060 46804 138664 46832
rect 137060 46792 137066 46804
rect 138658 46792 138664 46804
rect 138716 46792 138722 46844
rect 141050 46384 141056 46436
rect 141108 46424 141114 46436
rect 208394 46424 208400 46436
rect 141108 46396 208400 46424
rect 141108 46384 141114 46396
rect 208394 46384 208400 46396
rect 208452 46384 208458 46436
rect 144178 46316 144184 46368
rect 144236 46356 144242 46368
rect 233234 46356 233240 46368
rect 144236 46328 233240 46356
rect 144236 46316 144242 46328
rect 233234 46316 233240 46328
rect 233292 46316 233298 46368
rect 156230 46248 156236 46300
rect 156288 46288 156294 46300
rect 391934 46288 391940 46300
rect 156288 46260 391940 46288
rect 156288 46248 156294 46260
rect 391934 46248 391940 46260
rect 391992 46248 391998 46300
rect 138290 46180 138296 46232
rect 138348 46220 138354 46232
rect 156598 46220 156604 46232
rect 138348 46192 156604 46220
rect 138348 46180 138354 46192
rect 156598 46180 156604 46192
rect 156656 46180 156662 46232
rect 163130 46180 163136 46232
rect 163188 46220 163194 46232
rect 491294 46220 491300 46232
rect 163188 46192 491300 46220
rect 163188 46180 163194 46192
rect 491294 46180 491300 46192
rect 491352 46180 491358 46232
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 173986 45540 173992 45552
rect 3568 45512 173992 45540
rect 3568 45500 3574 45512
rect 173986 45500 173992 45512
rect 174044 45500 174050 45552
rect 142522 45024 142528 45076
rect 142580 45064 142586 45076
rect 218146 45064 218152 45076
rect 142580 45036 218152 45064
rect 142580 45024 142586 45036
rect 218146 45024 218152 45036
rect 218204 45024 218210 45076
rect 148134 44956 148140 45008
rect 148192 44996 148198 45008
rect 289814 44996 289820 45008
rect 148192 44968 289820 44996
rect 148192 44956 148198 44968
rect 289814 44956 289820 44968
rect 289872 44956 289878 45008
rect 171870 44888 171876 44940
rect 171928 44928 171934 44940
rect 397454 44928 397460 44940
rect 171928 44900 397460 44928
rect 171928 44888 171934 44900
rect 397454 44888 397460 44900
rect 397512 44888 397518 44940
rect 81434 44820 81440 44872
rect 81492 44860 81498 44872
rect 131390 44860 131396 44872
rect 81492 44832 131396 44860
rect 81492 44820 81498 44832
rect 131390 44820 131396 44832
rect 131448 44820 131454 44872
rect 168742 44820 168748 44872
rect 168800 44860 168806 44872
rect 553394 44860 553400 44872
rect 168800 44832 553400 44860
rect 168800 44820 168806 44832
rect 553394 44820 553400 44832
rect 553452 44820 553458 44872
rect 148042 43528 148048 43580
rect 148100 43568 148106 43580
rect 285674 43568 285680 43580
rect 148100 43540 285680 43568
rect 148100 43528 148106 43540
rect 285674 43528 285680 43540
rect 285732 43528 285738 43580
rect 171502 43460 171508 43512
rect 171560 43500 171566 43512
rect 432046 43500 432052 43512
rect 171560 43472 432052 43500
rect 171560 43460 171566 43472
rect 432046 43460 432052 43472
rect 432104 43460 432110 43512
rect 88334 43392 88340 43444
rect 88392 43432 88398 43444
rect 125226 43432 125232 43444
rect 88392 43404 125232 43432
rect 88392 43392 88398 43404
rect 125226 43392 125232 43404
rect 125284 43392 125290 43444
rect 169662 43392 169668 43444
rect 169720 43432 169726 43444
rect 563054 43432 563060 43444
rect 169720 43404 563060 43432
rect 169720 43392 169726 43404
rect 563054 43392 563060 43404
rect 563112 43392 563118 43444
rect 139486 42168 139492 42220
rect 139544 42208 139550 42220
rect 187694 42208 187700 42220
rect 139544 42180 187700 42208
rect 139544 42168 139550 42180
rect 187694 42168 187700 42180
rect 187752 42168 187758 42220
rect 157702 42100 157708 42152
rect 157760 42140 157766 42152
rect 415486 42140 415492 42152
rect 157760 42112 415492 42140
rect 157760 42100 157766 42112
rect 415486 42100 415492 42112
rect 415544 42100 415550 42152
rect 169938 42032 169944 42084
rect 169996 42072 170002 42084
rect 572806 42072 572812 42084
rect 169996 42044 572812 42072
rect 169996 42032 170002 42044
rect 572806 42032 572812 42044
rect 572864 42032 572870 42084
rect 152274 40740 152280 40792
rect 152332 40780 152338 40792
rect 345014 40780 345020 40792
rect 152332 40752 345020 40780
rect 152332 40740 152338 40752
rect 345014 40740 345020 40752
rect 345072 40740 345078 40792
rect 169846 40672 169852 40724
rect 169904 40712 169910 40724
rect 569954 40712 569960 40724
rect 169904 40684 569960 40712
rect 169904 40672 169910 40684
rect 569954 40672 569960 40684
rect 570012 40672 570018 40724
rect 153378 39448 153384 39500
rect 153436 39488 153442 39500
rect 357526 39488 357532 39500
rect 153436 39460 357532 39488
rect 153436 39448 153442 39460
rect 357526 39448 357532 39460
rect 357584 39448 357590 39500
rect 157610 39380 157616 39432
rect 157668 39420 157674 39432
rect 409874 39420 409880 39432
rect 157668 39392 409880 39420
rect 157668 39380 157674 39392
rect 409874 39380 409880 39392
rect 409932 39380 409938 39432
rect 166074 39312 166080 39364
rect 166132 39352 166138 39364
rect 527174 39352 527180 39364
rect 166132 39324 527180 39352
rect 166132 39312 166138 39324
rect 527174 39312 527180 39324
rect 527232 39312 527238 39364
rect 157518 37952 157524 38004
rect 157576 37992 157582 38004
rect 419534 37992 419540 38004
rect 157576 37964 419540 37992
rect 157576 37952 157582 37964
rect 419534 37952 419540 37964
rect 419592 37952 419598 38004
rect 164602 37884 164608 37936
rect 164660 37924 164666 37936
rect 503714 37924 503720 37936
rect 164660 37896 503720 37924
rect 164660 37884 164666 37896
rect 503714 37884 503720 37896
rect 503772 37884 503778 37936
rect 31754 36524 31760 36576
rect 31812 36564 31818 36576
rect 122374 36564 122380 36576
rect 31812 36536 122380 36564
rect 31812 36524 31818 36536
rect 122374 36524 122380 36536
rect 122432 36524 122438 36576
rect 27614 35164 27620 35216
rect 27672 35204 27678 35216
rect 127250 35204 127256 35216
rect 27672 35176 127256 35204
rect 27672 35164 27678 35176
rect 127250 35164 127256 35176
rect 127308 35164 127314 35216
rect 163038 35164 163044 35216
rect 163096 35204 163102 35216
rect 487154 35204 487160 35216
rect 163096 35176 487160 35204
rect 163096 35164 163102 35176
rect 487154 35164 487160 35176
rect 487212 35164 487218 35216
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 21450 33096 21456 33108
rect 2924 33068 21456 33096
rect 2924 33056 2930 33068
rect 21450 33056 21456 33068
rect 21508 33056 21514 33108
rect 147858 32444 147864 32496
rect 147916 32484 147922 32496
rect 291194 32484 291200 32496
rect 147916 32456 291200 32484
rect 147916 32444 147922 32456
rect 291194 32444 291200 32456
rect 291252 32444 291258 32496
rect 147950 32376 147956 32428
rect 148008 32416 148014 32428
rect 293954 32416 293960 32428
rect 148008 32388 293960 32416
rect 148008 32376 148014 32388
rect 293954 32376 293960 32388
rect 294012 32376 294018 32428
rect 140958 31356 140964 31408
rect 141016 31396 141022 31408
rect 205634 31396 205640 31408
rect 141016 31368 205640 31396
rect 141016 31356 141022 31368
rect 205634 31356 205640 31368
rect 205692 31356 205698 31408
rect 142430 31288 142436 31340
rect 142488 31328 142494 31340
rect 216674 31328 216680 31340
rect 142488 31300 216680 31328
rect 142488 31288 142494 31300
rect 216674 31288 216680 31300
rect 216732 31288 216738 31340
rect 144086 31220 144092 31272
rect 144144 31260 144150 31272
rect 237374 31260 237380 31272
rect 144144 31232 237380 31260
rect 144144 31220 144150 31232
rect 237374 31220 237380 31232
rect 237432 31220 237438 31272
rect 164510 31152 164516 31204
rect 164568 31192 164574 31204
rect 499574 31192 499580 31204
rect 164568 31164 499580 31192
rect 164568 31152 164574 31164
rect 499574 31152 499580 31164
rect 499632 31152 499638 31204
rect 167362 31084 167368 31136
rect 167420 31124 167426 31136
rect 535454 31124 535460 31136
rect 167420 31096 535460 31124
rect 167420 31084 167426 31096
rect 535454 31084 535460 31096
rect 535512 31084 535518 31136
rect 169754 31016 169760 31068
rect 169812 31056 169818 31068
rect 574094 31056 574100 31068
rect 169812 31028 574100 31056
rect 169812 31016 169818 31028
rect 574094 31016 574100 31028
rect 574152 31016 574158 31068
rect 150710 29792 150716 29844
rect 150768 29832 150774 29844
rect 324406 29832 324412 29844
rect 150768 29804 324412 29832
rect 150768 29792 150774 29804
rect 324406 29792 324412 29804
rect 324464 29792 324470 29844
rect 152182 29724 152188 29776
rect 152240 29764 152246 29776
rect 339494 29764 339500 29776
rect 152240 29736 339500 29764
rect 152240 29724 152246 29736
rect 339494 29724 339500 29736
rect 339552 29724 339558 29776
rect 153102 29656 153108 29708
rect 153160 29696 153166 29708
rect 346394 29696 346400 29708
rect 153160 29668 346400 29696
rect 153160 29656 153166 29668
rect 346394 29656 346400 29668
rect 346452 29656 346458 29708
rect 158898 29588 158904 29640
rect 158956 29628 158962 29640
rect 427814 29628 427820 29640
rect 158956 29600 427820 29628
rect 158956 29588 158962 29600
rect 427814 29588 427820 29600
rect 427872 29588 427878 29640
rect 150618 28364 150624 28416
rect 150676 28404 150682 28416
rect 321554 28404 321560 28416
rect 150676 28376 321560 28404
rect 150676 28364 150682 28376
rect 321554 28364 321560 28376
rect 321612 28364 321618 28416
rect 153286 28296 153292 28348
rect 153344 28336 153350 28348
rect 360194 28336 360200 28348
rect 153344 28308 360200 28336
rect 153344 28296 153350 28308
rect 360194 28296 360200 28308
rect 360252 28296 360258 28348
rect 172146 28228 172152 28280
rect 172204 28268 172210 28280
rect 418154 28268 418160 28280
rect 172204 28240 418160 28268
rect 172204 28228 172210 28240
rect 418154 28228 418160 28240
rect 418212 28228 418218 28280
rect 145282 26936 145288 26988
rect 145340 26976 145346 26988
rect 258074 26976 258080 26988
rect 145340 26948 258080 26976
rect 145340 26936 145346 26948
rect 258074 26936 258080 26948
rect 258132 26936 258138 26988
rect 154758 26868 154764 26920
rect 154816 26908 154822 26920
rect 378134 26908 378140 26920
rect 154816 26880 378140 26908
rect 154816 26868 154822 26880
rect 378134 26868 378140 26880
rect 378192 26868 378198 26920
rect 143994 25644 144000 25696
rect 144052 25684 144058 25696
rect 235994 25684 236000 25696
rect 144052 25656 236000 25684
rect 144052 25644 144058 25656
rect 235994 25644 236000 25656
rect 236052 25644 236058 25696
rect 145190 25576 145196 25628
rect 145248 25616 145254 25628
rect 251266 25616 251272 25628
rect 145248 25588 251272 25616
rect 145248 25576 145254 25588
rect 251266 25576 251272 25588
rect 251324 25576 251330 25628
rect 154666 25508 154672 25560
rect 154724 25548 154730 25560
rect 385034 25548 385040 25560
rect 154724 25520 385040 25548
rect 154724 25508 154730 25520
rect 385034 25508 385040 25520
rect 385092 25508 385098 25560
rect 142338 24216 142344 24268
rect 142396 24256 142402 24268
rect 222194 24256 222200 24268
rect 142396 24228 222200 24256
rect 142396 24216 142402 24228
rect 222194 24216 222200 24228
rect 222252 24216 222258 24268
rect 147766 24148 147772 24200
rect 147824 24188 147830 24200
rect 292666 24188 292672 24200
rect 147824 24160 292672 24188
rect 147824 24148 147830 24160
rect 292666 24148 292672 24160
rect 292724 24148 292730 24200
rect 106274 24080 106280 24132
rect 106332 24120 106338 24132
rect 132862 24120 132868 24132
rect 106332 24092 132868 24120
rect 106332 24080 106338 24092
rect 132862 24080 132868 24092
rect 132920 24080 132926 24132
rect 165982 24080 165988 24132
rect 166040 24120 166046 24132
rect 524414 24120 524420 24132
rect 166040 24092 524420 24120
rect 166040 24080 166046 24092
rect 524414 24080 524420 24092
rect 524472 24080 524478 24132
rect 139394 22992 139400 23044
rect 139452 23032 139458 23044
rect 186314 23032 186320 23044
rect 139452 23004 186320 23032
rect 139452 22992 139458 23004
rect 186314 22992 186320 23004
rect 186372 22992 186378 23044
rect 150526 22924 150532 22976
rect 150584 22964 150590 22976
rect 328454 22964 328460 22976
rect 150584 22936 328460 22964
rect 150584 22924 150590 22936
rect 328454 22924 328460 22936
rect 328512 22924 328518 22976
rect 67634 22856 67640 22908
rect 67692 22896 67698 22908
rect 130102 22896 130108 22908
rect 67692 22868 130108 22896
rect 67692 22856 67698 22868
rect 130102 22856 130108 22868
rect 130160 22856 130166 22908
rect 157426 22856 157432 22908
rect 157484 22896 157490 22908
rect 416774 22896 416780 22908
rect 157484 22868 416780 22896
rect 157484 22856 157490 22868
rect 416774 22856 416780 22868
rect 416832 22856 416838 22908
rect 60826 22788 60832 22840
rect 60884 22828 60890 22840
rect 129182 22828 129188 22840
rect 60884 22800 129188 22828
rect 60884 22788 60890 22800
rect 129182 22788 129188 22800
rect 129240 22788 129246 22840
rect 165890 22788 165896 22840
rect 165948 22828 165954 22840
rect 521654 22828 521660 22840
rect 165948 22800 521660 22828
rect 165948 22788 165954 22800
rect 521654 22788 521660 22800
rect 521712 22788 521718 22840
rect 3510 22720 3516 22772
rect 3568 22760 3574 22772
rect 179690 22760 179696 22772
rect 3568 22732 179696 22760
rect 3568 22720 3574 22732
rect 179690 22720 179696 22732
rect 179748 22720 179754 22772
rect 184198 22720 184204 22772
rect 184256 22760 184262 22772
rect 580166 22760 580172 22772
rect 184256 22732 580172 22760
rect 184256 22720 184262 22732
rect 580166 22720 580172 22732
rect 580224 22720 580230 22772
rect 135714 21632 135720 21684
rect 135772 21672 135778 21684
rect 139394 21672 139400 21684
rect 135772 21644 139400 21672
rect 135772 21632 135778 21644
rect 139394 21632 139400 21644
rect 139452 21632 139458 21684
rect 138198 21564 138204 21616
rect 138256 21604 138262 21616
rect 168650 21604 168656 21616
rect 138256 21576 168656 21604
rect 138256 21564 138262 21576
rect 168650 21564 168656 21576
rect 168708 21564 168714 21616
rect 154574 21496 154580 21548
rect 154632 21536 154638 21548
rect 379514 21536 379520 21548
rect 154632 21508 379520 21536
rect 154632 21496 154638 21508
rect 379514 21496 379520 21508
rect 379572 21496 379578 21548
rect 136910 21428 136916 21480
rect 136968 21468 136974 21480
rect 147766 21468 147772 21480
rect 136968 21440 147772 21468
rect 136968 21428 136974 21440
rect 147766 21428 147772 21440
rect 147824 21428 147830 21480
rect 172054 21428 172060 21480
rect 172112 21468 172118 21480
rect 404354 21468 404360 21480
rect 172112 21440 404360 21468
rect 172112 21428 172118 21440
rect 404354 21428 404360 21440
rect 404412 21428 404418 21480
rect 38654 21360 38660 21412
rect 38712 21400 38718 21412
rect 120810 21400 120816 21412
rect 38712 21372 120816 21400
rect 38712 21360 38718 21372
rect 120810 21360 120816 21372
rect 120868 21360 120874 21412
rect 168558 21360 168564 21412
rect 168616 21400 168622 21412
rect 556154 21400 556160 21412
rect 168616 21372 556160 21400
rect 168616 21360 168622 21372
rect 556154 21360 556160 21372
rect 556212 21360 556218 21412
rect 143902 20204 143908 20256
rect 143960 20244 143966 20256
rect 241514 20244 241520 20256
rect 143960 20216 241520 20244
rect 143960 20204 143966 20216
rect 241514 20204 241520 20216
rect 241572 20204 241578 20256
rect 145098 20136 145104 20188
rect 145156 20176 145162 20188
rect 262214 20176 262220 20188
rect 145156 20148 262220 20176
rect 145156 20136 145162 20148
rect 262214 20136 262220 20148
rect 262272 20136 262278 20188
rect 151998 20068 152004 20120
rect 152056 20108 152062 20120
rect 343634 20108 343640 20120
rect 152056 20080 343640 20108
rect 152056 20068 152062 20080
rect 343634 20068 343640 20080
rect 343692 20068 343698 20120
rect 124214 20000 124220 20052
rect 124272 20040 124278 20052
rect 134058 20040 134064 20052
rect 124272 20012 134064 20040
rect 124272 20000 124278 20012
rect 134058 20000 134064 20012
rect 134116 20000 134122 20052
rect 145006 20000 145012 20052
rect 145064 20040 145070 20052
rect 255314 20040 255320 20052
rect 145064 20012 255320 20040
rect 145064 20000 145070 20012
rect 255314 20000 255320 20012
rect 255372 20000 255378 20052
rect 255958 20000 255964 20052
rect 256016 20040 256022 20052
rect 456794 20040 456800 20052
rect 256016 20012 456800 20040
rect 256016 20000 256022 20012
rect 456794 20000 456800 20012
rect 456852 20000 456858 20052
rect 99374 19932 99380 19984
rect 99432 19972 99438 19984
rect 132770 19972 132776 19984
rect 99432 19944 132776 19972
rect 99432 19932 99438 19944
rect 132770 19932 132776 19944
rect 132828 19932 132834 19984
rect 156138 19932 156144 19984
rect 156196 19972 156202 19984
rect 400214 19972 400220 19984
rect 156196 19944 400220 19972
rect 156196 19932 156202 19944
rect 400214 19932 400220 19944
rect 400272 19932 400278 19984
rect 140866 18776 140872 18828
rect 140924 18816 140930 18828
rect 198734 18816 198740 18828
rect 140924 18788 198740 18816
rect 140924 18776 140930 18788
rect 198734 18776 198740 18788
rect 198792 18776 198798 18828
rect 158806 18708 158812 18760
rect 158864 18748 158870 18760
rect 429194 18748 429200 18760
rect 158864 18720 429200 18748
rect 158864 18708 158870 18720
rect 429194 18708 429200 18720
rect 429252 18708 429258 18760
rect 168374 18640 168380 18692
rect 168432 18680 168438 18692
rect 556246 18680 556252 18692
rect 168432 18652 556252 18680
rect 168432 18640 168438 18652
rect 556246 18640 556252 18652
rect 556304 18640 556310 18692
rect 168466 18572 168472 18624
rect 168524 18612 168530 18624
rect 560294 18612 560300 18624
rect 168524 18584 560300 18612
rect 168524 18572 168530 18584
rect 560294 18572 560300 18584
rect 560352 18572 560358 18624
rect 160462 17416 160468 17468
rect 160520 17456 160526 17468
rect 445754 17456 445760 17468
rect 160520 17428 445760 17456
rect 160520 17416 160526 17428
rect 445754 17416 445760 17428
rect 445812 17416 445818 17468
rect 160370 17348 160376 17400
rect 160428 17388 160434 17400
rect 452654 17388 452660 17400
rect 160428 17360 452660 17388
rect 160428 17348 160434 17360
rect 452654 17348 452660 17360
rect 452712 17348 452718 17400
rect 162946 17280 162952 17332
rect 163004 17320 163010 17332
rect 492674 17320 492680 17332
rect 163004 17292 492680 17320
rect 163004 17280 163010 17292
rect 492674 17280 492680 17292
rect 492732 17280 492738 17332
rect 167270 17212 167276 17264
rect 167328 17252 167334 17264
rect 540974 17252 540980 17264
rect 167328 17224 540980 17252
rect 167328 17212 167334 17224
rect 540974 17212 540980 17224
rect 541032 17212 541038 17264
rect 151906 16124 151912 16176
rect 151964 16164 151970 16176
rect 342898 16164 342904 16176
rect 151964 16136 342904 16164
rect 151964 16124 151970 16136
rect 342898 16124 342904 16136
rect 342956 16124 342962 16176
rect 160186 16056 160192 16108
rect 160244 16096 160250 16108
rect 448606 16096 448612 16108
rect 160244 16068 448612 16096
rect 160244 16056 160250 16068
rect 448606 16056 448612 16068
rect 448664 16056 448670 16108
rect 160278 15988 160284 16040
rect 160336 16028 160342 16040
rect 454034 16028 454040 16040
rect 160336 16000 454040 16028
rect 160336 15988 160342 16000
rect 454034 15988 454040 16000
rect 454092 15988 454098 16040
rect 165706 15920 165712 15972
rect 165764 15960 165770 15972
rect 517882 15960 517888 15972
rect 165764 15932 517888 15960
rect 165764 15920 165770 15932
rect 517882 15920 517888 15932
rect 517940 15920 517946 15972
rect 165798 15852 165804 15904
rect 165856 15892 165862 15904
rect 523770 15892 523776 15904
rect 165856 15864 523776 15892
rect 165856 15852 165862 15864
rect 523770 15852 523776 15864
rect 523828 15852 523834 15904
rect 144914 14764 144920 14816
rect 144972 14804 144978 14816
rect 254210 14804 254216 14816
rect 144972 14776 254216 14804
rect 144972 14764 144978 14776
rect 254210 14764 254216 14776
rect 254268 14764 254274 14816
rect 149790 14696 149796 14748
rect 149848 14736 149854 14748
rect 305546 14736 305552 14748
rect 149848 14708 305552 14736
rect 149848 14696 149854 14708
rect 305546 14696 305552 14708
rect 305604 14696 305610 14748
rect 149698 14628 149704 14680
rect 149756 14668 149762 14680
rect 307754 14668 307760 14680
rect 149756 14640 307760 14668
rect 149756 14628 149762 14640
rect 307754 14628 307760 14640
rect 307812 14628 307818 14680
rect 124122 14560 124128 14612
rect 124180 14600 124186 14612
rect 312170 14600 312176 14612
rect 124180 14572 312176 14600
rect 124180 14560 124186 14572
rect 312170 14560 312176 14572
rect 312228 14560 312234 14612
rect 315298 14560 315304 14612
rect 315356 14600 315362 14612
rect 475746 14600 475752 14612
rect 315356 14572 475752 14600
rect 315356 14560 315362 14572
rect 475746 14560 475752 14572
rect 475804 14560 475810 14612
rect 156046 14492 156052 14544
rect 156104 14532 156110 14544
rect 398926 14532 398932 14544
rect 156104 14504 398932 14532
rect 156104 14492 156110 14504
rect 398926 14492 398932 14504
rect 398984 14492 398990 14544
rect 165614 14424 165620 14476
rect 165672 14464 165678 14476
rect 520274 14464 520280 14476
rect 165672 14436 520280 14464
rect 165672 14424 165678 14436
rect 520274 14424 520280 14436
rect 520332 14424 520338 14476
rect 15930 13064 15936 13116
rect 15988 13104 15994 13116
rect 113818 13104 113824 13116
rect 15988 13076 113824 13104
rect 15988 13064 15994 13076
rect 113818 13064 113824 13076
rect 113876 13064 113882 13116
rect 140774 12316 140780 12368
rect 140832 12356 140838 12368
rect 202690 12356 202696 12368
rect 140832 12328 202696 12356
rect 140832 12316 140838 12328
rect 202690 12316 202696 12328
rect 202748 12316 202754 12368
rect 147030 12248 147036 12300
rect 147088 12288 147094 12300
rect 273254 12288 273260 12300
rect 147088 12260 273260 12288
rect 147088 12248 147094 12260
rect 273254 12248 273260 12260
rect 273312 12248 273318 12300
rect 146938 12180 146944 12232
rect 146996 12220 147002 12232
rect 276658 12220 276664 12232
rect 146996 12192 276664 12220
rect 146996 12180 147002 12192
rect 276658 12180 276664 12192
rect 276716 12180 276722 12232
rect 147674 12112 147680 12164
rect 147732 12152 147738 12164
rect 287330 12152 287336 12164
rect 147732 12124 287336 12152
rect 147732 12112 147738 12124
rect 287330 12112 287336 12124
rect 287388 12112 287394 12164
rect 149514 12044 149520 12096
rect 149572 12084 149578 12096
rect 311434 12084 311440 12096
rect 149572 12056 311440 12084
rect 149572 12044 149578 12056
rect 311434 12044 311440 12056
rect 311492 12044 311498 12096
rect 149606 11976 149612 12028
rect 149664 12016 149670 12028
rect 314654 12016 314660 12028
rect 149664 11988 314660 12016
rect 149664 11976 149670 11988
rect 314654 11976 314660 11988
rect 314712 11976 314718 12028
rect 160002 11908 160008 11960
rect 160060 11948 160066 11960
rect 435082 11948 435088 11960
rect 160060 11920 435088 11948
rect 160060 11908 160066 11920
rect 435082 11908 435088 11920
rect 435140 11908 435146 11960
rect 160094 11840 160100 11892
rect 160152 11880 160158 11892
rect 447410 11880 447416 11892
rect 160152 11852 447416 11880
rect 160152 11840 160158 11852
rect 447410 11840 447416 11852
rect 447468 11840 447474 11892
rect 140406 11772 140412 11824
rect 140464 11812 140470 11824
rect 156138 11812 156144 11824
rect 140464 11784 156144 11812
rect 140464 11772 140470 11784
rect 156138 11772 156144 11784
rect 156196 11772 156202 11824
rect 162026 11772 162032 11824
rect 162084 11812 162090 11824
rect 463970 11812 463976 11824
rect 162084 11784 463976 11812
rect 162084 11772 162090 11784
rect 463970 11772 463976 11784
rect 464028 11772 464034 11824
rect 136818 11704 136824 11756
rect 136876 11744 136882 11756
rect 153746 11744 153752 11756
rect 136876 11716 153752 11744
rect 136876 11704 136882 11716
rect 153746 11704 153752 11716
rect 153804 11704 153810 11756
rect 161934 11704 161940 11756
rect 161992 11744 161998 11756
rect 470594 11744 470600 11756
rect 161992 11716 470600 11744
rect 161992 11704 161998 11716
rect 470594 11704 470600 11716
rect 470652 11704 470658 11756
rect 173526 11636 173532 11688
rect 173584 11676 173590 11688
rect 173710 11676 173716 11688
rect 173584 11648 173716 11676
rect 173584 11636 173590 11648
rect 173710 11636 173716 11648
rect 173768 11636 173774 11688
rect 110506 10412 110512 10464
rect 110564 10452 110570 10464
rect 125134 10452 125140 10464
rect 110564 10424 125140 10452
rect 110564 10412 110570 10424
rect 125134 10412 125140 10424
rect 125192 10412 125198 10464
rect 25314 10344 25320 10396
rect 25372 10384 25378 10396
rect 106918 10384 106924 10396
rect 25372 10356 106924 10384
rect 25372 10344 25378 10356
rect 106918 10344 106924 10356
rect 106976 10344 106982 10396
rect 117314 10344 117320 10396
rect 117372 10384 117378 10396
rect 134426 10384 134432 10396
rect 117372 10356 134432 10384
rect 117372 10344 117378 10356
rect 134426 10344 134432 10356
rect 134484 10344 134490 10396
rect 44266 10276 44272 10328
rect 44324 10316 44330 10328
rect 128538 10316 128544 10328
rect 44324 10288 128544 10316
rect 44324 10276 44330 10288
rect 128538 10276 128544 10288
rect 128596 10276 128602 10328
rect 138106 10276 138112 10328
rect 138164 10316 138170 10328
rect 166074 10316 166080 10328
rect 138164 10288 166080 10316
rect 138164 10276 138170 10288
rect 166074 10276 166080 10288
rect 166132 10276 166138 10328
rect 146846 9596 146852 9648
rect 146904 9636 146910 9648
rect 272426 9636 272432 9648
rect 146904 9608 272432 9636
rect 146904 9596 146910 9608
rect 272426 9596 272432 9608
rect 272484 9596 272490 9648
rect 146662 9528 146668 9580
rect 146720 9568 146726 9580
rect 276014 9568 276020 9580
rect 146720 9540 276020 9568
rect 146720 9528 146726 9540
rect 276014 9528 276020 9540
rect 276072 9528 276078 9580
rect 149422 9460 149428 9512
rect 149480 9500 149486 9512
rect 304350 9500 304356 9512
rect 149480 9472 304356 9500
rect 149480 9460 149486 9472
rect 304350 9460 304356 9472
rect 304408 9460 304414 9512
rect 149330 9392 149336 9444
rect 149388 9432 149394 9444
rect 307938 9432 307944 9444
rect 149388 9404 307944 9432
rect 149388 9392 149394 9404
rect 307938 9392 307944 9404
rect 307996 9392 308002 9444
rect 171410 9324 171416 9376
rect 171468 9364 171474 9376
rect 411898 9364 411904 9376
rect 171468 9336 411904 9364
rect 171468 9324 171474 9336
rect 411898 9324 411904 9336
rect 411956 9324 411962 9376
rect 157334 9256 157340 9308
rect 157392 9296 157398 9308
rect 414290 9296 414296 9308
rect 157392 9268 414296 9296
rect 157392 9256 157398 9268
rect 414290 9256 414296 9268
rect 414348 9256 414354 9308
rect 161658 9188 161664 9240
rect 161716 9228 161722 9240
rect 466270 9228 466276 9240
rect 161716 9200 466276 9228
rect 161716 9188 161722 9200
rect 466270 9188 466276 9200
rect 466328 9188 466334 9240
rect 161750 9120 161756 9172
rect 161808 9160 161814 9172
rect 469858 9160 469864 9172
rect 161808 9132 469864 9160
rect 161808 9120 161814 9132
rect 469858 9120 469864 9132
rect 469916 9120 469922 9172
rect 34790 9052 34796 9104
rect 34848 9092 34854 9104
rect 127802 9092 127808 9104
rect 34848 9064 127808 9092
rect 34848 9052 34854 9064
rect 127802 9052 127808 9064
rect 127860 9052 127866 9104
rect 161842 9052 161848 9104
rect 161900 9092 161906 9104
rect 473446 9092 473452 9104
rect 161900 9064 473452 9092
rect 161900 9052 161906 9064
rect 473446 9052 473452 9064
rect 473504 9052 473510 9104
rect 24210 8984 24216 9036
rect 24268 9024 24274 9036
rect 122282 9024 122288 9036
rect 24268 8996 122288 9024
rect 24268 8984 24274 8996
rect 122282 8984 122288 8996
rect 122340 8984 122346 9036
rect 164418 8984 164424 9036
rect 164476 9024 164482 9036
rect 510062 9024 510068 9036
rect 164476 8996 510068 9024
rect 164476 8984 164482 8996
rect 510062 8984 510068 8996
rect 510120 8984 510126 9036
rect 9950 8916 9956 8968
rect 10008 8956 10014 8968
rect 125962 8956 125968 8968
rect 10008 8928 125968 8956
rect 10008 8916 10014 8928
rect 125962 8916 125968 8928
rect 126020 8916 126026 8968
rect 167178 8916 167184 8968
rect 167236 8956 167242 8968
rect 539594 8956 539600 8968
rect 167236 8928 539600 8956
rect 167236 8916 167242 8928
rect 539594 8916 539600 8928
rect 539652 8916 539658 8968
rect 146754 8848 146760 8900
rect 146812 8888 146818 8900
rect 268838 8888 268844 8900
rect 146812 8860 268844 8888
rect 146812 8848 146818 8860
rect 268838 8848 268844 8860
rect 268896 8848 268902 8900
rect 105722 7828 105728 7880
rect 105780 7868 105786 7880
rect 132954 7868 132960 7880
rect 105780 7840 132960 7868
rect 105780 7828 105786 7840
rect 132954 7828 132960 7840
rect 133012 7828 133018 7880
rect 98638 7760 98644 7812
rect 98696 7800 98702 7812
rect 133138 7800 133144 7812
rect 98696 7772 133144 7800
rect 98696 7760 98702 7772
rect 133138 7760 133144 7772
rect 133196 7760 133202 7812
rect 27706 7692 27712 7744
rect 27764 7732 27770 7744
rect 127342 7732 127348 7744
rect 27764 7704 127348 7732
rect 27764 7692 27770 7704
rect 127342 7692 127348 7704
rect 127400 7692 127406 7744
rect 23014 7624 23020 7676
rect 23072 7664 23078 7676
rect 127526 7664 127532 7676
rect 23072 7636 127532 7664
rect 23072 7624 23078 7636
rect 127526 7624 127532 7636
rect 127584 7624 127590 7676
rect 150434 7624 150440 7676
rect 150492 7664 150498 7676
rect 330386 7664 330392 7676
rect 150492 7636 330392 7664
rect 150492 7624 150498 7636
rect 330386 7624 330392 7636
rect 330444 7624 330450 7676
rect 18230 7556 18236 7608
rect 18288 7596 18294 7608
rect 125870 7596 125876 7608
rect 18288 7568 125876 7596
rect 18288 7556 18294 7568
rect 125870 7556 125876 7568
rect 125928 7556 125934 7608
rect 164326 7556 164332 7608
rect 164384 7596 164390 7608
rect 506474 7596 506480 7608
rect 164384 7568 506480 7596
rect 164384 7556 164390 7568
rect 506474 7556 506480 7568
rect 506532 7556 506538 7608
rect 146478 6808 146484 6860
rect 146536 6848 146542 6860
rect 278314 6848 278320 6860
rect 146536 6820 278320 6848
rect 146536 6808 146542 6820
rect 278314 6808 278320 6820
rect 278372 6808 278378 6860
rect 149238 6740 149244 6792
rect 149296 6780 149302 6792
rect 310238 6780 310244 6792
rect 149296 6752 310244 6780
rect 149296 6740 149302 6752
rect 310238 6740 310244 6752
rect 310296 6740 310302 6792
rect 149146 6672 149152 6724
rect 149204 6712 149210 6724
rect 313826 6712 313832 6724
rect 149204 6684 313832 6712
rect 149204 6672 149210 6684
rect 313826 6672 313832 6684
rect 313884 6672 313890 6724
rect 172330 6604 172336 6656
rect 172388 6644 172394 6656
rect 342162 6644 342168 6656
rect 172388 6616 342168 6644
rect 172388 6604 172394 6616
rect 342162 6604 342168 6616
rect 342220 6604 342226 6656
rect 151814 6536 151820 6588
rect 151872 6576 151878 6588
rect 338666 6576 338672 6588
rect 151872 6548 338672 6576
rect 151872 6536 151878 6548
rect 338666 6536 338672 6548
rect 338724 6536 338730 6588
rect 84470 6468 84476 6520
rect 84528 6508 84534 6520
rect 131298 6508 131304 6520
rect 84528 6480 131304 6508
rect 84528 6468 84534 6480
rect 131298 6468 131304 6480
rect 131356 6468 131362 6520
rect 153194 6468 153200 6520
rect 153252 6508 153258 6520
rect 364610 6508 364616 6520
rect 153252 6480 364616 6508
rect 153252 6468 153258 6480
rect 364610 6468 364616 6480
rect 364668 6468 364674 6520
rect 80882 6400 80888 6452
rect 80940 6440 80946 6452
rect 131666 6440 131672 6452
rect 80940 6412 131672 6440
rect 80940 6400 80946 6412
rect 131666 6400 131672 6412
rect 131724 6400 131730 6452
rect 155954 6400 155960 6452
rect 156012 6440 156018 6452
rect 394234 6440 394240 6452
rect 156012 6412 394240 6440
rect 156012 6400 156018 6412
rect 394234 6400 394240 6412
rect 394292 6400 394298 6452
rect 78582 6332 78588 6384
rect 78640 6372 78646 6384
rect 128998 6372 129004 6384
rect 78640 6344 129004 6372
rect 78640 6332 78646 6344
rect 128998 6332 129004 6344
rect 129056 6332 129062 6384
rect 161566 6332 161572 6384
rect 161624 6372 161630 6384
rect 462774 6372 462780 6384
rect 161624 6344 462780 6372
rect 161624 6332 161630 6344
rect 462774 6332 462780 6344
rect 462832 6332 462838 6384
rect 70302 6264 70308 6316
rect 70360 6304 70366 6316
rect 130010 6304 130016 6316
rect 70360 6276 130016 6304
rect 70360 6264 70366 6276
rect 130010 6264 130016 6276
rect 130068 6264 130074 6316
rect 161474 6264 161480 6316
rect 161532 6304 161538 6316
rect 467466 6304 467472 6316
rect 161532 6276 467472 6304
rect 161532 6264 161538 6276
rect 467466 6264 467472 6276
rect 467524 6264 467530 6316
rect 63218 6196 63224 6248
rect 63276 6236 63282 6248
rect 130470 6236 130476 6248
rect 63276 6208 130476 6236
rect 63276 6196 63282 6208
rect 130470 6196 130476 6208
rect 130528 6196 130534 6248
rect 164234 6196 164240 6248
rect 164292 6236 164298 6248
rect 502978 6236 502984 6248
rect 164292 6208 502984 6236
rect 164292 6196 164298 6208
rect 502978 6196 502984 6208
rect 503036 6196 503042 6248
rect 538858 6196 538864 6248
rect 538916 6236 538922 6248
rect 580994 6236 581000 6248
rect 538916 6208 581000 6236
rect 538916 6196 538922 6208
rect 580994 6196 581000 6208
rect 581052 6196 581058 6248
rect 13538 6128 13544 6180
rect 13596 6168 13602 6180
rect 126514 6168 126520 6180
rect 13596 6140 126520 6168
rect 13596 6128 13602 6140
rect 126514 6128 126520 6140
rect 126572 6128 126578 6180
rect 167086 6128 167092 6180
rect 167144 6168 167150 6180
rect 545482 6168 545488 6180
rect 167144 6140 545488 6168
rect 167144 6128 167150 6140
rect 545482 6128 545488 6140
rect 545540 6128 545546 6180
rect 146570 6060 146576 6112
rect 146628 6100 146634 6112
rect 274818 6100 274824 6112
rect 146628 6072 274824 6100
rect 146628 6060 146634 6072
rect 274818 6060 274824 6072
rect 274876 6060 274882 6112
rect 146386 5992 146392 6044
rect 146444 6032 146450 6044
rect 270034 6032 270040 6044
rect 146444 6004 270040 6032
rect 146444 5992 146450 6004
rect 270034 5992 270040 6004
rect 270092 5992 270098 6044
rect 85666 5108 85672 5160
rect 85724 5148 85730 5160
rect 131574 5148 131580 5160
rect 85724 5120 131580 5148
rect 85724 5108 85730 5120
rect 131574 5108 131580 5120
rect 131632 5108 131638 5160
rect 66714 5040 66720 5092
rect 66772 5080 66778 5092
rect 130286 5080 130292 5092
rect 66772 5052 130292 5080
rect 66772 5040 66778 5052
rect 130286 5040 130292 5052
rect 130344 5040 130350 5092
rect 52546 4972 52552 5024
rect 52604 5012 52610 5024
rect 128722 5012 128728 5024
rect 52604 4984 128728 5012
rect 52604 4972 52610 4984
rect 128722 4972 128728 4984
rect 128780 4972 128786 5024
rect 138014 4972 138020 5024
rect 138072 5012 138078 5024
rect 167178 5012 167184 5024
rect 138072 4984 167184 5012
rect 138072 4972 138078 4984
rect 167178 4972 167184 4984
rect 167236 4972 167242 5024
rect 6454 4904 6460 4956
rect 6512 4944 6518 4956
rect 17218 4944 17224 4956
rect 6512 4916 17224 4944
rect 6512 4904 6518 4916
rect 17218 4904 17224 4916
rect 17276 4904 17282 4956
rect 48958 4904 48964 4956
rect 49016 4944 49022 4956
rect 128906 4944 128912 4956
rect 49016 4916 128912 4944
rect 49016 4904 49022 4916
rect 128906 4904 128912 4916
rect 128964 4904 128970 4956
rect 143810 4904 143816 4956
rect 143868 4944 143874 4956
rect 234614 4944 234620 4956
rect 143868 4916 234620 4944
rect 143868 4904 143874 4916
rect 234614 4904 234620 4916
rect 234672 4904 234678 4956
rect 8754 4836 8760 4888
rect 8812 4876 8818 4888
rect 126330 4876 126336 4888
rect 8812 4848 126336 4876
rect 8812 4836 8818 4848
rect 126330 4836 126336 4848
rect 126388 4836 126394 4888
rect 137922 4836 137928 4888
rect 137980 4876 137986 4888
rect 151814 4876 151820 4888
rect 137980 4848 151820 4876
rect 137980 4836 137986 4848
rect 151814 4836 151820 4848
rect 151872 4836 151878 4888
rect 162854 4836 162860 4888
rect 162912 4876 162918 4888
rect 486418 4876 486424 4888
rect 162912 4848 486424 4876
rect 162912 4836 162918 4848
rect 486418 4836 486424 4848
rect 486476 4836 486482 4888
rect 5258 4768 5264 4820
rect 5316 4808 5322 4820
rect 126054 4808 126060 4820
rect 5316 4780 126060 4808
rect 5316 4768 5322 4780
rect 126054 4768 126060 4780
rect 126112 4768 126118 4820
rect 136726 4768 136732 4820
rect 136784 4808 136790 4820
rect 157794 4808 157800 4820
rect 136784 4780 157800 4808
rect 136784 4768 136790 4780
rect 157794 4768 157800 4780
rect 157852 4768 157858 4820
rect 168282 4768 168288 4820
rect 168340 4808 168346 4820
rect 538398 4808 538404 4820
rect 168340 4780 538404 4808
rect 168340 4768 168346 4780
rect 538398 4768 538404 4780
rect 538456 4768 538462 4820
rect 138934 4360 138940 4412
rect 138992 4400 138998 4412
rect 143534 4400 143540 4412
rect 138992 4372 143540 4400
rect 138992 4360 138998 4372
rect 143534 4360 143540 4372
rect 143592 4360 143598 4412
rect 125870 4088 125876 4140
rect 125928 4128 125934 4140
rect 134518 4128 134524 4140
rect 125928 4100 134524 4128
rect 125928 4088 125934 4100
rect 134518 4088 134524 4100
rect 134576 4088 134582 4140
rect 142246 4088 142252 4140
rect 142304 4128 142310 4140
rect 221550 4128 221556 4140
rect 142304 4100 221556 4128
rect 142304 4088 142310 4100
rect 221550 4088 221556 4100
rect 221608 4088 221614 4140
rect 143718 4020 143724 4072
rect 143776 4060 143782 4072
rect 235810 4060 235816 4072
rect 143776 4032 235816 4060
rect 143776 4020 143782 4032
rect 235810 4020 235816 4032
rect 235868 4020 235874 4072
rect 144546 3952 144552 4004
rect 144604 3992 144610 4004
rect 239306 3992 239312 4004
rect 144604 3964 239312 3992
rect 144604 3952 144610 3964
rect 239306 3952 239312 3964
rect 239364 3952 239370 4004
rect 117682 3884 117688 3936
rect 117740 3924 117746 3936
rect 122190 3924 122196 3936
rect 117740 3896 122196 3924
rect 117740 3884 117746 3896
rect 122190 3884 122196 3896
rect 122248 3884 122254 3936
rect 143626 3884 143632 3936
rect 143684 3924 143690 3936
rect 242894 3924 242900 3936
rect 143684 3896 242900 3924
rect 143684 3884 143690 3896
rect 242894 3884 242900 3896
rect 242952 3884 242958 3936
rect 251174 3884 251180 3936
rect 251232 3924 251238 3936
rect 252370 3924 252376 3936
rect 251232 3896 252376 3924
rect 251232 3884 251238 3896
rect 252370 3884 252376 3896
rect 252428 3884 252434 3936
rect 259454 3884 259460 3936
rect 259512 3924 259518 3936
rect 260650 3924 260656 3936
rect 259512 3896 260656 3924
rect 259512 3884 259518 3896
rect 260650 3884 260656 3896
rect 260708 3884 260714 3936
rect 77386 3816 77392 3868
rect 77444 3856 77450 3868
rect 123478 3856 123484 3868
rect 77444 3828 123484 3856
rect 77444 3816 77450 3828
rect 123478 3816 123484 3828
rect 123536 3816 123542 3868
rect 128170 3816 128176 3868
rect 128228 3856 128234 3868
rect 131758 3856 131764 3868
rect 128228 3828 131764 3856
rect 128228 3816 128234 3828
rect 131758 3816 131764 3828
rect 131816 3816 131822 3868
rect 140222 3816 140228 3868
rect 140280 3856 140286 3868
rect 144730 3856 144736 3868
rect 140280 3828 144736 3856
rect 140280 3816 140286 3828
rect 144730 3816 144736 3828
rect 144788 3816 144794 3868
rect 146294 3816 146300 3868
rect 146352 3856 146358 3868
rect 271230 3856 271236 3868
rect 146352 3828 271236 3856
rect 146352 3816 146358 3828
rect 271230 3816 271236 3828
rect 271288 3816 271294 3868
rect 284294 3816 284300 3868
rect 284352 3856 284358 3868
rect 285030 3856 285036 3868
rect 284352 3828 285036 3856
rect 284352 3816 284358 3828
rect 285030 3816 285036 3828
rect 285088 3816 285094 3868
rect 299566 3816 299572 3868
rect 299624 3856 299630 3868
rect 300762 3856 300768 3868
rect 299624 3828 300768 3856
rect 299624 3816 299630 3828
rect 300762 3816 300768 3828
rect 300820 3816 300826 3868
rect 64322 3748 64328 3800
rect 64380 3788 64386 3800
rect 126238 3788 126244 3800
rect 64380 3760 126244 3788
rect 64380 3748 64386 3760
rect 126238 3748 126244 3760
rect 126296 3748 126302 3800
rect 138658 3748 138664 3800
rect 138716 3788 138722 3800
rect 145926 3788 145932 3800
rect 138716 3760 145932 3788
rect 138716 3748 138722 3760
rect 145926 3748 145932 3760
rect 145984 3748 145990 3800
rect 149054 3748 149060 3800
rect 149112 3788 149118 3800
rect 306742 3788 306748 3800
rect 149112 3760 306748 3788
rect 149112 3748 149118 3760
rect 306742 3748 306748 3760
rect 306800 3748 306806 3800
rect 47854 3680 47860 3732
rect 47912 3720 47918 3732
rect 123570 3720 123576 3732
rect 47912 3692 123576 3720
rect 47912 3680 47918 3692
rect 123570 3680 123576 3692
rect 123628 3680 123634 3732
rect 131758 3680 131764 3732
rect 131816 3720 131822 3732
rect 135622 3720 135628 3732
rect 131816 3692 135628 3720
rect 131816 3680 131822 3692
rect 135622 3680 135628 3692
rect 135680 3680 135686 3732
rect 142890 3680 142896 3732
rect 142948 3720 142954 3732
rect 155402 3720 155408 3732
rect 142948 3692 155408 3720
rect 142948 3680 142954 3692
rect 155402 3680 155408 3692
rect 155460 3680 155466 3732
rect 156598 3680 156604 3732
rect 156656 3720 156662 3732
rect 168374 3720 168380 3732
rect 156656 3692 168380 3720
rect 156656 3680 156662 3692
rect 168374 3680 168380 3692
rect 168432 3680 168438 3732
rect 173526 3680 173532 3732
rect 173584 3720 173590 3732
rect 178126 3720 178132 3732
rect 173584 3692 178132 3720
rect 173584 3680 173590 3692
rect 178126 3680 178132 3692
rect 178184 3680 178190 3732
rect 184934 3680 184940 3732
rect 184992 3720 184998 3732
rect 186130 3720 186136 3732
rect 184992 3692 186136 3720
rect 184992 3680 184998 3692
rect 186130 3680 186136 3692
rect 186188 3680 186194 3732
rect 186222 3680 186228 3732
rect 186280 3720 186286 3732
rect 468662 3720 468668 3732
rect 186280 3692 468668 3720
rect 186280 3680 186286 3692
rect 468662 3680 468668 3692
rect 468720 3680 468726 3732
rect 43070 3612 43076 3664
rect 43128 3652 43134 3664
rect 125042 3652 125048 3664
rect 43128 3624 125048 3652
rect 43128 3612 43134 3624
rect 125042 3612 125048 3624
rect 125100 3612 125106 3664
rect 133782 3612 133788 3664
rect 133840 3652 133846 3664
rect 147122 3652 147128 3664
rect 133840 3624 147128 3652
rect 133840 3612 133846 3624
rect 147122 3612 147128 3624
rect 147180 3612 147186 3664
rect 155218 3612 155224 3664
rect 155276 3652 155282 3664
rect 160094 3652 160100 3664
rect 155276 3624 160100 3652
rect 155276 3612 155282 3624
rect 160094 3612 160100 3624
rect 160152 3612 160158 3664
rect 160738 3612 160744 3664
rect 160796 3652 160802 3664
rect 173158 3652 173164 3664
rect 160796 3624 173164 3652
rect 160796 3612 160802 3624
rect 173158 3612 173164 3624
rect 173216 3612 173222 3664
rect 173250 3612 173256 3664
rect 173308 3652 173314 3664
rect 461578 3652 461584 3664
rect 173308 3624 461584 3652
rect 173308 3612 173314 3624
rect 461578 3612 461584 3624
rect 461636 3612 461642 3664
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 117682 3584 117688 3596
rect 2924 3556 117688 3584
rect 2924 3544 2930 3556
rect 117682 3544 117688 3556
rect 117740 3544 117746 3596
rect 119890 3544 119896 3596
rect 119948 3584 119954 3596
rect 122098 3584 122104 3596
rect 119948 3556 122104 3584
rect 119948 3544 119954 3556
rect 122098 3544 122104 3556
rect 122156 3544 122162 3596
rect 135254 3544 135260 3596
rect 135312 3584 135318 3596
rect 136082 3584 136088 3596
rect 135312 3556 136088 3584
rect 135312 3544 135318 3556
rect 136082 3544 136088 3556
rect 136140 3544 136146 3596
rect 140130 3544 140136 3596
rect 140188 3584 140194 3596
rect 140188 3556 142154 3584
rect 140188 3544 140194 3556
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 4798 3516 4804 3528
rect 624 3488 4804 3516
rect 624 3476 630 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 124858 3516 124864 3528
rect 6886 3488 124864 3516
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 6886 3448 6914 3488
rect 124858 3476 124864 3488
rect 124916 3476 124922 3528
rect 126974 3476 126980 3528
rect 127032 3516 127038 3528
rect 129090 3516 129096 3528
rect 127032 3488 129096 3516
rect 127032 3476 127038 3488
rect 129090 3476 129096 3488
rect 129148 3476 129154 3528
rect 140314 3476 140320 3528
rect 140372 3516 140378 3528
rect 141234 3516 141240 3528
rect 140372 3488 141240 3516
rect 140372 3476 140378 3488
rect 141234 3476 141240 3488
rect 141292 3476 141298 3528
rect 142126 3516 142154 3556
rect 144270 3544 144276 3596
rect 144328 3584 144334 3596
rect 162486 3584 162492 3596
rect 144328 3556 162492 3584
rect 144328 3544 144334 3556
rect 162486 3544 162492 3556
rect 162544 3544 162550 3596
rect 173342 3544 173348 3596
rect 173400 3584 173406 3596
rect 173400 3556 175596 3584
rect 173400 3544 173406 3556
rect 163682 3516 163688 3528
rect 142126 3488 163688 3516
rect 163682 3476 163688 3488
rect 163740 3476 163746 3528
rect 174538 3476 174544 3528
rect 174596 3516 174602 3528
rect 175458 3516 175464 3528
rect 174596 3488 175464 3516
rect 174596 3476 174602 3488
rect 175458 3476 175464 3488
rect 175516 3476 175522 3528
rect 175568 3516 175596 3556
rect 176654 3544 176660 3596
rect 176712 3584 176718 3596
rect 177850 3584 177856 3596
rect 176712 3556 177856 3584
rect 176712 3544 176718 3556
rect 177850 3544 177856 3556
rect 177908 3544 177914 3596
rect 472250 3584 472256 3596
rect 177960 3556 472256 3584
rect 177960 3516 177988 3556
rect 472250 3544 472256 3556
rect 472308 3544 472314 3596
rect 479334 3516 479340 3528
rect 175568 3488 177988 3516
rect 178052 3488 479340 3516
rect 1728 3420 6914 3448
rect 1728 3408 1734 3420
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 124950 3448 124956 3460
rect 11204 3420 124956 3448
rect 11204 3408 11210 3420
rect 124950 3408 124956 3420
rect 125008 3408 125014 3460
rect 140038 3408 140044 3460
rect 140096 3448 140102 3460
rect 170766 3448 170772 3460
rect 140096 3420 170772 3448
rect 140096 3408 140102 3420
rect 170766 3408 170772 3420
rect 170824 3408 170830 3460
rect 173434 3408 173440 3460
rect 173492 3448 173498 3460
rect 178052 3448 178080 3488
rect 479334 3476 479340 3488
rect 479392 3476 479398 3528
rect 481634 3476 481640 3528
rect 481692 3516 481698 3528
rect 482462 3516 482468 3528
rect 481692 3488 482468 3516
rect 481692 3476 481698 3488
rect 482462 3476 482468 3488
rect 482520 3476 482526 3528
rect 514754 3476 514760 3528
rect 514812 3516 514818 3528
rect 515582 3516 515588 3528
rect 514812 3488 515588 3516
rect 514812 3476 514818 3488
rect 515582 3476 515588 3488
rect 515640 3476 515646 3528
rect 173492 3420 178080 3448
rect 173492 3408 173498 3420
rect 178126 3408 178132 3460
rect 178184 3448 178190 3460
rect 491110 3448 491116 3460
rect 178184 3420 491116 3448
rect 178184 3408 178190 3420
rect 491110 3408 491116 3420
rect 491168 3408 491174 3460
rect 44174 3340 44180 3392
rect 44232 3380 44238 3392
rect 45094 3380 45100 3392
rect 44232 3352 45100 3380
rect 44232 3340 44238 3352
rect 45094 3340 45100 3352
rect 45152 3340 45158 3392
rect 60734 3340 60740 3392
rect 60792 3380 60798 3392
rect 61654 3380 61660 3392
rect 60792 3352 61660 3380
rect 60792 3340 60798 3352
rect 61654 3340 61660 3352
rect 61712 3340 61718 3392
rect 93854 3340 93860 3392
rect 93912 3380 93918 3392
rect 94774 3380 94780 3392
rect 93912 3352 94780 3380
rect 93912 3340 93918 3352
rect 94774 3340 94780 3352
rect 94832 3340 94838 3392
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111610 3380 111616 3392
rect 110472 3352 111616 3380
rect 110472 3340 110478 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 142154 3340 142160 3392
rect 142212 3380 142218 3392
rect 218054 3380 218060 3392
rect 142212 3352 218060 3380
rect 142212 3340 142218 3352
rect 218054 3340 218060 3352
rect 218112 3340 218118 3392
rect 307754 3340 307760 3392
rect 307812 3380 307818 3392
rect 309042 3380 309048 3392
rect 307812 3352 309048 3380
rect 307812 3340 307818 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 324406 3340 324412 3392
rect 324464 3380 324470 3392
rect 325602 3380 325608 3392
rect 324464 3352 325608 3380
rect 324464 3340 324470 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 349246 3340 349252 3392
rect 349304 3380 349310 3392
rect 350442 3380 350448 3392
rect 349304 3352 350448 3380
rect 349304 3340 349310 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 357434 3340 357440 3392
rect 357492 3380 357498 3392
rect 358722 3380 358728 3392
rect 357492 3352 358728 3380
rect 357492 3340 357498 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 365714 3340 365720 3392
rect 365772 3380 365778 3392
rect 367002 3380 367008 3392
rect 365772 3352 367008 3380
rect 365772 3340 365778 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382274 3340 382280 3392
rect 382332 3380 382338 3392
rect 383562 3380 383568 3392
rect 382332 3352 383568 3380
rect 382332 3340 382338 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 390554 3340 390560 3392
rect 390612 3380 390618 3392
rect 391842 3380 391848 3392
rect 390612 3352 391848 3380
rect 390612 3340 390618 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 407206 3340 407212 3392
rect 407264 3380 407270 3392
rect 408402 3380 408408 3392
rect 407264 3352 408408 3380
rect 407264 3340 407270 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 138842 3272 138848 3324
rect 138900 3312 138906 3324
rect 150618 3312 150624 3324
rect 138900 3284 150624 3312
rect 138900 3272 138906 3284
rect 150618 3272 150624 3284
rect 150676 3272 150682 3324
rect 200298 3312 200304 3324
rect 178236 3284 200304 3312
rect 138750 3204 138756 3256
rect 138808 3244 138814 3256
rect 149514 3244 149520 3256
rect 138808 3216 149520 3244
rect 138808 3204 138814 3216
rect 149514 3204 149520 3216
rect 149572 3204 149578 3256
rect 172238 3204 172244 3256
rect 172296 3244 172302 3256
rect 178236 3244 178264 3284
rect 200298 3272 200304 3284
rect 200356 3272 200362 3324
rect 172296 3216 178264 3244
rect 172296 3204 172302 3216
rect 181438 3204 181444 3256
rect 181496 3244 181502 3256
rect 186222 3244 186228 3256
rect 181496 3216 186228 3244
rect 181496 3204 181502 3216
rect 186222 3204 186228 3216
rect 186280 3204 186286 3256
rect 118786 3136 118792 3188
rect 118844 3176 118850 3188
rect 120718 3176 120724 3188
rect 118844 3148 120724 3176
rect 118844 3136 118850 3148
rect 120718 3136 120724 3148
rect 120776 3136 120782 3188
rect 129366 3136 129372 3188
rect 129424 3176 129430 3188
rect 134610 3176 134616 3188
rect 129424 3148 134616 3176
rect 129424 3136 129430 3148
rect 134610 3136 134616 3148
rect 134668 3136 134674 3188
rect 135530 3136 135536 3188
rect 135588 3176 135594 3188
rect 137646 3176 137652 3188
rect 135588 3148 137652 3176
rect 135588 3136 135594 3148
rect 137646 3136 137652 3148
rect 137704 3136 137710 3188
rect 144454 3136 144460 3188
rect 144512 3176 144518 3188
rect 153010 3176 153016 3188
rect 144512 3148 153016 3176
rect 144512 3136 144518 3148
rect 153010 3136 153016 3148
rect 153068 3136 153074 3188
rect 172054 3136 172060 3188
rect 172112 3176 172118 3188
rect 182542 3176 182548 3188
rect 172112 3148 182548 3176
rect 172112 3136 172118 3148
rect 182542 3136 182548 3148
rect 182600 3136 182606 3188
rect 135438 3068 135444 3120
rect 135496 3108 135502 3120
rect 138842 3108 138848 3120
rect 135496 3080 138848 3108
rect 135496 3068 135502 3080
rect 138842 3068 138848 3080
rect 138900 3068 138906 3120
rect 153838 3068 153844 3120
rect 153896 3108 153902 3120
rect 161290 3108 161296 3120
rect 153896 3080 161296 3108
rect 153896 3068 153902 3080
rect 161290 3068 161296 3080
rect 161348 3068 161354 3120
rect 432046 2048 432052 2100
rect 432104 2088 432110 2100
rect 433242 2088 433248 2100
rect 432104 2060 433248 2088
rect 432104 2048 432110 2060
rect 433242 2048 433248 2060
rect 433300 2048 433306 2100
rect 415394 1912 415400 1964
rect 415452 1952 415458 1964
rect 416682 1952 416688 1964
rect 415452 1924 416688 1952
rect 415452 1912 415458 1924
rect 416682 1912 416688 1924
rect 416740 1912 416746 1964
rect 440234 1912 440240 1964
rect 440292 1952 440298 1964
rect 441522 1952 441528 1964
rect 440292 1924 441528 1952
rect 440292 1912 440298 1924
rect 441522 1912 441528 1924
rect 441580 1912 441586 1964
rect 456794 1912 456800 1964
rect 456852 1952 456858 1964
rect 458082 1952 458088 1964
rect 456852 1924 458088 1952
rect 456852 1912 456858 1924
rect 458082 1912 458088 1924
rect 458140 1912 458146 1964
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 405004 700408 405056 700460
rect 413652 700408 413704 700460
rect 364984 700340 365036 700392
rect 397552 700340 397604 700392
rect 403624 700340 403676 700392
rect 478512 700340 478564 700392
rect 292580 700272 292632 700324
rect 300124 700272 300176 700324
rect 348792 700272 348844 700324
rect 396632 700272 396684 700324
rect 400864 700272 400916 700324
rect 543464 700272 543516 700324
rect 233884 697552 233936 697604
rect 235172 697552 235224 697604
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 284944 697552 284996 697604
rect 292580 697552 292632 697604
rect 182180 694764 182232 694816
rect 201500 694764 201552 694816
rect 160744 692044 160796 692096
rect 169668 692044 169720 692096
rect 180064 690208 180116 690260
rect 182180 690208 182232 690260
rect 279424 687488 279476 687540
rect 284944 687488 284996 687540
rect 230848 684428 230900 684480
rect 233884 684496 233936 684548
rect 2780 683680 2832 683732
rect 4804 683680 4856 683732
rect 399484 683136 399536 683188
rect 580172 683136 580224 683188
rect 229744 681708 229796 681760
rect 230848 681708 230900 681760
rect 147772 678036 147824 678088
rect 153200 678036 153252 678088
rect 147036 675520 147088 675572
rect 147772 675520 147824 675572
rect 272524 674840 272576 674892
rect 279424 674840 279476 674892
rect 159456 674772 159508 674824
rect 160744 674772 160796 674824
rect 266360 674092 266412 674144
rect 275284 674092 275336 674144
rect 413284 670692 413336 670744
rect 580172 670692 580224 670744
rect 157340 668584 157392 668636
rect 159456 668584 159508 668636
rect 145564 667836 145616 667888
rect 147036 667836 147088 667888
rect 150440 665796 150492 665848
rect 157340 665796 157392 665848
rect 228364 663756 228416 663808
rect 229744 663756 229796 663808
rect 146944 662396 146996 662448
rect 150440 662396 150492 662448
rect 173164 662396 173216 662448
rect 180064 662396 180116 662448
rect 275284 661852 275336 661904
rect 278044 661852 278096 661904
rect 260104 658928 260156 658980
rect 272524 658928 272576 658980
rect 215944 658180 215996 658232
rect 218060 658180 218112 658232
rect 142804 657976 142856 658028
rect 145564 657976 145616 658028
rect 331220 655732 331272 655784
rect 335360 655732 335412 655784
rect 282920 653692 282972 653744
rect 286324 653692 286376 653744
rect 138388 652672 138440 652724
rect 142804 652740 142856 652792
rect 167000 652740 167052 652792
rect 173164 652740 173216 652792
rect 222844 652740 222896 652792
rect 228364 652740 228416 652792
rect 335360 652740 335412 652792
rect 341524 652740 341576 652792
rect 278044 652060 278096 652112
rect 281448 652060 281500 652112
rect 165344 650020 165396 650072
rect 167000 650020 167052 650072
rect 213184 650020 213236 650072
rect 215944 650020 215996 650072
rect 281448 647164 281500 647216
rect 285680 647164 285732 647216
rect 159364 646484 159416 646536
rect 165344 646484 165396 646536
rect 135904 644376 135956 644428
rect 138388 644444 138440 644496
rect 285680 642404 285732 642456
rect 289084 642404 289136 642456
rect 286324 642336 286376 642388
rect 294604 642336 294656 642388
rect 221556 640296 221608 640348
rect 222844 640296 222896 640348
rect 133144 639548 133196 639600
rect 159364 639548 159416 639600
rect 210424 638596 210476 638648
rect 213184 638596 213236 638648
rect 220084 638392 220136 638444
rect 221556 638392 221608 638444
rect 3332 632068 3384 632120
rect 7564 632068 7616 632120
rect 133236 630640 133288 630692
rect 135904 630640 135956 630692
rect 531964 630640 532016 630692
rect 579988 630640 580040 630692
rect 289084 630164 289136 630216
rect 295340 630164 295392 630216
rect 254584 626560 254636 626612
rect 260104 626560 260156 626612
rect 341524 626560 341576 626612
rect 347044 626560 347096 626612
rect 295340 625540 295392 625592
rect 298100 625540 298152 625592
rect 129740 623772 129792 623824
rect 133236 623772 133288 623824
rect 113824 623024 113876 623076
rect 133144 623024 133196 623076
rect 129004 620984 129056 621036
rect 129740 620984 129792 621036
rect 298100 620304 298152 620356
rect 305644 620304 305696 620356
rect 145564 618876 145616 618928
rect 146944 618876 146996 618928
rect 108304 611940 108356 611992
rect 113824 611940 113876 611992
rect 143540 608472 143592 608524
rect 145564 608472 145616 608524
rect 294604 607860 294656 607912
rect 300124 607860 300176 607912
rect 305644 606432 305696 606484
rect 310888 606432 310940 606484
rect 142804 604460 142856 604512
rect 143540 604460 143592 604512
rect 310888 600244 310940 600296
rect 315304 600244 315356 600296
rect 79324 592628 79376 592680
rect 108304 592628 108356 592680
rect 347044 592560 347096 592612
rect 353944 592560 353996 592612
rect 249064 587188 249116 587240
rect 254584 587188 254636 587240
rect 315304 587120 315356 587172
rect 319076 587120 319128 587172
rect 141424 586508 141476 586560
rect 142804 586508 142856 586560
rect 319076 582972 319128 583024
rect 333980 582972 334032 583024
rect 218704 580932 218756 580984
rect 220084 580932 220136 580984
rect 3332 579776 3384 579828
rect 8944 579776 8996 579828
rect 333980 577464 334032 577516
rect 340144 577464 340196 577516
rect 353944 577464 353996 577516
rect 360844 577464 360896 577516
rect 530584 576852 530636 576904
rect 580172 576852 580224 576904
rect 109684 576104 109736 576156
rect 141424 576104 141476 576156
rect 204904 573248 204956 573300
rect 210424 573248 210476 573300
rect 300124 572908 300176 572960
rect 302884 572908 302936 572960
rect 340144 569168 340196 569220
rect 352564 569168 352616 569220
rect 302884 562980 302936 563032
rect 307024 562980 307076 563032
rect 202144 562300 202196 562352
rect 204904 562300 204956 562352
rect 108304 561008 108356 561060
rect 109684 561008 109736 561060
rect 239404 560940 239456 560992
rect 249064 560940 249116 560992
rect 106280 556180 106332 556232
rect 108304 556180 108356 556232
rect 195980 556180 196032 556232
rect 202144 556180 202196 556232
rect 104164 551488 104216 551540
rect 106280 551488 106332 551540
rect 191196 550808 191248 550860
rect 195980 550808 196032 550860
rect 188344 547884 188396 547936
rect 191196 547884 191248 547936
rect 352564 547136 352616 547188
rect 364984 547136 365036 547188
rect 217416 545096 217468 545148
rect 218704 545096 218756 545148
rect 215944 542988 215996 543040
rect 217416 542988 217468 543040
rect 233884 542308 233936 542360
rect 239404 542308 239456 542360
rect 127624 540880 127676 540932
rect 129004 540880 129056 540932
rect 214564 535440 214616 535492
rect 215944 535440 215996 535492
rect 307024 534692 307076 534744
rect 344284 534692 344336 534744
rect 126244 529864 126296 529916
rect 127624 529864 127676 529916
rect 360844 528572 360896 528624
rect 366364 528572 366416 528624
rect 2964 527144 3016 527196
rect 10324 527144 10376 527196
rect 101404 527144 101456 527196
rect 104164 527144 104216 527196
rect 526444 524424 526496 524476
rect 580172 524424 580224 524476
rect 185584 523472 185636 523524
rect 188344 523472 188396 523524
rect 124220 520208 124272 520260
rect 126244 520208 126296 520260
rect 225604 519528 225656 519580
rect 233884 519528 233936 519580
rect 344284 519528 344336 519580
rect 349712 519528 349764 519580
rect 176660 518168 176712 518220
rect 185584 518168 185636 518220
rect 98644 516128 98696 516180
rect 101404 516128 101456 516180
rect 3332 514768 3384 514820
rect 25504 514768 25556 514820
rect 123484 514768 123536 514820
rect 124220 514768 124272 514820
rect 349712 514700 349764 514752
rect 355324 514700 355376 514752
rect 163504 514020 163556 514072
rect 176660 514020 176712 514072
rect 211804 513272 211856 513324
rect 214564 513272 214616 513324
rect 210424 508512 210476 508564
rect 225604 508512 225656 508564
rect 157984 507832 158036 507884
rect 163504 507832 163556 507884
rect 3240 500964 3292 501016
rect 43444 500964 43496 501016
rect 203524 498176 203576 498228
rect 210424 498176 210476 498228
rect 366364 494708 366416 494760
rect 374644 494708 374696 494760
rect 73160 487772 73212 487824
rect 79324 487772 79376 487824
rect 355324 485800 355376 485852
rect 359832 485800 359884 485852
rect 149704 485052 149756 485104
rect 157984 485052 158036 485104
rect 374644 485052 374696 485104
rect 384028 485052 384080 485104
rect 65524 484372 65576 484424
rect 73160 484372 73212 484424
rect 384028 480904 384080 480956
rect 393964 480904 394016 480956
rect 359832 480700 359884 480752
rect 364340 480700 364392 480752
rect 364340 476076 364392 476128
rect 370596 476076 370648 476128
rect 3056 474716 3108 474768
rect 18604 474716 18656 474768
rect 97264 473016 97316 473068
rect 98644 473016 98696 473068
rect 525064 470568 525116 470620
rect 579988 470568 580040 470620
rect 364984 469820 365036 469872
rect 370504 469820 370556 469872
rect 95884 469208 95936 469260
rect 97264 469208 97316 469260
rect 393964 469208 394016 469260
rect 396540 469208 396592 469260
rect 370596 465944 370648 465996
rect 373264 465944 373316 465996
rect 210424 463360 210476 463412
rect 211804 463360 211856 463412
rect 3332 462340 3384 462392
rect 28264 462340 28316 462392
rect 141424 461592 141476 461644
rect 149704 461592 149756 461644
rect 373264 453296 373316 453348
rect 393964 453296 394016 453348
rect 62120 452616 62172 452668
rect 65524 452616 65576 452668
rect 49608 449148 49660 449200
rect 62120 449148 62172 449200
rect 3332 448536 3384 448588
rect 37924 448536 37976 448588
rect 45008 446360 45060 446412
rect 49608 446360 49660 446412
rect 94504 445680 94556 445732
rect 95884 445680 95936 445732
rect 208400 438880 208452 438932
rect 210424 438880 210476 438932
rect 207664 435344 207716 435396
rect 208400 435344 208452 435396
rect 396724 430584 396776 430636
rect 580080 430584 580132 430636
rect 200672 429156 200724 429208
rect 203524 429156 203576 429208
rect 370504 424328 370556 424380
rect 389824 424328 389876 424380
rect 2964 422288 3016 422340
rect 13084 422288 13136 422340
rect 93124 422288 93176 422340
rect 94504 422288 94556 422340
rect 198004 422288 198056 422340
rect 200672 422288 200724 422340
rect 122104 420180 122156 420232
rect 123484 420180 123536 420232
rect 410524 418140 410576 418192
rect 580080 418140 580132 418192
rect 193864 415352 193916 415404
rect 198004 415352 198056 415404
rect 91100 413924 91152 413976
rect 93124 413924 93176 413976
rect 3332 409844 3384 409896
rect 32404 409844 32456 409896
rect 87696 408416 87748 408468
rect 91100 408484 91152 408536
rect 84200 405628 84252 405680
rect 87696 405696 87748 405748
rect 203892 404268 203944 404320
rect 207664 404336 207716 404388
rect 417424 404336 417476 404388
rect 580080 404336 580132 404388
rect 393964 404268 394016 404320
rect 397000 404268 397052 404320
rect 131764 402228 131816 402280
rect 141424 402228 141476 402280
rect 84200 401616 84252 401668
rect 119344 401616 119396 401668
rect 122104 401616 122156 401668
rect 82452 401548 82504 401600
rect 389824 399100 389876 399152
rect 392584 399100 392636 399152
rect 116584 398828 116636 398880
rect 119344 398828 119396 398880
rect 201408 397672 201460 397724
rect 203892 397672 203944 397724
rect 3332 397468 3384 397520
rect 39304 397468 39356 397520
rect 80704 397468 80756 397520
rect 82452 397468 82504 397520
rect 69664 396720 69716 396772
rect 136640 396720 136692 396772
rect 198740 393320 198792 393372
rect 201408 393320 201460 393372
rect 194508 389172 194560 389224
rect 198740 389172 198792 389224
rect 73804 388424 73856 388476
rect 80704 388424 80756 388476
rect 68284 384956 68336 385008
rect 69664 384956 69716 385008
rect 191840 384616 191892 384668
rect 194508 384616 194560 384668
rect 177304 384276 177356 384328
rect 193864 384276 193916 384328
rect 189724 382236 189776 382288
rect 191840 382236 191892 382288
rect 396816 378156 396868 378208
rect 580080 378156 580132 378208
rect 3332 371220 3384 371272
rect 14464 371220 14516 371272
rect 392584 371152 392636 371204
rect 395344 371152 395396 371204
rect 114928 370744 114980 370796
rect 116584 370744 116636 370796
rect 71044 369860 71096 369912
rect 73804 369860 73856 369912
rect 112444 367752 112496 367804
rect 114928 367752 114980 367804
rect 409144 364352 409196 364404
rect 579804 364352 579856 364404
rect 69664 362924 69716 362976
rect 71044 362924 71096 362976
rect 186320 362856 186372 362908
rect 189724 362924 189776 362976
rect 182364 360136 182416 360188
rect 186320 360204 186372 360256
rect 65432 358776 65484 358828
rect 68284 358776 68336 358828
rect 64144 358096 64196 358148
rect 65432 358096 65484 358148
rect 3332 357416 3384 357468
rect 26884 357416 26936 357468
rect 123484 357008 123536 357060
rect 131764 357008 131816 357060
rect 179420 354628 179472 354680
rect 182364 354696 182416 354748
rect 111064 353268 111116 353320
rect 112444 353268 112496 353320
rect 414664 351908 414716 351960
rect 580080 351908 580132 351960
rect 175004 346332 175056 346384
rect 179420 346400 179472 346452
rect 3332 345040 3384 345092
rect 43536 345040 43588 345092
rect 66260 343612 66312 343664
rect 69664 343612 69716 343664
rect 109776 343612 109828 343664
rect 111064 343612 111116 343664
rect 117964 343612 118016 343664
rect 123484 343612 123536 343664
rect 108304 340008 108356 340060
rect 109776 340008 109828 340060
rect 171876 339464 171928 339516
rect 175004 339464 175056 339516
rect 64236 336744 64288 336796
rect 66168 336744 66220 336796
rect 165436 335452 165488 335504
rect 171876 335452 171928 335504
rect 162860 332596 162912 332648
rect 165436 332596 165488 332648
rect 79324 331848 79376 331900
rect 117964 331848 118016 331900
rect 157984 331168 158036 331220
rect 162860 331236 162912 331288
rect 68284 320832 68336 320884
rect 79324 320832 79376 320884
rect 154764 320084 154816 320136
rect 157984 320152 158036 320204
rect 166264 319404 166316 319456
rect 177304 319404 177356 319456
rect 62764 318860 62816 318912
rect 64144 318860 64196 318912
rect 3148 318792 3200 318844
rect 17224 318792 17276 318844
rect 153200 318384 153252 318436
rect 154764 318384 154816 318436
rect 152464 314644 152516 314696
rect 153200 314644 153252 314696
rect 407764 311856 407816 311908
rect 580080 311856 580132 311908
rect 153844 311108 153896 311160
rect 166264 311108 166316 311160
rect 102784 305600 102836 305652
rect 108304 305600 108356 305652
rect 61384 303628 61436 303680
rect 64236 303628 64288 303680
rect 133144 302880 133196 302932
rect 153844 302880 153896 302932
rect 61476 299412 61528 299464
rect 62764 299412 62816 299464
rect 400956 298120 401008 298172
rect 580080 298120 580132 298172
rect 60096 297712 60148 297764
rect 61384 297712 61436 297764
rect 60004 293972 60056 294024
rect 61476 293972 61528 294024
rect 124496 293224 124548 293276
rect 133144 293224 133196 293276
rect 65616 292544 65668 292596
rect 68284 292544 68336 292596
rect 58624 290504 58676 290556
rect 60096 290504 60148 290556
rect 65524 290436 65576 290488
rect 104900 290436 104952 290488
rect 101404 290368 101456 290420
rect 102784 290368 102836 290420
rect 122104 288396 122156 288448
rect 124496 288396 124548 288448
rect 50528 286288 50580 286340
rect 65616 286288 65668 286340
rect 56600 285676 56652 285728
rect 58624 285676 58676 285728
rect 57980 282888 58032 282940
rect 60004 282888 60056 282940
rect 55864 282072 55916 282124
rect 56600 282072 56652 282124
rect 45836 279216 45888 279268
rect 50528 279216 50580 279268
rect 54484 278740 54536 278792
rect 57888 278740 57940 278792
rect 62764 277992 62816 278044
rect 101404 277992 101456 278044
rect 118884 277584 118936 277636
rect 122104 277584 122156 277636
rect 63500 276020 63552 276072
rect 65524 276020 65576 276072
rect 53840 275272 53892 275324
rect 55864 275272 55916 275324
rect 112444 273912 112496 273964
rect 118884 273912 118936 273964
rect 50988 271872 51040 271924
rect 53840 271872 53892 271924
rect 396908 271872 396960 271924
rect 579804 271872 579856 271924
rect 58532 268608 58584 268660
rect 63408 268608 63460 268660
rect 46940 268064 46992 268116
rect 50988 268064 51040 268116
rect 3240 266364 3292 266416
rect 21364 266364 21416 266416
rect 53104 266364 53156 266416
rect 54484 266364 54536 266416
rect 56140 266364 56192 266416
rect 58532 266364 58584 266416
rect 45192 264120 45244 264172
rect 46848 264120 46900 264172
rect 151084 263236 151136 263288
rect 152464 263236 152516 263288
rect 54484 262760 54536 262812
rect 56140 262760 56192 262812
rect 60004 262760 60056 262812
rect 62764 262760 62816 262812
rect 93124 261468 93176 261520
rect 112444 261468 112496 261520
rect 406384 258068 406436 258120
rect 579988 258068 580040 258120
rect 57612 255280 57664 255332
rect 60004 255280 60056 255332
rect 143080 255280 143132 255332
rect 151084 255280 151136 255332
rect 3332 253920 3384 253972
rect 35164 253920 35216 253972
rect 49608 253920 49660 253972
rect 53104 253920 53156 253972
rect 140044 252288 140096 252340
rect 143080 252288 143132 252340
rect 50252 251132 50304 251184
rect 54484 251200 54536 251252
rect 46204 249296 46256 249348
rect 49608 249296 49660 249348
rect 51080 248344 51132 248396
rect 57612 248412 57664 248464
rect 45376 244876 45428 244928
rect 50988 244876 51040 244928
rect 80060 244876 80112 244928
rect 93124 244876 93176 244928
rect 138020 244400 138072 244452
rect 140044 244400 140096 244452
rect 399576 244264 399628 244316
rect 579988 244264 580040 244316
rect 47492 243176 47544 243228
rect 50252 243176 50304 243228
rect 44916 240864 44968 240916
rect 71780 240864 71832 240916
rect 45284 240796 45336 240848
rect 88340 240796 88392 240848
rect 45836 240728 45888 240780
rect 138020 240728 138072 240780
rect 45652 240592 45704 240644
rect 47492 240592 47544 240644
rect 2780 240320 2832 240372
rect 4896 240320 4948 240372
rect 45468 240184 45520 240236
rect 46204 240184 46256 240236
rect 395344 240048 395396 240100
rect 396448 240048 396500 240100
rect 45560 239368 45612 239420
rect 80060 239776 80112 239828
rect 44824 238824 44876 238876
rect 45744 238824 45796 238876
rect 45100 238756 45152 238808
rect 45836 238756 45888 238808
rect 45192 233180 45244 233232
rect 45836 233180 45888 233232
rect 45468 232908 45520 232960
rect 86224 232364 86276 232416
rect 394148 232364 394200 232416
rect 397000 232364 397052 232416
rect 393964 231820 394016 231872
rect 580080 231820 580132 231872
rect 3700 231140 3752 231192
rect 180800 231140 180852 231192
rect 384396 231140 384448 231192
rect 396448 231140 396500 231192
rect 45836 231072 45888 231124
rect 49700 231072 49752 231124
rect 118608 231072 118660 231124
rect 397552 231072 397604 231124
rect 45376 231004 45428 231056
rect 150440 231004 150492 231056
rect 86224 230800 86276 230852
rect 88892 230800 88944 230852
rect 45560 230460 45612 230512
rect 390560 230460 390612 230512
rect 394148 230460 394200 230512
rect 54484 230392 54536 230444
rect 163504 229780 163556 229832
rect 176660 229780 176712 229832
rect 45100 229712 45152 229764
rect 53104 229712 53156 229764
rect 120816 229712 120868 229764
rect 580724 229712 580776 229764
rect 150440 229440 150492 229492
rect 153200 229440 153252 229492
rect 49700 229100 49752 229152
rect 52460 229032 52512 229084
rect 166264 228420 166316 228472
rect 296720 228420 296772 228472
rect 53104 228352 53156 228404
rect 58900 228352 58952 228404
rect 117228 228352 117280 228404
rect 143540 228352 143592 228404
rect 161388 228352 161440 228404
rect 386512 228352 386564 228404
rect 391940 228352 391992 228404
rect 396540 228352 396592 228404
rect 3056 227740 3108 227792
rect 140044 227740 140096 227792
rect 144920 227740 144972 227792
rect 146484 227740 146536 227792
rect 44824 227196 44876 227248
rect 47400 227196 47452 227248
rect 120724 226992 120776 227044
rect 580172 226992 580224 227044
rect 153200 226516 153252 226568
rect 155960 226516 156012 226568
rect 52460 226312 52512 226364
rect 56692 226244 56744 226296
rect 387800 225020 387852 225072
rect 390468 225020 390520 225072
rect 88892 224952 88944 225004
rect 45008 224884 45060 224936
rect 47584 224884 47636 224936
rect 387064 224952 387116 225004
rect 391940 224952 391992 225004
rect 91100 224884 91152 224936
rect 58900 224204 58952 224256
rect 63500 224204 63552 224256
rect 118700 224204 118752 224256
rect 580816 224204 580868 224256
rect 155960 223524 156012 223576
rect 157984 223524 158036 223576
rect 56692 222164 56744 222216
rect 60648 222096 60700 222148
rect 383660 221824 383712 221876
rect 387800 221824 387852 221876
rect 47400 220736 47452 220788
rect 49608 220736 49660 220788
rect 63500 220124 63552 220176
rect 68284 220124 68336 220176
rect 3884 220056 3936 220108
rect 179512 220056 179564 220108
rect 91100 219444 91152 219496
rect 95148 219376 95200 219428
rect 54484 218220 54536 218272
rect 56692 218220 56744 218272
rect 382280 218084 382332 218136
rect 383660 218084 383712 218136
rect 192484 218016 192536 218068
rect 580172 218016 580224 218068
rect 60648 217744 60700 217796
rect 64144 217744 64196 217796
rect 95148 216588 95200 216640
rect 98092 216588 98144 216640
rect 49700 214752 49752 214804
rect 53104 214752 53156 214804
rect 3332 213936 3384 213988
rect 22744 213936 22796 213988
rect 98092 213868 98144 213920
rect 104164 213868 104216 213920
rect 56692 212440 56744 212492
rect 58716 212440 58768 212492
rect 104164 211760 104216 211812
rect 108304 211760 108356 211812
rect 378784 209720 378836 209772
rect 382280 209788 382332 209840
rect 4068 209040 4120 209092
rect 180892 209040 180944 209092
rect 58716 208360 58768 208412
rect 61384 208360 61436 208412
rect 157984 208360 158036 208412
rect 162124 208292 162176 208344
rect 53104 207000 53156 207052
rect 55864 206932 55916 206984
rect 384304 205708 384356 205760
rect 387064 205708 387116 205760
rect 122104 205640 122156 205692
rect 580172 205640 580224 205692
rect 45652 205164 45704 205216
rect 49608 205164 49660 205216
rect 64144 204212 64196 204264
rect 65524 204212 65576 204264
rect 155224 203532 155276 203584
rect 266360 203532 266412 203584
rect 49608 202784 49660 202836
rect 53840 202784 53892 202836
rect 153200 202104 153252 202156
rect 236000 202104 236052 202156
rect 47584 201424 47636 201476
rect 50344 201424 50396 201476
rect 155960 200744 156012 200796
rect 166264 200744 166316 200796
rect 140044 199384 140096 199436
rect 164240 199384 164292 199436
rect 148968 198024 149020 198076
rect 207020 198024 207072 198076
rect 159824 197956 159876 198008
rect 356060 197956 356112 198008
rect 376024 197344 376076 197396
rect 378784 197344 378836 197396
rect 53840 197276 53892 197328
rect 57704 197276 57756 197328
rect 65524 196664 65576 196716
rect 66904 196664 66956 196716
rect 158260 196596 158312 196648
rect 327080 196596 327132 196648
rect 162124 195984 162176 196036
rect 56600 195916 56652 195968
rect 138112 195916 138164 195968
rect 166264 195916 166316 195968
rect 86960 195848 87012 195900
rect 139400 195848 139452 195900
rect 150348 195644 150400 195696
rect 165436 195644 165488 195696
rect 379520 193740 379572 193792
rect 384396 193740 384448 193792
rect 57704 193128 57756 193180
rect 61752 193128 61804 193180
rect 151636 191088 151688 191140
rect 371884 191088 371936 191140
rect 379520 191088 379572 191140
rect 50344 190884 50396 190936
rect 57244 190884 57296 190936
rect 2964 187688 3016 187740
rect 119344 187688 119396 187740
rect 61752 184832 61804 184884
rect 64972 184832 65024 184884
rect 68284 184832 68336 184884
rect 72424 184832 72476 184884
rect 66904 183472 66956 183524
rect 68284 183472 68336 183524
rect 55864 182112 55916 182164
rect 58624 182112 58676 182164
rect 64972 181432 65024 181484
rect 75184 181432 75236 181484
rect 144460 180684 144512 180736
rect 146116 180684 146168 180736
rect 162124 180888 162176 180940
rect 161664 180548 161716 180600
rect 9588 180072 9640 180124
rect 136824 180276 136876 180328
rect 136640 180072 136692 180124
rect 141240 180072 141292 180124
rect 143540 179596 143592 179648
rect 72424 179324 72476 179376
rect 75736 179324 75788 179376
rect 122840 178780 122892 178832
rect 136640 178780 136692 178832
rect 121460 178644 121512 178696
rect 137008 178644 137060 178696
rect 144184 178644 144236 178696
rect 159088 178508 159140 178560
rect 161664 178508 161716 178560
rect 166264 178236 166316 178288
rect 167644 178236 167696 178288
rect 189724 178032 189776 178084
rect 580172 178032 580224 178084
rect 61384 177964 61436 178016
rect 65892 177964 65944 178016
rect 140780 177828 140832 177880
rect 141608 177828 141660 177880
rect 124220 177284 124272 177336
rect 137100 177284 137152 177336
rect 75736 176944 75788 176996
rect 77300 176944 77352 176996
rect 159088 176196 159140 176248
rect 3332 176060 3384 176112
rect 9588 176060 9640 176112
rect 125600 175992 125652 176044
rect 137192 175992 137244 176044
rect 128360 175924 128412 175976
rect 137284 175924 137336 175976
rect 355324 175924 355376 175976
rect 371884 175924 371936 175976
rect 159088 175584 159140 175636
rect 165528 174972 165580 175024
rect 163136 174700 163188 174752
rect 165528 174700 165580 174752
rect 3700 174088 3752 174140
rect 179420 174088 179472 174140
rect 77300 173884 77352 173936
rect 65892 173816 65944 173868
rect 66904 173816 66956 173868
rect 133880 173884 133932 173936
rect 135260 173884 135312 173936
rect 81348 173816 81400 173868
rect 140780 173816 140832 173868
rect 141608 173816 141660 173868
rect 131120 173204 131172 173256
rect 137376 173204 137428 173256
rect 126980 173136 127032 173188
rect 140780 173136 140832 173188
rect 135260 172388 135312 172440
rect 138940 172388 138992 172440
rect 132500 172184 132552 172236
rect 137468 172184 137520 172236
rect 138020 171912 138072 171964
rect 140964 171912 141016 171964
rect 160008 171028 160060 171080
rect 163872 171028 163924 171080
rect 57244 170076 57296 170128
rect 60648 170076 60700 170128
rect 35164 168988 35216 169040
rect 182272 168988 182324 169040
rect 68284 168580 68336 168632
rect 69756 168580 69808 168632
rect 60648 166608 60700 166660
rect 62120 166608 62172 166660
rect 130384 165588 130436 165640
rect 580172 165588 580224 165640
rect 69756 165520 69808 165572
rect 71044 165520 71096 165572
rect 81440 165520 81492 165572
rect 83464 165520 83516 165572
rect 163872 165520 163924 165572
rect 166264 165520 166316 165572
rect 167644 165520 167696 165572
rect 169024 165520 169076 165572
rect 26884 164840 26936 164892
rect 182364 164840 182416 164892
rect 162860 164772 162912 164824
rect 163596 164772 163648 164824
rect 75184 163480 75236 163532
rect 86224 163480 86276 163532
rect 345664 163480 345716 163532
rect 355324 163480 355376 163532
rect 3332 162868 3384 162920
rect 108396 162868 108448 162920
rect 66904 162800 66956 162852
rect 68284 162800 68336 162852
rect 62120 162188 62172 162240
rect 87604 162188 87656 162240
rect 32404 162120 32456 162172
rect 182732 162120 182784 162172
rect 3516 160692 3568 160744
rect 179604 160692 179656 160744
rect 373264 160012 373316 160064
rect 376024 160080 376076 160132
rect 58624 159400 58676 159452
rect 81440 159400 81492 159452
rect 23480 159332 23532 159384
rect 180984 159332 181036 159384
rect 81440 157972 81492 158024
rect 84752 157972 84804 158024
rect 83464 157292 83516 157344
rect 84844 157292 84896 157344
rect 84752 156612 84804 156664
rect 89076 156612 89128 156664
rect 118240 156612 118292 156664
rect 417424 156612 417476 156664
rect 118332 155184 118384 155236
rect 414664 155184 414716 155236
rect 87604 154504 87656 154556
rect 90364 154504 90416 154556
rect 118516 153824 118568 153876
rect 400956 153824 401008 153876
rect 71044 153144 71096 153196
rect 73804 153144 73856 153196
rect 118424 152464 118476 152516
rect 399576 152464 399628 152516
rect 381544 151852 381596 151904
rect 384304 151852 384356 151904
rect 181444 151784 181496 151836
rect 579988 151784 580040 151836
rect 118792 151036 118844 151088
rect 580540 151036 580592 151088
rect 165436 150900 165488 150952
rect 167736 150900 167788 150952
rect 89076 149812 89128 149864
rect 91008 149812 91060 149864
rect 319444 149744 319496 149796
rect 345664 149744 345716 149796
rect 121000 149676 121052 149728
rect 429200 149676 429252 149728
rect 86224 149200 86276 149252
rect 88984 149200 89036 149252
rect 3516 149064 3568 149116
rect 178684 149064 178736 149116
rect 91008 148996 91060 149048
rect 92480 148996 92532 149048
rect 166264 147296 166316 147348
rect 168380 147296 168432 147348
rect 169024 146888 169076 146940
rect 175188 146888 175240 146940
rect 108304 146208 108356 146260
rect 109684 146208 109736 146260
rect 118976 145528 119028 145580
rect 494060 145528 494112 145580
rect 373356 144236 373408 144288
rect 381544 144236 381596 144288
rect 118884 144168 118936 144220
rect 558920 144168 558972 144220
rect 175280 143556 175332 143608
rect 151820 143488 151872 143540
rect 157432 143488 157484 143540
rect 167736 143488 167788 143540
rect 169944 143488 169996 143540
rect 178224 143488 178276 143540
rect 164056 143420 164108 143472
rect 166080 143420 166132 143472
rect 137744 143148 137796 143200
rect 139400 143148 139452 143200
rect 162768 143080 162820 143132
rect 166172 143080 166224 143132
rect 162860 142944 162912 142996
rect 174636 142944 174688 142996
rect 150440 142876 150492 142928
rect 154580 142876 154632 142928
rect 164240 142876 164292 142928
rect 176200 142876 176252 142928
rect 92480 142808 92532 142860
rect 104900 142808 104952 142860
rect 118148 142808 118200 142860
rect 130384 142808 130436 142860
rect 163136 142808 163188 142860
rect 178040 142808 178092 142860
rect 149060 142128 149112 142180
rect 152740 142128 152792 142180
rect 45284 141516 45336 141568
rect 182456 141516 182508 141568
rect 28264 141448 28316 141500
rect 182548 141448 182600 141500
rect 104900 141380 104952 141432
rect 107660 141380 107712 141432
rect 117964 141380 118016 141432
rect 413284 141380 413336 141432
rect 107660 140088 107712 140140
rect 181536 140088 181588 140140
rect 25504 140020 25556 140072
rect 182640 140020 182692 140072
rect 88984 139476 89036 139528
rect 91376 139476 91428 139528
rect 118056 139476 118108 139528
rect 122104 139476 122156 139528
rect 3700 139408 3752 139460
rect 181076 139408 181128 139460
rect 316684 139408 316736 139460
rect 319444 139408 319496 139460
rect 178224 139340 178276 139392
rect 180156 139340 180208 139392
rect 178684 139272 178736 139324
rect 182180 139272 182232 139324
rect 188344 137980 188396 138032
rect 580172 137980 580224 138032
rect 21456 136688 21508 136740
rect 117320 136688 117372 136740
rect 3516 136620 3568 136672
rect 120908 136620 120960 136672
rect 3516 135940 3568 135992
rect 3700 135940 3752 135992
rect 90364 135872 90416 135924
rect 105544 135872 105596 135924
rect 97264 135260 97316 135312
rect 117320 135260 117372 135312
rect 18696 133900 18748 133952
rect 117320 133900 117372 133952
rect 108396 133832 108448 133884
rect 117412 133832 117464 133884
rect 91376 132812 91428 132864
rect 94228 132812 94280 132864
rect 22744 132404 22796 132456
rect 117320 132404 117372 132456
rect 84844 131724 84896 131776
rect 86316 131724 86368 131776
rect 369860 131112 369912 131164
rect 373264 131112 373316 131164
rect 21364 131044 21416 131096
rect 117320 131044 117372 131096
rect 86316 130840 86368 130892
rect 87604 130840 87656 130892
rect 109684 129752 109736 129804
rect 111064 129752 111116 129804
rect 17224 129684 17276 129736
rect 117320 129684 117372 129736
rect 355968 129004 356020 129056
rect 369860 129004 369912 129056
rect 14464 128256 14516 128308
rect 117320 128256 117372 128308
rect 68284 127576 68336 127628
rect 71044 127576 71096 127628
rect 328920 127576 328972 127628
rect 355968 127576 356020 127628
rect 13084 126896 13136 126948
rect 117320 126896 117372 126948
rect 94228 126828 94280 126880
rect 100024 126828 100076 126880
rect 105544 126828 105596 126880
rect 109684 126828 109736 126880
rect 326712 126012 326764 126064
rect 328920 126012 328972 126064
rect 180064 125604 180116 125656
rect 579804 125604 579856 125656
rect 73804 124788 73856 124840
rect 75828 124788 75880 124840
rect 322940 124448 322992 124500
rect 326712 124448 326764 124500
rect 18604 124108 18656 124160
rect 117320 124108 117372 124160
rect 367744 123632 367796 123684
rect 373356 123632 373408 123684
rect 304264 123428 304316 123480
rect 322940 123428 322992 123480
rect 10324 122748 10376 122800
rect 117320 122748 117372 122800
rect 109684 122476 109736 122528
rect 113824 122476 113876 122528
rect 87604 121796 87656 121848
rect 91008 121796 91060 121848
rect 8944 121388 8996 121440
rect 117320 121388 117372 121440
rect 7564 120028 7616 120080
rect 117320 120028 117372 120080
rect 91100 119892 91152 119944
rect 93124 119892 93176 119944
rect 181536 119824 181588 119876
rect 182272 119824 182324 119876
rect 75920 119076 75972 119128
rect 78588 119076 78640 119128
rect 4804 118600 4856 118652
rect 117320 118600 117372 118652
rect 71044 117920 71096 117972
rect 77300 117920 77352 117972
rect 40040 117240 40092 117292
rect 117320 117240 117372 117292
rect 77300 116016 77352 116068
rect 79324 116016 79376 116068
rect 100024 115880 100076 115932
rect 117320 115880 117372 115932
rect 180156 114520 180208 114572
rect 78588 114452 78640 114504
rect 117320 114452 117372 114504
rect 182180 114452 182232 114504
rect 93124 113092 93176 113144
rect 117320 113092 117372 113144
rect 79324 112412 79376 112464
rect 88248 112412 88300 112464
rect 180156 111800 180208 111852
rect 580172 111800 580224 111852
rect 2964 111732 3016 111784
rect 18696 111732 18748 111784
rect 88248 111732 88300 111784
rect 117320 111732 117372 111784
rect 111064 109012 111116 109064
rect 112444 109012 112496 109064
rect 113824 109012 113876 109064
rect 120632 109012 120684 109064
rect 183284 107584 183336 107636
rect 304264 107584 304316 107636
rect 183284 106224 183336 106276
rect 396632 106224 396684 106276
rect 183284 104796 183336 104848
rect 405004 104796 405056 104848
rect 183284 103436 183336 103488
rect 403624 103436 403676 103488
rect 112444 103096 112496 103148
rect 115388 103096 115440 103148
rect 183284 102076 183336 102128
rect 400864 102076 400916 102128
rect 183192 100648 183244 100700
rect 399484 100648 399536 100700
rect 115388 100308 115440 100360
rect 117320 100308 117372 100360
rect 182824 99356 182876 99408
rect 580172 99356 580224 99408
rect 183192 99288 183244 99340
rect 531964 99288 532016 99340
rect 117320 97928 117372 97980
rect 120816 97928 120868 97980
rect 183192 97928 183244 97980
rect 530584 97928 530636 97980
rect 183192 96568 183244 96620
rect 526444 96568 526496 96620
rect 183468 95140 183520 95192
rect 525064 95140 525116 95192
rect 183468 93780 183520 93832
rect 410524 93780 410576 93832
rect 183468 92420 183520 92472
rect 409144 92420 409196 92472
rect 183468 90992 183520 91044
rect 407764 90992 407816 91044
rect 183468 89632 183520 89684
rect 406384 89632 406436 89684
rect 305644 88952 305696 89004
rect 316684 88952 316736 89004
rect 183468 88272 183520 88324
rect 192484 88272 192536 88324
rect 182548 86504 182600 86556
rect 189724 86504 189776 86556
rect 182732 84872 182784 84924
rect 188344 84872 188396 84924
rect 3332 84192 3384 84244
rect 120264 84192 120316 84244
rect 293960 83444 294012 83496
rect 305644 83444 305696 83496
rect 178960 82084 179012 82136
rect 580264 82084 580316 82136
rect 179420 80792 179472 80844
rect 580448 80792 580500 80844
rect 118608 80724 118660 80776
rect 579988 80724 580040 80776
rect 120816 80588 120868 80640
rect 121828 80588 121880 80640
rect 125140 80316 125192 80368
rect 124772 80248 124824 80300
rect 124956 80180 125008 80232
rect 123576 80112 123628 80164
rect 123300 80044 123352 80096
rect 123208 79976 123260 80028
rect 122196 79908 122248 79960
rect 125738 79908 125790 79960
rect 126106 79908 126158 79960
rect 126290 79908 126342 79960
rect 126474 79908 126526 79960
rect 124864 79772 124916 79824
rect 125646 79772 125698 79824
rect 43536 79704 43588 79756
rect 116860 79704 116912 79756
rect 123024 79704 123076 79756
rect 126198 79840 126250 79892
rect 126244 79704 126296 79756
rect 126750 79908 126802 79960
rect 126566 79840 126618 79892
rect 126658 79840 126710 79892
rect 126520 79704 126572 79756
rect 126612 79636 126664 79688
rect 39304 79568 39356 79620
rect 125140 79568 125192 79620
rect 126152 79568 126204 79620
rect 126336 79568 126388 79620
rect 120908 79500 120960 79552
rect 125600 79500 125652 79552
rect 125692 79500 125744 79552
rect 126796 79500 126848 79552
rect 127210 79908 127262 79960
rect 127486 79908 127538 79960
rect 127302 79840 127354 79892
rect 127394 79840 127446 79892
rect 127118 79772 127170 79824
rect 127072 79636 127124 79688
rect 127762 79840 127814 79892
rect 127440 79704 127492 79756
rect 127348 79636 127400 79688
rect 127624 79568 127676 79620
rect 127716 79568 127768 79620
rect 116860 79432 116912 79484
rect 120264 79364 120316 79416
rect 126336 79432 126388 79484
rect 127946 79908 127998 79960
rect 128130 79908 128182 79960
rect 128498 79908 128550 79960
rect 128774 79908 128826 79960
rect 129234 79908 129286 79960
rect 130338 79908 130390 79960
rect 128314 79840 128366 79892
rect 128866 79840 128918 79892
rect 128084 79704 128136 79756
rect 128360 79704 128412 79756
rect 128452 79704 128504 79756
rect 128728 79704 128780 79756
rect 127992 79636 128044 79688
rect 128268 79568 128320 79620
rect 129142 79840 129194 79892
rect 129418 79840 129470 79892
rect 129602 79840 129654 79892
rect 129694 79840 129746 79892
rect 129188 79704 129240 79756
rect 129556 79704 129608 79756
rect 129096 79636 129148 79688
rect 129878 79772 129930 79824
rect 128820 79500 128872 79552
rect 129556 79500 129608 79552
rect 129648 79500 129700 79552
rect 130522 79908 130574 79960
rect 130614 79908 130666 79960
rect 130982 79908 131034 79960
rect 131258 79908 131310 79960
rect 131350 79908 131402 79960
rect 131442 79908 131494 79960
rect 131994 79908 132046 79960
rect 132454 79908 132506 79960
rect 130016 79500 130068 79552
rect 3976 79296 4028 79348
rect 119344 79160 119396 79212
rect 129004 79364 129056 79416
rect 129556 79364 129608 79416
rect 130890 79772 130942 79824
rect 131258 79772 131310 79824
rect 130752 79500 130804 79552
rect 131304 79636 131356 79688
rect 131396 79568 131448 79620
rect 131488 79500 131540 79552
rect 132086 79840 132138 79892
rect 132362 79840 132414 79892
rect 132270 79772 132322 79824
rect 132224 79568 132276 79620
rect 132638 79908 132690 79960
rect 132730 79908 132782 79960
rect 133190 79908 133242 79960
rect 133466 79908 133518 79960
rect 133558 79908 133610 79960
rect 133742 79908 133794 79960
rect 133834 79908 133886 79960
rect 133926 79908 133978 79960
rect 134110 79908 134162 79960
rect 134294 79908 134346 79960
rect 134386 79908 134438 79960
rect 134478 79908 134530 79960
rect 132500 79772 132552 79824
rect 132592 79704 132644 79756
rect 132776 79636 132828 79688
rect 133098 79840 133150 79892
rect 133006 79772 133058 79824
rect 133052 79636 133104 79688
rect 133696 79704 133748 79756
rect 133880 79772 133932 79824
rect 134064 79772 134116 79824
rect 134156 79772 134208 79824
rect 133972 79704 134024 79756
rect 134248 79704 134300 79756
rect 133420 79636 133472 79688
rect 133512 79636 133564 79688
rect 133144 79568 133196 79620
rect 134754 79908 134806 79960
rect 134846 79908 134898 79960
rect 134938 79908 134990 79960
rect 132132 79500 132184 79552
rect 132316 79500 132368 79552
rect 132868 79500 132920 79552
rect 133788 79500 133840 79552
rect 134800 79772 134852 79824
rect 135398 79908 135450 79960
rect 135582 79908 135634 79960
rect 135766 79908 135818 79960
rect 135444 79772 135496 79824
rect 134708 79500 134760 79552
rect 135260 79500 135312 79552
rect 135628 79500 135680 79552
rect 136134 79908 136186 79960
rect 136226 79908 136278 79960
rect 137882 79908 137934 79960
rect 138526 79908 138578 79960
rect 138894 79908 138946 79960
rect 138986 79908 139038 79960
rect 139078 79908 139130 79960
rect 136042 79840 136094 79892
rect 135904 79636 135956 79688
rect 137146 79840 137198 79892
rect 137422 79840 137474 79892
rect 137606 79840 137658 79892
rect 136180 79636 136232 79688
rect 137100 79636 137152 79688
rect 138250 79840 138302 79892
rect 137928 79772 137980 79824
rect 138204 79704 138256 79756
rect 137560 79636 137612 79688
rect 137928 79636 137980 79688
rect 136088 79568 136140 79620
rect 138710 79772 138762 79824
rect 138848 79772 138900 79824
rect 138756 79636 138808 79688
rect 139216 79636 139268 79688
rect 138664 79568 138716 79620
rect 139032 79568 139084 79620
rect 139906 79908 139958 79960
rect 139722 79840 139774 79892
rect 140366 79908 140418 79960
rect 140458 79908 140510 79960
rect 140090 79840 140142 79892
rect 140182 79840 140234 79892
rect 139584 79636 139636 79688
rect 139768 79636 139820 79688
rect 130844 79432 130896 79484
rect 130568 79364 130620 79416
rect 133972 79432 134024 79484
rect 135168 79432 135220 79484
rect 139952 79636 140004 79688
rect 140550 79840 140602 79892
rect 140642 79840 140694 79892
rect 140412 79772 140464 79824
rect 140504 79704 140556 79756
rect 140734 79772 140786 79824
rect 140596 79636 140648 79688
rect 140320 79568 140372 79620
rect 141378 79908 141430 79960
rect 141654 79908 141706 79960
rect 141746 79908 141798 79960
rect 141838 79908 141890 79960
rect 142206 79908 142258 79960
rect 142298 79908 142350 79960
rect 142390 79908 142442 79960
rect 141010 79840 141062 79892
rect 141102 79840 141154 79892
rect 140872 79636 140924 79688
rect 140964 79568 141016 79620
rect 140136 79500 140188 79552
rect 140320 79432 140372 79484
rect 141562 79840 141614 79892
rect 141424 79636 141476 79688
rect 141976 79636 142028 79688
rect 142574 79908 142626 79960
rect 142666 79908 142718 79960
rect 143126 79908 143178 79960
rect 143218 79908 143270 79960
rect 143678 79908 143730 79960
rect 143862 79908 143914 79960
rect 144230 79908 144282 79960
rect 144414 79908 144466 79960
rect 142436 79772 142488 79824
rect 142528 79772 142580 79824
rect 142620 79772 142672 79824
rect 143172 79772 143224 79824
rect 142160 79636 142212 79688
rect 141700 79500 141752 79552
rect 141792 79432 141844 79484
rect 132684 79364 132736 79416
rect 139124 79364 139176 79416
rect 141148 79364 141200 79416
rect 142252 79568 142304 79620
rect 142344 79568 142396 79620
rect 143632 79704 143684 79756
rect 143724 79636 143776 79688
rect 144138 79840 144190 79892
rect 143954 79772 144006 79824
rect 144000 79636 144052 79688
rect 144184 79704 144236 79756
rect 144368 79704 144420 79756
rect 144690 79908 144742 79960
rect 145150 79908 145202 79960
rect 145242 79908 145294 79960
rect 145334 79908 145386 79960
rect 145426 79908 145478 79960
rect 145610 79908 145662 79960
rect 144782 79840 144834 79892
rect 144598 79772 144650 79824
rect 144460 79636 144512 79688
rect 145288 79772 145340 79824
rect 144736 79704 144788 79756
rect 145196 79704 145248 79756
rect 144644 79636 144696 79688
rect 145104 79636 145156 79688
rect 144552 79568 144604 79620
rect 145380 79568 145432 79620
rect 146162 79908 146214 79960
rect 145978 79840 146030 79892
rect 145748 79568 145800 79620
rect 146116 79636 146168 79688
rect 145932 79500 145984 79552
rect 146530 79908 146582 79960
rect 146484 79704 146536 79756
rect 146806 79908 146858 79960
rect 146898 79908 146950 79960
rect 147082 79908 147134 79960
rect 147818 79908 147870 79960
rect 148002 79908 148054 79960
rect 147542 79840 147594 79892
rect 146944 79636 146996 79688
rect 147128 79636 147180 79688
rect 147634 79772 147686 79824
rect 147588 79636 147640 79688
rect 146576 79568 146628 79620
rect 146852 79568 146904 79620
rect 148554 79908 148606 79960
rect 148646 79908 148698 79960
rect 149014 79908 149066 79960
rect 148370 79840 148422 79892
rect 148462 79840 148514 79892
rect 147956 79636 148008 79688
rect 148232 79636 148284 79688
rect 148048 79568 148100 79620
rect 147680 79500 147732 79552
rect 148738 79772 148790 79824
rect 149382 79908 149434 79960
rect 149658 79908 149710 79960
rect 149842 79908 149894 79960
rect 150486 79908 150538 79960
rect 150762 79908 150814 79960
rect 150854 79908 150906 79960
rect 150946 79908 150998 79960
rect 151038 79908 151090 79960
rect 151314 79908 151366 79960
rect 149290 79840 149342 79892
rect 148416 79636 148468 79688
rect 148692 79636 148744 79688
rect 148968 79636 149020 79688
rect 149152 79636 149204 79688
rect 149612 79704 149664 79756
rect 149428 79636 149480 79688
rect 149244 79568 149296 79620
rect 149934 79840 149986 79892
rect 150302 79840 150354 79892
rect 150026 79772 150078 79824
rect 149888 79636 149940 79688
rect 150256 79636 150308 79688
rect 149980 79568 150032 79620
rect 150532 79568 150584 79620
rect 150808 79568 150860 79620
rect 151406 79840 151458 79892
rect 151268 79704 151320 79756
rect 151360 79704 151412 79756
rect 151084 79568 151136 79620
rect 148600 79500 148652 79552
rect 150992 79500 151044 79552
rect 152050 79908 152102 79960
rect 152142 79908 152194 79960
rect 152418 79908 152470 79960
rect 152786 79908 152838 79960
rect 152878 79908 152930 79960
rect 152970 79908 153022 79960
rect 153154 79908 153206 79960
rect 153246 79908 153298 79960
rect 153338 79908 153390 79960
rect 153614 79908 153666 79960
rect 152050 79772 152102 79824
rect 152280 79636 152332 79688
rect 152510 79840 152562 79892
rect 152694 79840 152746 79892
rect 152556 79704 152608 79756
rect 152878 79772 152930 79824
rect 153062 79840 153114 79892
rect 152832 79636 152884 79688
rect 151912 79568 151964 79620
rect 152648 79568 152700 79620
rect 153016 79636 153068 79688
rect 152464 79500 152516 79552
rect 152740 79500 152792 79552
rect 152924 79500 152976 79552
rect 153706 79772 153758 79824
rect 153384 79704 153436 79756
rect 153660 79636 153712 79688
rect 154074 79908 154126 79960
rect 154166 79908 154218 79960
rect 154258 79908 154310 79960
rect 154350 79908 154402 79960
rect 154534 79908 154586 79960
rect 154810 79908 154862 79960
rect 154902 79908 154954 79960
rect 155270 79908 155322 79960
rect 155454 79908 155506 79960
rect 155546 79908 155598 79960
rect 153890 79840 153942 79892
rect 154028 79704 154080 79756
rect 153936 79636 153988 79688
rect 153752 79568 153804 79620
rect 153844 79500 153896 79552
rect 154212 79772 154264 79824
rect 154580 79772 154632 79824
rect 154718 79772 154770 79824
rect 154304 79704 154356 79756
rect 154488 79568 154540 79620
rect 155086 79840 155138 79892
rect 154856 79704 154908 79756
rect 155224 79772 155276 79824
rect 155316 79772 155368 79824
rect 155040 79704 155092 79756
rect 155132 79704 155184 79756
rect 155730 79840 155782 79892
rect 155914 79908 155966 79960
rect 156006 79908 156058 79960
rect 155868 79772 155920 79824
rect 155500 79636 155552 79688
rect 155684 79636 155736 79688
rect 154948 79568 155000 79620
rect 155408 79568 155460 79620
rect 155960 79568 156012 79620
rect 156374 79908 156426 79960
rect 156466 79908 156518 79960
rect 156328 79568 156380 79620
rect 155592 79500 155644 79552
rect 156650 79908 156702 79960
rect 156742 79908 156794 79960
rect 156834 79908 156886 79960
rect 156604 79704 156656 79756
rect 157202 79908 157254 79960
rect 157478 79908 157530 79960
rect 157662 79908 157714 79960
rect 157754 79908 157806 79960
rect 157938 79908 157990 79960
rect 156926 79840 156978 79892
rect 157018 79840 157070 79892
rect 156880 79636 156932 79688
rect 156512 79500 156564 79552
rect 156788 79568 156840 79620
rect 157294 79840 157346 79892
rect 157432 79772 157484 79824
rect 157156 79636 157208 79688
rect 157064 79568 157116 79620
rect 157524 79568 157576 79620
rect 156972 79500 157024 79552
rect 157846 79840 157898 79892
rect 157708 79772 157760 79824
rect 158030 79840 158082 79892
rect 174452 80588 174504 80640
rect 174544 80588 174596 80640
rect 580724 80656 580776 80708
rect 178040 80588 178092 80640
rect 580632 80588 580684 80640
rect 174728 80520 174780 80572
rect 158214 79772 158266 79824
rect 157892 79636 157944 79688
rect 158122 79636 158174 79688
rect 157984 79568 158036 79620
rect 158766 79840 158818 79892
rect 158490 79772 158542 79824
rect 158720 79704 158772 79756
rect 159042 79908 159094 79960
rect 159686 79908 159738 79960
rect 158444 79636 158496 79688
rect 158536 79636 158588 79688
rect 158076 79500 158128 79552
rect 158260 79500 158312 79552
rect 159410 79840 159462 79892
rect 159502 79840 159554 79892
rect 159594 79840 159646 79892
rect 159364 79636 159416 79688
rect 159456 79568 159508 79620
rect 159548 79568 159600 79620
rect 159364 79500 159416 79552
rect 160054 79840 160106 79892
rect 160146 79840 160198 79892
rect 160422 79840 160474 79892
rect 159870 79772 159922 79824
rect 159824 79636 159876 79688
rect 159916 79636 159968 79688
rect 160468 79704 160520 79756
rect 160698 79908 160750 79960
rect 160882 79908 160934 79960
rect 160974 79908 161026 79960
rect 161158 79840 161210 79892
rect 174636 80384 174688 80436
rect 554780 80316 554832 80368
rect 161342 79908 161394 79960
rect 161434 79908 161486 79960
rect 161112 79704 161164 79756
rect 161204 79704 161256 79756
rect 161020 79636 161072 79688
rect 160560 79568 160612 79620
rect 160744 79568 160796 79620
rect 161802 79908 161854 79960
rect 161894 79772 161946 79824
rect 161572 79636 161624 79688
rect 160652 79500 160704 79552
rect 161388 79500 161440 79552
rect 161848 79636 161900 79688
rect 162170 79908 162222 79960
rect 162630 79908 162682 79960
rect 162078 79840 162130 79892
rect 162262 79840 162314 79892
rect 144092 79432 144144 79484
rect 161572 79432 161624 79484
rect 161664 79432 161716 79484
rect 161940 79500 161992 79552
rect 162124 79432 162176 79484
rect 162446 79772 162498 79824
rect 174912 80248 174964 80300
rect 252560 80248 252612 80300
rect 174728 80180 174780 80232
rect 320180 80180 320232 80232
rect 163366 79908 163418 79960
rect 163642 79908 163694 79960
rect 163734 79908 163786 79960
rect 164286 79908 164338 79960
rect 164562 79908 164614 79960
rect 164746 79908 164798 79960
rect 163182 79840 163234 79892
rect 162676 79636 162728 79688
rect 162768 79636 162820 79688
rect 162400 79568 162452 79620
rect 163274 79772 163326 79824
rect 163550 79772 163602 79824
rect 163228 79636 163280 79688
rect 163320 79636 163372 79688
rect 163826 79840 163878 79892
rect 164194 79840 164246 79892
rect 163780 79704 163832 79756
rect 163596 79568 163648 79620
rect 163872 79636 163924 79688
rect 164424 79636 164476 79688
rect 164148 79568 164200 79620
rect 164930 79772 164982 79824
rect 164700 79704 164752 79756
rect 164884 79636 164936 79688
rect 165390 79908 165442 79960
rect 165482 79908 165534 79960
rect 165666 79908 165718 79960
rect 165850 79908 165902 79960
rect 166034 79908 166086 79960
rect 167414 79908 167466 79960
rect 165114 79840 165166 79892
rect 165298 79840 165350 79892
rect 164056 79500 164108 79552
rect 164976 79568 165028 79620
rect 165206 79772 165258 79824
rect 165482 79772 165534 79824
rect 165712 79772 165764 79824
rect 166862 79840 166914 79892
rect 166126 79772 166178 79824
rect 166310 79772 166362 79824
rect 165252 79636 165304 79688
rect 165528 79636 165580 79688
rect 165896 79636 165948 79688
rect 166540 79636 166592 79688
rect 167230 79772 167282 79824
rect 167276 79636 167328 79688
rect 168242 79908 168294 79960
rect 168702 79908 168754 79960
rect 168886 79908 168938 79960
rect 167598 79840 167650 79892
rect 167874 79772 167926 79824
rect 165160 79568 165212 79620
rect 165436 79568 165488 79620
rect 166816 79568 166868 79620
rect 167460 79568 167512 79620
rect 167828 79636 167880 79688
rect 168196 79772 168248 79824
rect 168288 79636 168340 79688
rect 168380 79636 168432 79688
rect 169990 79908 170042 79960
rect 170082 79908 170134 79960
rect 170174 79908 170226 79960
rect 170358 79908 170410 79960
rect 169162 79840 169214 79892
rect 169530 79840 169582 79892
rect 169622 79840 169674 79892
rect 169346 79772 169398 79824
rect 169438 79772 169490 79824
rect 169392 79636 169444 79688
rect 169484 79636 169536 79688
rect 169668 79636 169720 79688
rect 170128 79704 170180 79756
rect 170036 79636 170088 79688
rect 170220 79636 170272 79688
rect 170312 79636 170364 79688
rect 169116 79568 169168 79620
rect 169300 79568 169352 79620
rect 169576 79568 169628 79620
rect 164424 79500 164476 79552
rect 162492 79432 162544 79484
rect 169576 79432 169628 79484
rect 143540 79364 143592 79416
rect 159088 79364 159140 79416
rect 137284 79296 137336 79348
rect 126980 79228 127032 79280
rect 140780 79228 140832 79280
rect 142896 79296 142948 79348
rect 161296 79364 161348 79416
rect 169944 79296 169996 79348
rect 170910 79908 170962 79960
rect 170542 79840 170594 79892
rect 170726 79840 170778 79892
rect 171002 79772 171054 79824
rect 170588 79636 170640 79688
rect 171048 79636 171100 79688
rect 171370 79840 171422 79892
rect 174452 80112 174504 80164
rect 426440 80112 426492 80164
rect 171554 79908 171606 79960
rect 171416 79636 171468 79688
rect 171232 79568 171284 79620
rect 172106 79772 172158 79824
rect 171692 79636 171744 79688
rect 172750 79908 172802 79960
rect 172842 79908 172894 79960
rect 173302 79908 173354 79960
rect 173394 79908 173446 79960
rect 173578 79908 173630 79960
rect 172060 79568 172112 79620
rect 172612 79568 172664 79620
rect 172934 79840 172986 79892
rect 173026 79840 173078 79892
rect 172980 79704 173032 79756
rect 172888 79568 172940 79620
rect 173302 79704 173354 79756
rect 173486 79840 173538 79892
rect 177396 80044 177448 80096
rect 182180 80044 182232 80096
rect 184204 80044 184256 80096
rect 174130 79908 174182 79960
rect 174360 79908 174412 79960
rect 174636 79908 174688 79960
rect 173854 79772 173906 79824
rect 174452 79772 174504 79824
rect 498200 79840 498252 79892
rect 514760 79772 514812 79824
rect 173762 79704 173814 79756
rect 173348 79568 173400 79620
rect 173440 79568 173492 79620
rect 170772 79500 170824 79552
rect 173624 79500 173676 79552
rect 170864 79432 170916 79484
rect 171140 79432 171192 79484
rect 180156 79636 180208 79688
rect 170772 79296 170824 79348
rect 171784 79364 171836 79416
rect 181444 79364 181496 79416
rect 184940 79364 184992 79416
rect 580356 79364 580408 79416
rect 174360 79296 174412 79348
rect 177396 79296 177448 79348
rect 580908 79296 580960 79348
rect 146668 79228 146720 79280
rect 147680 79228 147732 79280
rect 157800 79228 157852 79280
rect 161572 79228 161624 79280
rect 164424 79228 164476 79280
rect 164700 79228 164752 79280
rect 128636 79160 128688 79212
rect 128912 79160 128964 79212
rect 129004 79160 129056 79212
rect 130844 79160 130896 79212
rect 131028 79160 131080 79212
rect 134340 79160 134392 79212
rect 135168 79160 135220 79212
rect 170404 79160 170456 79212
rect 171232 79228 171284 79280
rect 174084 79228 174136 79280
rect 174268 79228 174320 79280
rect 288440 79228 288492 79280
rect 173992 79160 174044 79212
rect 125968 79092 126020 79144
rect 126244 79092 126296 79144
rect 127256 79092 127308 79144
rect 137284 79092 137336 79144
rect 140780 79092 140832 79144
rect 142896 79092 142948 79144
rect 146668 79092 146720 79144
rect 126980 79024 127032 79076
rect 139124 79024 139176 79076
rect 143540 79024 143592 79076
rect 158352 79092 158404 79144
rect 161204 79092 161256 79144
rect 161572 79092 161624 79144
rect 161940 79092 161992 79144
rect 162216 79092 162268 79144
rect 324320 79092 324372 79144
rect 158812 79024 158864 79076
rect 159364 79024 159416 79076
rect 164700 79024 164752 79076
rect 135168 78956 135220 79008
rect 125600 78888 125652 78940
rect 127256 78888 127308 78940
rect 132684 78888 132736 78940
rect 144092 78956 144144 79008
rect 150440 78956 150492 79008
rect 150900 78956 150952 79008
rect 157800 78956 157852 79008
rect 166264 78956 166316 79008
rect 150992 78888 151044 78940
rect 158812 78888 158864 78940
rect 159364 78888 159416 78940
rect 172428 79024 172480 79076
rect 172704 79024 172756 79076
rect 293960 79024 294012 79076
rect 167368 78956 167420 79008
rect 167736 78956 167788 79008
rect 169300 78956 169352 79008
rect 169668 78956 169720 79008
rect 172520 78956 172572 79008
rect 367744 78956 367796 79008
rect 133604 78752 133656 78804
rect 138020 78752 138072 78804
rect 138112 78752 138164 78804
rect 138388 78752 138440 78804
rect 140320 78752 140372 78804
rect 140780 78752 140832 78804
rect 132684 78684 132736 78736
rect 132960 78684 133012 78736
rect 125048 78548 125100 78600
rect 133420 78616 133472 78668
rect 125416 78412 125468 78464
rect 133052 78412 133104 78464
rect 133512 78412 133564 78464
rect 146668 78684 146720 78736
rect 147036 78684 147088 78736
rect 138388 78616 138440 78668
rect 139952 78616 140004 78668
rect 140320 78616 140372 78668
rect 146484 78616 146536 78668
rect 147220 78616 147272 78668
rect 147680 78616 147732 78668
rect 147864 78616 147916 78668
rect 155868 78820 155920 78872
rect 160836 78820 160888 78872
rect 161204 78820 161256 78872
rect 165988 78820 166040 78872
rect 172796 78888 172848 78940
rect 172888 78888 172940 78940
rect 173900 78888 173952 78940
rect 174084 78888 174136 78940
rect 393964 78888 394016 78940
rect 159456 78752 159508 78804
rect 430580 78820 430632 78872
rect 169944 78752 169996 78804
rect 173348 78752 173400 78804
rect 151912 78684 151964 78736
rect 153108 78684 153160 78736
rect 154856 78684 154908 78736
rect 162400 78684 162452 78736
rect 151084 78616 151136 78668
rect 158812 78616 158864 78668
rect 158996 78616 159048 78668
rect 159088 78616 159140 78668
rect 161296 78616 161348 78668
rect 136548 78548 136600 78600
rect 144460 78548 144512 78600
rect 145288 78548 145340 78600
rect 166264 78616 166316 78668
rect 164976 78548 165028 78600
rect 165252 78548 165304 78600
rect 167000 78548 167052 78600
rect 174268 78684 174320 78736
rect 168840 78616 168892 78668
rect 170772 78616 170824 78668
rect 171876 78616 171928 78668
rect 178040 78616 178092 78668
rect 171600 78548 171652 78600
rect 396816 78548 396868 78600
rect 139492 78480 139544 78532
rect 171784 78480 171836 78532
rect 172060 78480 172112 78532
rect 178960 78480 179012 78532
rect 140688 78412 140740 78464
rect 195980 78412 196032 78464
rect 133696 78344 133748 78396
rect 140780 78344 140832 78396
rect 141332 78344 141384 78396
rect 145196 78344 145248 78396
rect 147312 78344 147364 78396
rect 150716 78344 150768 78396
rect 150900 78344 150952 78396
rect 159548 78344 159600 78396
rect 160008 78344 160060 78396
rect 160836 78344 160888 78396
rect 161020 78344 161072 78396
rect 161112 78344 161164 78396
rect 255964 78344 256016 78396
rect 132960 78276 133012 78328
rect 145840 78276 145892 78328
rect 150808 78276 150860 78328
rect 153660 78276 153712 78328
rect 157248 78276 157300 78328
rect 158628 78276 158680 78328
rect 158996 78276 159048 78328
rect 162584 78276 162636 78328
rect 315304 78276 315356 78328
rect 106924 78208 106976 78260
rect 127440 78208 127492 78260
rect 133696 78208 133748 78260
rect 137008 78208 137060 78260
rect 140872 78208 140924 78260
rect 141332 78208 141384 78260
rect 156420 78208 156472 78260
rect 161020 78208 161072 78260
rect 164792 78208 164844 78260
rect 341524 78208 341576 78260
rect 110420 78140 110472 78192
rect 123116 78140 123168 78192
rect 141056 78140 141108 78192
rect 89720 78072 89772 78124
rect 132500 78072 132552 78124
rect 140412 78072 140464 78124
rect 148784 78072 148836 78124
rect 71780 78004 71832 78056
rect 126152 78004 126204 78056
rect 132776 78004 132828 78056
rect 133328 78004 133380 78056
rect 149060 78140 149112 78192
rect 151544 78140 151596 78192
rect 152464 78140 152516 78192
rect 154856 78140 154908 78192
rect 155316 78140 155368 78192
rect 157340 78140 157392 78192
rect 157708 78140 157760 78192
rect 163688 78140 163740 78192
rect 480260 78140 480312 78192
rect 162216 78072 162268 78124
rect 163136 78072 163188 78124
rect 163504 78072 163556 78124
rect 167184 78072 167236 78124
rect 532700 78072 532752 78124
rect 152464 78004 152516 78056
rect 153476 78004 153528 78056
rect 153660 78004 153712 78056
rect 154488 78004 154540 78056
rect 155132 78004 155184 78056
rect 156512 78004 156564 78056
rect 53840 77936 53892 77988
rect 129740 77936 129792 77988
rect 123668 77868 123720 77920
rect 134708 77936 134760 77988
rect 139768 77936 139820 77988
rect 132868 77868 132920 77920
rect 133328 77868 133380 77920
rect 137652 77868 137704 77920
rect 140412 77868 140464 77920
rect 154580 77936 154632 77988
rect 155040 77936 155092 77988
rect 156052 77936 156104 77988
rect 156604 77936 156656 77988
rect 157708 77936 157760 77988
rect 157984 77936 158036 77988
rect 165988 78004 166040 78056
rect 170680 78004 170732 78056
rect 538864 78004 538916 78056
rect 131120 77800 131172 77852
rect 133880 77800 133932 77852
rect 140964 77800 141016 77852
rect 141700 77800 141752 77852
rect 143540 77800 143592 77852
rect 144368 77800 144420 77852
rect 149152 77800 149204 77852
rect 149888 77800 149940 77852
rect 153292 77800 153344 77852
rect 153752 77800 153804 77852
rect 155040 77732 155092 77784
rect 155408 77732 155460 77784
rect 157616 77732 157668 77784
rect 174452 77936 174504 77988
rect 171416 77868 171468 77920
rect 581000 77936 581052 77988
rect 171968 77800 172020 77852
rect 125140 77664 125192 77716
rect 134064 77664 134116 77716
rect 134524 77664 134576 77716
rect 135352 77664 135404 77716
rect 149428 77664 149480 77716
rect 149888 77664 149940 77716
rect 171876 77732 171928 77784
rect 171416 77664 171468 77716
rect 136640 77596 136692 77648
rect 139124 77596 139176 77648
rect 144920 77596 144972 77648
rect 157064 77596 157116 77648
rect 160100 77596 160152 77648
rect 171692 77596 171744 77648
rect 123116 77528 123168 77580
rect 131028 77528 131080 77580
rect 141792 77528 141844 77580
rect 172244 77528 172296 77580
rect 172796 77528 172848 77580
rect 396724 77528 396776 77580
rect 147956 77460 148008 77512
rect 167000 77460 167052 77512
rect 122932 77392 122984 77444
rect 130108 77392 130160 77444
rect 133880 77392 133932 77444
rect 135996 77392 136048 77444
rect 150532 77392 150584 77444
rect 158352 77392 158404 77444
rect 164424 77392 164476 77444
rect 169024 77460 169076 77512
rect 171784 77460 171836 77512
rect 178040 77460 178092 77512
rect 145012 77324 145064 77376
rect 145748 77324 145800 77376
rect 155868 77324 155920 77376
rect 156604 77324 156656 77376
rect 161112 77324 161164 77376
rect 172152 77324 172204 77376
rect 129004 77256 129056 77308
rect 131672 77256 131724 77308
rect 135720 77256 135772 77308
rect 135996 77256 136048 77308
rect 139952 77256 140004 77308
rect 140228 77256 140280 77308
rect 151912 77256 151964 77308
rect 152188 77256 152240 77308
rect 154212 77256 154264 77308
rect 157984 77256 158036 77308
rect 160652 77256 160704 77308
rect 166908 77256 166960 77308
rect 169024 77256 169076 77308
rect 171692 77256 171744 77308
rect 121828 77188 121880 77240
rect 123944 77188 123996 77240
rect 131396 77188 131448 77240
rect 131948 77188 132000 77240
rect 139492 77188 139544 77240
rect 140136 77188 140188 77240
rect 153476 77188 153528 77240
rect 154028 77188 154080 77240
rect 162216 77188 162268 77240
rect 197360 77188 197412 77240
rect 139308 77120 139360 77172
rect 140596 77120 140648 77172
rect 142252 77120 142304 77172
rect 213920 77120 213972 77172
rect 126980 77052 127032 77104
rect 129188 77052 129240 77104
rect 131304 77052 131356 77104
rect 132132 77052 132184 77104
rect 143172 77052 143224 77104
rect 226340 77052 226392 77104
rect 143448 76984 143500 77036
rect 231860 76984 231912 77036
rect 129188 76916 129240 76968
rect 129924 76916 129976 76968
rect 144184 76916 144236 76968
rect 240140 76916 240192 76968
rect 122104 76848 122156 76900
rect 134800 76848 134852 76900
rect 138296 76848 138348 76900
rect 138572 76848 138624 76900
rect 150808 76848 150860 76900
rect 260840 76848 260892 76900
rect 129924 76780 129976 76832
rect 130200 76780 130252 76832
rect 146300 76780 146352 76832
rect 267740 76780 267792 76832
rect 102140 76712 102192 76764
rect 132408 76712 132460 76764
rect 142252 76712 142304 76764
rect 142712 76712 142764 76764
rect 147772 76712 147824 76764
rect 284300 76712 284352 76764
rect 86960 76644 87012 76696
rect 132316 76644 132368 76696
rect 145104 76644 145156 76696
rect 145380 76644 145432 76696
rect 152556 76644 152608 76696
rect 153108 76644 153160 76696
rect 156144 76644 156196 76696
rect 156880 76644 156932 76696
rect 157524 76644 157576 76696
rect 296720 76644 296772 76696
rect 44180 76576 44232 76628
rect 120908 76576 120960 76628
rect 130200 76576 130252 76628
rect 130568 76576 130620 76628
rect 142344 76576 142396 76628
rect 142804 76576 142856 76628
rect 146024 76576 146076 76628
rect 146760 76576 146812 76628
rect 147956 76576 148008 76628
rect 148416 76576 148468 76628
rect 151544 76576 151596 76628
rect 30380 76508 30432 76560
rect 137560 76508 137612 76560
rect 144460 76508 144512 76560
rect 156328 76576 156380 76628
rect 156512 76576 156564 76628
rect 157432 76576 157484 76628
rect 158168 76576 158220 76628
rect 302240 76576 302292 76628
rect 171232 76508 171284 76560
rect 374000 76508 374052 76560
rect 126336 76440 126388 76492
rect 130108 76440 130160 76492
rect 130660 76440 130712 76492
rect 141148 76440 141200 76492
rect 141516 76440 141568 76492
rect 142160 76440 142212 76492
rect 142620 76440 142672 76492
rect 147772 76440 147824 76492
rect 148600 76440 148652 76492
rect 152464 76440 152516 76492
rect 162216 76440 162268 76492
rect 153200 76372 153252 76424
rect 157524 76372 157576 76424
rect 145380 76304 145432 76356
rect 145656 76304 145708 76356
rect 162492 76304 162544 76356
rect 173256 76304 173308 76356
rect 153200 76236 153252 76288
rect 153936 76236 153988 76288
rect 157524 76236 157576 76288
rect 158260 76236 158312 76288
rect 161940 76236 161992 76288
rect 162124 76236 162176 76288
rect 159088 76168 159140 76220
rect 159272 76168 159324 76220
rect 120908 76100 120960 76152
rect 128268 76100 128320 76152
rect 161756 76100 161808 76152
rect 162124 76100 162176 76152
rect 122288 76032 122340 76084
rect 127348 76032 127400 76084
rect 145104 76032 145156 76084
rect 145932 76032 145984 76084
rect 161572 76032 161624 76084
rect 167460 76032 167512 76084
rect 167920 76032 167972 76084
rect 155776 75964 155828 76016
rect 156972 75964 157024 76016
rect 161756 75964 161808 76016
rect 163136 75964 163188 76016
rect 163872 75964 163924 76016
rect 125876 75896 125928 75948
rect 126060 75896 126112 75948
rect 127256 75896 127308 75948
rect 127716 75896 127768 75948
rect 127900 75896 127952 75948
rect 128268 75896 128320 75948
rect 128912 75896 128964 75948
rect 129280 75896 129332 75948
rect 160100 75896 160152 75948
rect 160376 75896 160428 75948
rect 160468 75896 160520 75948
rect 160652 75896 160704 75948
rect 165804 75896 165856 75948
rect 166632 75896 166684 75948
rect 44916 75828 44968 75880
rect 173072 75828 173124 75880
rect 125048 75760 125100 75812
rect 125508 75760 125560 75812
rect 125600 75760 125652 75812
rect 172612 75760 172664 75812
rect 123944 75692 123996 75744
rect 171508 75692 171560 75744
rect 125876 75624 125928 75676
rect 126888 75624 126940 75676
rect 127348 75624 127400 75676
rect 127808 75624 127860 75676
rect 120724 75488 120776 75540
rect 133788 75624 133840 75676
rect 135444 75624 135496 75676
rect 136272 75624 136324 75676
rect 164700 75624 164752 75676
rect 165252 75624 165304 75676
rect 129740 75556 129792 75608
rect 135536 75556 135588 75608
rect 163044 75556 163096 75608
rect 163412 75556 163464 75608
rect 107660 75420 107712 75472
rect 131120 75488 131172 75540
rect 150992 75488 151044 75540
rect 322940 75488 322992 75540
rect 135536 75420 135588 75472
rect 136180 75420 136232 75472
rect 157248 75420 157300 75472
rect 361580 75420 361632 75472
rect 70400 75352 70452 75404
rect 130936 75352 130988 75404
rect 162952 75352 163004 75404
rect 163964 75352 164016 75404
rect 164148 75352 164200 75404
rect 60740 75284 60792 75336
rect 124956 75284 125008 75336
rect 137100 75284 137152 75336
rect 137284 75284 137336 75336
rect 138020 75284 138072 75336
rect 138480 75284 138532 75336
rect 160284 75284 160336 75336
rect 160836 75284 160888 75336
rect 164332 75284 164384 75336
rect 164700 75284 164752 75336
rect 166080 75284 166132 75336
rect 166724 75284 166776 75336
rect 166908 75352 166960 75404
rect 438860 75352 438912 75404
rect 490012 75284 490064 75336
rect 35900 75216 35952 75268
rect 6920 75148 6972 75200
rect 121092 75216 121144 75268
rect 125600 75216 125652 75268
rect 135812 75216 135864 75268
rect 136456 75216 136508 75268
rect 136824 75216 136876 75268
rect 137008 75216 137060 75268
rect 139400 75216 139452 75268
rect 139768 75216 139820 75268
rect 143632 75216 143684 75268
rect 144184 75216 144236 75268
rect 149244 75216 149296 75268
rect 149428 75216 149480 75268
rect 149520 75216 149572 75268
rect 149796 75216 149848 75268
rect 150808 75216 150860 75268
rect 151268 75216 151320 75268
rect 159180 75216 159232 75268
rect 159824 75216 159876 75268
rect 160376 75216 160428 75268
rect 160928 75216 160980 75268
rect 163044 75216 163096 75268
rect 163596 75216 163648 75268
rect 166264 75216 166316 75268
rect 166448 75216 166500 75268
rect 168472 75216 168524 75268
rect 168840 75216 168892 75268
rect 169944 75216 169996 75268
rect 170220 75216 170272 75268
rect 178684 75216 178736 75268
rect 506480 75216 506532 75268
rect 128360 75148 128412 75200
rect 135720 75148 135772 75200
rect 136364 75148 136416 75200
rect 136732 75148 136784 75200
rect 137100 75148 137152 75200
rect 138020 75148 138072 75200
rect 138664 75148 138716 75200
rect 150532 75148 150584 75200
rect 151176 75148 151228 75200
rect 164424 75148 164476 75200
rect 164976 75148 165028 75200
rect 165804 75148 165856 75200
rect 166540 75148 166592 75200
rect 169392 75148 169444 75200
rect 136824 75080 136876 75132
rect 137468 75080 137520 75132
rect 138204 75080 138256 75132
rect 138572 75080 138624 75132
rect 139400 75080 139452 75132
rect 140320 75080 140372 75132
rect 149244 75080 149296 75132
rect 149612 75080 149664 75132
rect 153016 75080 153068 75132
rect 154028 75080 154080 75132
rect 156328 75080 156380 75132
rect 156788 75080 156840 75132
rect 164332 75080 164384 75132
rect 164884 75080 164936 75132
rect 165160 75080 165212 75132
rect 178684 75080 178736 75132
rect 564440 75148 564492 75200
rect 123024 75012 123076 75064
rect 136732 75012 136784 75064
rect 137744 75012 137796 75064
rect 167092 75012 167144 75064
rect 167552 75012 167604 75064
rect 168472 75012 168524 75064
rect 169116 75012 169168 75064
rect 169760 75012 169812 75064
rect 170220 75012 170272 75064
rect 120816 74944 120868 74996
rect 128544 74944 128596 74996
rect 138204 74944 138256 74996
rect 138756 74944 138808 74996
rect 149612 74944 149664 74996
rect 149980 74944 150032 74996
rect 167092 74876 167144 74928
rect 167828 74876 167880 74928
rect 169760 74876 169812 74928
rect 170496 74876 170548 74928
rect 154672 74672 154724 74724
rect 155500 74672 155552 74724
rect 134616 74468 134668 74520
rect 135352 74468 135404 74520
rect 126244 74264 126296 74316
rect 129556 74264 129608 74316
rect 137928 74264 137980 74316
rect 142896 74264 142948 74316
rect 164056 74128 164108 74180
rect 173440 74128 173492 74180
rect 139216 74060 139268 74112
rect 173900 74060 173952 74112
rect 122840 73992 122892 74044
rect 135076 73992 135128 74044
rect 141976 73992 142028 74044
rect 209780 73992 209832 74044
rect 93952 73924 94004 73976
rect 133236 73924 133288 73976
rect 142988 73924 143040 73976
rect 223580 73924 223632 73976
rect 51080 73856 51132 73908
rect 129464 73856 129516 73908
rect 147312 73856 147364 73908
rect 251180 73856 251232 73908
rect 4804 73788 4856 73840
rect 125232 73788 125284 73840
rect 155316 73788 155368 73840
rect 357440 73788 357492 73840
rect 124772 73652 124824 73704
rect 125232 73652 125284 73704
rect 161480 73380 161532 73432
rect 161848 73380 161900 73432
rect 125048 73312 125100 73364
rect 127992 73312 128044 73364
rect 161848 73244 161900 73296
rect 162308 73244 162360 73296
rect 171140 73108 171192 73160
rect 580172 73108 580224 73160
rect 126152 73040 126204 73092
rect 126704 73040 126756 73092
rect 163780 72904 163832 72956
rect 173532 72904 173584 72956
rect 162032 72836 162084 72888
rect 181444 72836 181496 72888
rect 114560 72768 114612 72820
rect 133420 72768 133472 72820
rect 151084 72768 151136 72820
rect 325700 72768 325752 72820
rect 103520 72700 103572 72752
rect 133604 72700 133656 72752
rect 151452 72700 151504 72752
rect 332600 72700 332652 72752
rect 69020 72632 69072 72684
rect 130660 72632 130712 72684
rect 152004 72632 152056 72684
rect 340880 72632 340932 72684
rect 341524 72632 341576 72684
rect 465080 72632 465132 72684
rect 26240 72564 26292 72616
rect 127440 72564 127492 72616
rect 152740 72564 152792 72616
rect 347780 72564 347832 72616
rect 13820 72496 13872 72548
rect 123208 72496 123260 72548
rect 157984 72496 158036 72548
rect 368480 72496 368532 72548
rect 11060 72428 11112 72480
rect 126612 72428 126664 72480
rect 127440 72428 127492 72480
rect 128084 72428 128136 72480
rect 159456 72428 159508 72480
rect 382280 72428 382332 72480
rect 124956 72224 125008 72276
rect 125692 72224 125744 72276
rect 3424 71680 3476 71732
rect 97264 71680 97316 71732
rect 132684 71680 132736 71732
rect 135996 71680 136048 71732
rect 140596 71340 140648 71392
rect 176752 71340 176804 71392
rect 121460 71272 121512 71324
rect 134892 71272 134944 71324
rect 155592 71272 155644 71324
rect 367100 71272 367152 71324
rect 100760 71204 100812 71256
rect 133512 71204 133564 71256
rect 155224 71204 155276 71256
rect 382372 71204 382424 71256
rect 96620 71136 96672 71188
rect 133328 71136 133380 71188
rect 165252 71136 165304 71188
rect 505100 71136 505152 71188
rect 49700 71068 49752 71120
rect 126980 71068 127032 71120
rect 166632 71068 166684 71120
rect 518900 71068 518952 71120
rect 29000 71000 29052 71052
rect 128268 71000 128320 71052
rect 168288 71000 168340 71052
rect 539600 71000 539652 71052
rect 137284 70388 137336 70440
rect 138756 70388 138808 70440
rect 140044 70184 140096 70236
rect 184940 70184 184992 70236
rect 141516 70116 141568 70168
rect 209872 70116 209924 70168
rect 3424 70048 3476 70100
rect 174544 70048 174596 70100
rect 162400 69980 162452 70032
rect 375380 69980 375432 70032
rect 159364 69912 159416 69964
rect 437480 69912 437532 69964
rect 82820 69844 82872 69896
rect 131488 69844 131540 69896
rect 166356 69844 166408 69896
rect 523040 69844 523092 69896
rect 78680 69776 78732 69828
rect 131212 69776 131264 69828
rect 167736 69776 167788 69828
rect 536840 69776 536892 69828
rect 52460 69708 52512 69760
rect 128820 69708 128872 69760
rect 170772 69708 170824 69760
rect 558920 69708 558972 69760
rect 33140 69640 33192 69692
rect 127440 69640 127492 69692
rect 169484 69640 169536 69692
rect 564532 69640 564584 69692
rect 137192 68960 137244 69012
rect 138848 68960 138900 69012
rect 138664 68824 138716 68876
rect 171140 68824 171192 68876
rect 141424 68756 141476 68808
rect 202880 68756 202932 68808
rect 157064 68688 157116 68740
rect 249800 68688 249852 68740
rect 18604 68620 18656 68672
rect 183008 68620 183060 68672
rect 150992 68552 151044 68604
rect 332692 68552 332744 68604
rect 159272 68484 159324 68536
rect 431960 68484 432012 68536
rect 115940 68416 115992 68468
rect 134248 68416 134300 68468
rect 163504 68416 163556 68468
rect 481640 68416 481692 68468
rect 85580 68348 85632 68400
rect 132132 68348 132184 68400
rect 167644 68348 167696 68400
rect 543740 68348 543792 68400
rect 59360 68280 59412 68332
rect 129832 68280 129884 68332
rect 170588 68280 170640 68332
rect 550640 68280 550692 68332
rect 139952 67124 140004 67176
rect 189080 67124 189132 67176
rect 141332 67056 141384 67108
rect 207020 67056 207072 67108
rect 153752 66988 153804 67040
rect 356060 66988 356112 67040
rect 64880 66920 64932 66972
rect 130200 66920 130252 66972
rect 155132 66920 155184 66972
rect 374092 66920 374144 66972
rect 16580 66852 16632 66904
rect 126152 66852 126204 66904
rect 166264 66852 166316 66904
rect 525800 66852 525852 66904
rect 138572 66172 138624 66224
rect 140136 66172 140188 66224
rect 148324 65696 148376 65748
rect 292580 65696 292632 65748
rect 156604 65628 156656 65680
rect 390560 65628 390612 65680
rect 158352 65560 158404 65612
rect 396080 65560 396132 65612
rect 170220 65492 170272 65544
rect 568580 65492 568632 65544
rect 120080 64880 120132 64932
rect 123668 64880 123720 64932
rect 145564 64336 145616 64388
rect 256700 64336 256752 64388
rect 157984 64268 158036 64320
rect 412640 64268 412692 64320
rect 160836 64200 160888 64252
rect 444380 64200 444432 64252
rect 169024 64132 169076 64184
rect 561680 64132 561732 64184
rect 148692 62908 148744 62960
rect 190460 62908 190512 62960
rect 157892 62840 157944 62892
rect 408500 62840 408552 62892
rect 159180 62772 159232 62824
rect 440240 62772 440292 62824
rect 145472 61548 145524 61600
rect 259460 61548 259512 61600
rect 155040 61480 155092 61532
rect 380900 61480 380952 61532
rect 163412 61412 163464 61464
rect 481732 61412 481784 61464
rect 118332 61344 118384 61396
rect 580264 61344 580316 61396
rect 138480 60664 138532 60716
rect 144276 60664 144328 60716
rect 182824 60664 182876 60716
rect 580172 60664 580224 60716
rect 139768 60256 139820 60308
rect 179512 60256 179564 60308
rect 139860 60188 139912 60240
rect 183560 60188 183612 60240
rect 148232 60120 148284 60172
rect 295340 60120 295392 60172
rect 154948 60052 155000 60104
rect 376760 60052 376812 60104
rect 102232 59984 102284 60036
rect 125416 59984 125468 60036
rect 161112 59984 161164 60036
rect 390652 59984 390704 60036
rect 3056 59304 3108 59356
rect 18604 59304 18656 59356
rect 137100 59304 137152 59356
rect 140228 59304 140280 59356
rect 139676 58964 139728 59016
rect 180800 58964 180852 59016
rect 150900 58896 150952 58948
rect 327080 58896 327132 58948
rect 153660 58828 153712 58880
rect 358820 58828 358872 58880
rect 159088 58760 159140 58812
rect 433340 58760 433392 58812
rect 164792 58692 164844 58744
rect 507860 58692 507912 58744
rect 170128 58624 170180 58676
rect 572720 58624 572772 58676
rect 141240 57264 141292 57316
rect 201500 57264 201552 57316
rect 156512 57196 156564 57248
rect 394700 57196 394752 57248
rect 150808 55904 150860 55956
rect 331220 55904 331272 55956
rect 95240 55836 95292 55888
rect 125324 55836 125376 55888
rect 154856 55836 154908 55888
rect 383660 55836 383712 55888
rect 142712 54680 142764 54732
rect 219440 54680 219492 54732
rect 152372 54612 152424 54664
rect 349160 54612 349212 54664
rect 153568 54544 153620 54596
rect 362960 54544 363012 54596
rect 156420 54476 156472 54528
rect 398840 54476 398892 54528
rect 139584 53252 139636 53304
rect 185032 53252 185084 53304
rect 160744 53184 160796 53236
rect 455420 53184 455472 53236
rect 163320 53116 163372 53168
rect 488540 53116 488592 53168
rect 166172 53048 166224 53100
rect 516140 53048 516192 53100
rect 135812 52980 135864 53032
rect 140320 52980 140372 53032
rect 141148 51824 141200 51876
rect 204260 51824 204312 51876
rect 153476 51756 153528 51808
rect 365720 51756 365772 51808
rect 157800 51688 157852 51740
rect 415400 51688 415452 51740
rect 154028 50668 154080 50720
rect 353300 50668 353352 50720
rect 156328 50600 156380 50652
rect 401600 50600 401652 50652
rect 160652 50532 160704 50584
rect 448520 50532 448572 50584
rect 167552 50464 167604 50516
rect 534080 50464 534132 50516
rect 167460 50396 167512 50448
rect 542360 50396 542412 50448
rect 168932 50328 168984 50380
rect 557540 50328 557592 50380
rect 145380 49240 145432 49292
rect 259552 49240 259604 49292
rect 156972 49172 157024 49224
rect 389180 49172 389232 49224
rect 171692 49104 171744 49156
rect 425060 49104 425112 49156
rect 164700 49036 164752 49088
rect 498292 49036 498344 49088
rect 168840 48968 168892 49020
rect 552020 48968 552072 49020
rect 142620 47812 142672 47864
rect 215300 47812 215352 47864
rect 158996 47744 159048 47796
rect 436100 47744 436152 47796
rect 160560 47676 160612 47728
rect 451280 47676 451332 47728
rect 163228 47608 163280 47660
rect 484400 47608 484452 47660
rect 45560 47540 45612 47592
rect 120908 47540 120960 47592
rect 138388 47540 138440 47592
rect 153844 47540 153896 47592
rect 170036 47540 170088 47592
rect 571340 47540 571392 47592
rect 118424 46860 118476 46912
rect 580172 46860 580224 46912
rect 137008 46792 137060 46844
rect 138664 46792 138716 46844
rect 141056 46384 141108 46436
rect 208400 46384 208452 46436
rect 144184 46316 144236 46368
rect 233240 46316 233292 46368
rect 156236 46248 156288 46300
rect 391940 46248 391992 46300
rect 138296 46180 138348 46232
rect 156604 46180 156656 46232
rect 163136 46180 163188 46232
rect 491300 46180 491352 46232
rect 3516 45500 3568 45552
rect 173992 45500 174044 45552
rect 142528 45024 142580 45076
rect 218152 45024 218204 45076
rect 148140 44956 148192 45008
rect 289820 44956 289872 45008
rect 171876 44888 171928 44940
rect 397460 44888 397512 44940
rect 81440 44820 81492 44872
rect 131396 44820 131448 44872
rect 168748 44820 168800 44872
rect 553400 44820 553452 44872
rect 148048 43528 148100 43580
rect 285680 43528 285732 43580
rect 171508 43460 171560 43512
rect 432052 43460 432104 43512
rect 88340 43392 88392 43444
rect 125232 43392 125284 43444
rect 169668 43392 169720 43444
rect 563060 43392 563112 43444
rect 139492 42168 139544 42220
rect 187700 42168 187752 42220
rect 157708 42100 157760 42152
rect 415492 42100 415544 42152
rect 169944 42032 169996 42084
rect 572812 42032 572864 42084
rect 152280 40740 152332 40792
rect 345020 40740 345072 40792
rect 169852 40672 169904 40724
rect 569960 40672 570012 40724
rect 153384 39448 153436 39500
rect 357532 39448 357584 39500
rect 157616 39380 157668 39432
rect 409880 39380 409932 39432
rect 166080 39312 166132 39364
rect 527180 39312 527232 39364
rect 157524 37952 157576 38004
rect 419540 37952 419592 38004
rect 164608 37884 164660 37936
rect 503720 37884 503772 37936
rect 31760 36524 31812 36576
rect 122380 36524 122432 36576
rect 27620 35164 27672 35216
rect 127256 35164 127308 35216
rect 163044 35164 163096 35216
rect 487160 35164 487212 35216
rect 2872 33056 2924 33108
rect 21456 33056 21508 33108
rect 147864 32444 147916 32496
rect 291200 32444 291252 32496
rect 147956 32376 148008 32428
rect 293960 32376 294012 32428
rect 140964 31356 141016 31408
rect 205640 31356 205692 31408
rect 142436 31288 142488 31340
rect 216680 31288 216732 31340
rect 144092 31220 144144 31272
rect 237380 31220 237432 31272
rect 164516 31152 164568 31204
rect 499580 31152 499632 31204
rect 167368 31084 167420 31136
rect 535460 31084 535512 31136
rect 169760 31016 169812 31068
rect 574100 31016 574152 31068
rect 150716 29792 150768 29844
rect 324412 29792 324464 29844
rect 152188 29724 152240 29776
rect 339500 29724 339552 29776
rect 153108 29656 153160 29708
rect 346400 29656 346452 29708
rect 158904 29588 158956 29640
rect 427820 29588 427872 29640
rect 150624 28364 150676 28416
rect 321560 28364 321612 28416
rect 153292 28296 153344 28348
rect 360200 28296 360252 28348
rect 172152 28228 172204 28280
rect 418160 28228 418212 28280
rect 145288 26936 145340 26988
rect 258080 26936 258132 26988
rect 154764 26868 154816 26920
rect 378140 26868 378192 26920
rect 144000 25644 144052 25696
rect 236000 25644 236052 25696
rect 145196 25576 145248 25628
rect 251272 25576 251324 25628
rect 154672 25508 154724 25560
rect 385040 25508 385092 25560
rect 142344 24216 142396 24268
rect 222200 24216 222252 24268
rect 147772 24148 147824 24200
rect 292672 24148 292724 24200
rect 106280 24080 106332 24132
rect 132868 24080 132920 24132
rect 165988 24080 166040 24132
rect 524420 24080 524472 24132
rect 139400 22992 139452 23044
rect 186320 22992 186372 23044
rect 150532 22924 150584 22976
rect 328460 22924 328512 22976
rect 67640 22856 67692 22908
rect 130108 22856 130160 22908
rect 157432 22856 157484 22908
rect 416780 22856 416832 22908
rect 60832 22788 60884 22840
rect 129188 22788 129240 22840
rect 165896 22788 165948 22840
rect 521660 22788 521712 22840
rect 3516 22720 3568 22772
rect 179696 22720 179748 22772
rect 184204 22720 184256 22772
rect 580172 22720 580224 22772
rect 135720 21632 135772 21684
rect 139400 21632 139452 21684
rect 138204 21564 138256 21616
rect 168656 21564 168708 21616
rect 154580 21496 154632 21548
rect 379520 21496 379572 21548
rect 136916 21428 136968 21480
rect 147772 21428 147824 21480
rect 172060 21428 172112 21480
rect 404360 21428 404412 21480
rect 38660 21360 38712 21412
rect 120816 21360 120868 21412
rect 168564 21360 168616 21412
rect 556160 21360 556212 21412
rect 143908 20204 143960 20256
rect 241520 20204 241572 20256
rect 145104 20136 145156 20188
rect 262220 20136 262272 20188
rect 152004 20068 152056 20120
rect 343640 20068 343692 20120
rect 124220 20000 124272 20052
rect 134064 20000 134116 20052
rect 145012 20000 145064 20052
rect 255320 20000 255372 20052
rect 255964 20000 256016 20052
rect 456800 20000 456852 20052
rect 99380 19932 99432 19984
rect 132776 19932 132828 19984
rect 156144 19932 156196 19984
rect 400220 19932 400272 19984
rect 140872 18776 140924 18828
rect 198740 18776 198792 18828
rect 158812 18708 158864 18760
rect 429200 18708 429252 18760
rect 168380 18640 168432 18692
rect 556252 18640 556304 18692
rect 168472 18572 168524 18624
rect 560300 18572 560352 18624
rect 160468 17416 160520 17468
rect 445760 17416 445812 17468
rect 160376 17348 160428 17400
rect 452660 17348 452712 17400
rect 162952 17280 163004 17332
rect 492680 17280 492732 17332
rect 167276 17212 167328 17264
rect 540980 17212 541032 17264
rect 151912 16124 151964 16176
rect 342904 16124 342956 16176
rect 160192 16056 160244 16108
rect 448612 16056 448664 16108
rect 160284 15988 160336 16040
rect 454040 15988 454092 16040
rect 165712 15920 165764 15972
rect 517888 15920 517940 15972
rect 165804 15852 165856 15904
rect 523776 15852 523828 15904
rect 144920 14764 144972 14816
rect 254216 14764 254268 14816
rect 149796 14696 149848 14748
rect 305552 14696 305604 14748
rect 149704 14628 149756 14680
rect 307760 14628 307812 14680
rect 124128 14560 124180 14612
rect 312176 14560 312228 14612
rect 315304 14560 315356 14612
rect 475752 14560 475804 14612
rect 156052 14492 156104 14544
rect 398932 14492 398984 14544
rect 165620 14424 165672 14476
rect 520280 14424 520332 14476
rect 15936 13064 15988 13116
rect 113824 13064 113876 13116
rect 140780 12316 140832 12368
rect 202696 12316 202748 12368
rect 147036 12248 147088 12300
rect 273260 12248 273312 12300
rect 146944 12180 146996 12232
rect 276664 12180 276716 12232
rect 147680 12112 147732 12164
rect 287336 12112 287388 12164
rect 149520 12044 149572 12096
rect 311440 12044 311492 12096
rect 149612 11976 149664 12028
rect 314660 11976 314712 12028
rect 160008 11908 160060 11960
rect 435088 11908 435140 11960
rect 160100 11840 160152 11892
rect 447416 11840 447468 11892
rect 140412 11772 140464 11824
rect 156144 11772 156196 11824
rect 162032 11772 162084 11824
rect 463976 11772 464028 11824
rect 136824 11704 136876 11756
rect 153752 11704 153804 11756
rect 161940 11704 161992 11756
rect 470600 11704 470652 11756
rect 173532 11636 173584 11688
rect 173716 11636 173768 11688
rect 110512 10412 110564 10464
rect 125140 10412 125192 10464
rect 25320 10344 25372 10396
rect 106924 10344 106976 10396
rect 117320 10344 117372 10396
rect 134432 10344 134484 10396
rect 44272 10276 44324 10328
rect 128544 10276 128596 10328
rect 138112 10276 138164 10328
rect 166080 10276 166132 10328
rect 146852 9596 146904 9648
rect 272432 9596 272484 9648
rect 146668 9528 146720 9580
rect 276020 9528 276072 9580
rect 149428 9460 149480 9512
rect 304356 9460 304408 9512
rect 149336 9392 149388 9444
rect 307944 9392 307996 9444
rect 171416 9324 171468 9376
rect 411904 9324 411956 9376
rect 157340 9256 157392 9308
rect 414296 9256 414348 9308
rect 161664 9188 161716 9240
rect 466276 9188 466328 9240
rect 161756 9120 161808 9172
rect 469864 9120 469916 9172
rect 34796 9052 34848 9104
rect 127808 9052 127860 9104
rect 161848 9052 161900 9104
rect 473452 9052 473504 9104
rect 24216 8984 24268 9036
rect 122288 8984 122340 9036
rect 164424 8984 164476 9036
rect 510068 8984 510120 9036
rect 9956 8916 10008 8968
rect 125968 8916 126020 8968
rect 167184 8916 167236 8968
rect 539600 8916 539652 8968
rect 146760 8848 146812 8900
rect 268844 8848 268896 8900
rect 105728 7828 105780 7880
rect 132960 7828 133012 7880
rect 98644 7760 98696 7812
rect 133144 7760 133196 7812
rect 27712 7692 27764 7744
rect 127348 7692 127400 7744
rect 23020 7624 23072 7676
rect 127532 7624 127584 7676
rect 150440 7624 150492 7676
rect 330392 7624 330444 7676
rect 18236 7556 18288 7608
rect 125876 7556 125928 7608
rect 164332 7556 164384 7608
rect 506480 7556 506532 7608
rect 146484 6808 146536 6860
rect 278320 6808 278372 6860
rect 149244 6740 149296 6792
rect 310244 6740 310296 6792
rect 149152 6672 149204 6724
rect 313832 6672 313884 6724
rect 172336 6604 172388 6656
rect 342168 6604 342220 6656
rect 151820 6536 151872 6588
rect 338672 6536 338724 6588
rect 84476 6468 84528 6520
rect 131304 6468 131356 6520
rect 153200 6468 153252 6520
rect 364616 6468 364668 6520
rect 80888 6400 80940 6452
rect 131672 6400 131724 6452
rect 155960 6400 156012 6452
rect 394240 6400 394292 6452
rect 78588 6332 78640 6384
rect 129004 6332 129056 6384
rect 161572 6332 161624 6384
rect 462780 6332 462832 6384
rect 70308 6264 70360 6316
rect 130016 6264 130068 6316
rect 161480 6264 161532 6316
rect 467472 6264 467524 6316
rect 63224 6196 63276 6248
rect 130476 6196 130528 6248
rect 164240 6196 164292 6248
rect 502984 6196 503036 6248
rect 538864 6196 538916 6248
rect 581000 6196 581052 6248
rect 13544 6128 13596 6180
rect 126520 6128 126572 6180
rect 167092 6128 167144 6180
rect 545488 6128 545540 6180
rect 146576 6060 146628 6112
rect 274824 6060 274876 6112
rect 146392 5992 146444 6044
rect 270040 5992 270092 6044
rect 85672 5108 85724 5160
rect 131580 5108 131632 5160
rect 66720 5040 66772 5092
rect 130292 5040 130344 5092
rect 52552 4972 52604 5024
rect 128728 4972 128780 5024
rect 138020 4972 138072 5024
rect 167184 4972 167236 5024
rect 6460 4904 6512 4956
rect 17224 4904 17276 4956
rect 48964 4904 49016 4956
rect 128912 4904 128964 4956
rect 143816 4904 143868 4956
rect 234620 4904 234672 4956
rect 8760 4836 8812 4888
rect 126336 4836 126388 4888
rect 137928 4836 137980 4888
rect 151820 4836 151872 4888
rect 162860 4836 162912 4888
rect 486424 4836 486476 4888
rect 5264 4768 5316 4820
rect 126060 4768 126112 4820
rect 136732 4768 136784 4820
rect 157800 4768 157852 4820
rect 168288 4768 168340 4820
rect 538404 4768 538456 4820
rect 138940 4360 138992 4412
rect 143540 4360 143592 4412
rect 125876 4088 125928 4140
rect 134524 4088 134576 4140
rect 142252 4088 142304 4140
rect 221556 4088 221608 4140
rect 143724 4020 143776 4072
rect 235816 4020 235868 4072
rect 144552 3952 144604 4004
rect 239312 3952 239364 4004
rect 117688 3884 117740 3936
rect 122196 3884 122248 3936
rect 143632 3884 143684 3936
rect 242900 3884 242952 3936
rect 251180 3884 251232 3936
rect 252376 3884 252428 3936
rect 259460 3884 259512 3936
rect 260656 3884 260708 3936
rect 77392 3816 77444 3868
rect 123484 3816 123536 3868
rect 128176 3816 128228 3868
rect 131764 3816 131816 3868
rect 140228 3816 140280 3868
rect 144736 3816 144788 3868
rect 146300 3816 146352 3868
rect 271236 3816 271288 3868
rect 284300 3816 284352 3868
rect 285036 3816 285088 3868
rect 299572 3816 299624 3868
rect 300768 3816 300820 3868
rect 64328 3748 64380 3800
rect 126244 3748 126296 3800
rect 138664 3748 138716 3800
rect 145932 3748 145984 3800
rect 149060 3748 149112 3800
rect 306748 3748 306800 3800
rect 47860 3680 47912 3732
rect 123576 3680 123628 3732
rect 131764 3680 131816 3732
rect 135628 3680 135680 3732
rect 142896 3680 142948 3732
rect 155408 3680 155460 3732
rect 156604 3680 156656 3732
rect 168380 3680 168432 3732
rect 173532 3680 173584 3732
rect 178132 3680 178184 3732
rect 184940 3680 184992 3732
rect 186136 3680 186188 3732
rect 186228 3680 186280 3732
rect 468668 3680 468720 3732
rect 43076 3612 43128 3664
rect 125048 3612 125100 3664
rect 133788 3612 133840 3664
rect 147128 3612 147180 3664
rect 155224 3612 155276 3664
rect 160100 3612 160152 3664
rect 160744 3612 160796 3664
rect 173164 3612 173216 3664
rect 173256 3612 173308 3664
rect 461584 3612 461636 3664
rect 2872 3544 2924 3596
rect 117688 3544 117740 3596
rect 119896 3544 119948 3596
rect 122104 3544 122156 3596
rect 135260 3544 135312 3596
rect 136088 3544 136140 3596
rect 140136 3544 140188 3596
rect 572 3476 624 3528
rect 4804 3476 4856 3528
rect 1676 3408 1728 3460
rect 124864 3476 124916 3528
rect 126980 3476 127032 3528
rect 129096 3476 129148 3528
rect 140320 3476 140372 3528
rect 141240 3476 141292 3528
rect 144276 3544 144328 3596
rect 162492 3544 162544 3596
rect 173348 3544 173400 3596
rect 163688 3476 163740 3528
rect 174544 3476 174596 3528
rect 175464 3476 175516 3528
rect 176660 3544 176712 3596
rect 177856 3544 177908 3596
rect 472256 3544 472308 3596
rect 11152 3408 11204 3460
rect 124956 3408 125008 3460
rect 140044 3408 140096 3460
rect 170772 3408 170824 3460
rect 173440 3408 173492 3460
rect 479340 3476 479392 3528
rect 481640 3476 481692 3528
rect 482468 3476 482520 3528
rect 514760 3476 514812 3528
rect 515588 3476 515640 3528
rect 178132 3408 178184 3460
rect 491116 3408 491168 3460
rect 44180 3340 44232 3392
rect 45100 3340 45152 3392
rect 60740 3340 60792 3392
rect 61660 3340 61712 3392
rect 93860 3340 93912 3392
rect 94780 3340 94832 3392
rect 110420 3340 110472 3392
rect 111616 3340 111668 3392
rect 142160 3340 142212 3392
rect 218060 3340 218112 3392
rect 307760 3340 307812 3392
rect 309048 3340 309100 3392
rect 324412 3340 324464 3392
rect 325608 3340 325660 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 349252 3340 349304 3392
rect 350448 3340 350500 3392
rect 357440 3340 357492 3392
rect 358728 3340 358780 3392
rect 365720 3340 365772 3392
rect 367008 3340 367060 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 382280 3340 382332 3392
rect 383568 3340 383620 3392
rect 390560 3340 390612 3392
rect 391848 3340 391900 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 407212 3340 407264 3392
rect 408408 3340 408460 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 138848 3272 138900 3324
rect 150624 3272 150676 3324
rect 138756 3204 138808 3256
rect 149520 3204 149572 3256
rect 172244 3204 172296 3256
rect 200304 3272 200356 3324
rect 181444 3204 181496 3256
rect 186228 3204 186280 3256
rect 118792 3136 118844 3188
rect 120724 3136 120776 3188
rect 129372 3136 129424 3188
rect 134616 3136 134668 3188
rect 135536 3136 135588 3188
rect 137652 3136 137704 3188
rect 144460 3136 144512 3188
rect 153016 3136 153068 3188
rect 172060 3136 172112 3188
rect 182548 3136 182600 3188
rect 135444 3068 135496 3120
rect 138848 3068 138900 3120
rect 153844 3068 153896 3120
rect 161296 3068 161348 3120
rect 432052 2048 432104 2100
rect 433248 2048 433300 2100
rect 415400 1912 415452 1964
rect 416688 1912 416740 1964
rect 440240 1912 440292 1964
rect 441528 1912 441580 1964
rect 456800 1912 456852 1964
rect 458088 1912 458140 1964
<< metal2 >>
rect 6932 703582 7972 703610
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683738 2820 684247
rect 2780 683732 2832 683738
rect 2780 683674 2832 683680
rect 4804 683732 4856 683738
rect 4804 683674 4856 683680
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3332 632120 3384 632126
rect 3330 632088 3332 632097
rect 3384 632088 3386 632097
rect 3330 632023 3386 632032
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579834 3372 579935
rect 3332 579828 3384 579834
rect 3332 579770 3384 579776
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 3238 501800 3294 501809
rect 3238 501735 3294 501744
rect 3252 501022 3280 501735
rect 3240 501016 3292 501022
rect 3240 500958 3292 500964
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3344 462398 3372 462567
rect 3332 462392 3384 462398
rect 3332 462334 3384 462340
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3344 448594 3372 449511
rect 3332 448588 3384 448594
rect 3332 448530 3384 448536
rect 2962 423600 3018 423609
rect 2962 423535 3018 423544
rect 2976 422346 3004 423535
rect 2964 422340 3016 422346
rect 2964 422282 3016 422288
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3344 409902 3372 410479
rect 3332 409896 3384 409902
rect 3332 409838 3384 409844
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3344 357474 3372 358391
rect 3332 357468 3384 357474
rect 3332 357410 3384 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3146 319288 3202 319297
rect 3146 319223 3202 319232
rect 3160 318850 3188 319223
rect 3148 318844 3200 318850
rect 3148 318786 3200 318792
rect 3238 267200 3294 267209
rect 3238 267135 3294 267144
rect 3252 266422 3280 267135
rect 3240 266416 3292 266422
rect 3240 266358 3292 266364
rect 3330 254144 3386 254153
rect 3330 254079 3386 254088
rect 3344 253978 3372 254079
rect 3332 253972 3384 253978
rect 3332 253914 3384 253920
rect 2778 241088 2834 241097
rect 2778 241023 2834 241032
rect 2792 240378 2820 241023
rect 2780 240372 2832 240378
rect 2780 240314 2832 240320
rect 3054 228032 3110 228041
rect 3054 227967 3110 227976
rect 3068 227798 3096 227967
rect 3056 227792 3108 227798
rect 3056 227734 3108 227740
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3344 213994 3372 214911
rect 3332 213988 3384 213994
rect 3332 213930 3384 213936
rect 2962 188864 3018 188873
rect 2962 188799 3018 188808
rect 2976 187746 3004 188799
rect 2964 187740 3016 187746
rect 2964 187682 3016 187688
rect 3332 176112 3384 176118
rect 3332 176054 3384 176060
rect 3344 175953 3372 176054
rect 3330 175944 3386 175953
rect 3330 175879 3386 175888
rect 3332 162920 3384 162926
rect 3330 162888 3332 162897
rect 3384 162888 3386 162897
rect 3330 162823 3386 162832
rect 2964 111784 3016 111790
rect 2964 111726 3016 111732
rect 2976 110673 3004 111726
rect 2962 110664 3018 110673
rect 2962 110599 3018 110608
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 3344 84250 3372 84623
rect 3332 84244 3384 84250
rect 3332 84186 3384 84192
rect 3436 78849 3464 658135
rect 3528 160750 3556 671191
rect 3698 619168 3754 619177
rect 3698 619103 3754 619112
rect 3606 606112 3662 606121
rect 3606 606047 3662 606056
rect 3516 160744 3568 160750
rect 3516 160686 3568 160692
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3528 149122 3556 149767
rect 3516 149116 3568 149122
rect 3516 149058 3568 149064
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3528 136678 3556 136711
rect 3516 136672 3568 136678
rect 3516 136614 3568 136620
rect 3516 135992 3568 135998
rect 3516 135934 3568 135940
rect 3528 97617 3556 135934
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3620 78985 3648 606047
rect 3712 231198 3740 619103
rect 3882 566944 3938 566953
rect 3882 566879 3938 566888
rect 3790 553888 3846 553897
rect 3790 553823 3846 553832
rect 3700 231192 3752 231198
rect 3700 231134 3752 231140
rect 3698 201920 3754 201929
rect 3698 201855 3754 201864
rect 3712 174146 3740 201855
rect 3700 174140 3752 174146
rect 3700 174082 3752 174088
rect 3700 139460 3752 139466
rect 3700 139402 3752 139408
rect 3712 135998 3740 139402
rect 3700 135992 3752 135998
rect 3700 135934 3752 135940
rect 3804 79121 3832 553823
rect 3896 220114 3924 566879
rect 4066 306232 4122 306241
rect 4066 306167 4122 306176
rect 3974 293176 4030 293185
rect 3974 293111 4030 293120
rect 3884 220108 3936 220114
rect 3884 220050 3936 220056
rect 3988 79354 4016 293111
rect 4080 209098 4108 306167
rect 4068 209092 4120 209098
rect 4068 209034 4120 209040
rect 4816 118658 4844 683674
rect 4896 240372 4948 240378
rect 4896 240314 4948 240320
rect 4804 118652 4856 118658
rect 4804 118594 4856 118600
rect 3976 79348 4028 79354
rect 3976 79290 4028 79296
rect 3790 79112 3846 79121
rect 3790 79047 3846 79056
rect 3606 78976 3662 78985
rect 3606 78911 3662 78920
rect 3422 78840 3478 78849
rect 3422 78775 3478 78784
rect 4908 78577 4936 240314
rect 6932 79257 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 7564 632120 7616 632126
rect 7564 632062 7616 632068
rect 7576 120086 7604 632062
rect 8944 579828 8996 579834
rect 8944 579770 8996 579776
rect 8956 121446 8984 579770
rect 10324 527196 10376 527202
rect 10324 527138 10376 527144
rect 9588 180124 9640 180130
rect 9588 180066 9640 180072
rect 9600 176118 9628 180066
rect 9588 176112 9640 176118
rect 9588 176054 9640 176060
rect 10336 122806 10364 527138
rect 18604 474768 18656 474774
rect 18604 474710 18656 474716
rect 13084 422340 13136 422346
rect 13084 422282 13136 422288
rect 13096 126954 13124 422282
rect 14464 371272 14516 371278
rect 14464 371214 14516 371220
rect 14476 128314 14504 371214
rect 17224 318844 17276 318850
rect 17224 318786 17276 318792
rect 17236 129742 17264 318786
rect 17224 129736 17276 129742
rect 17224 129678 17276 129684
rect 14464 128308 14516 128314
rect 14464 128250 14516 128256
rect 13084 126948 13136 126954
rect 13084 126890 13136 126896
rect 18616 124166 18644 474710
rect 21364 266416 21416 266422
rect 21364 266358 21416 266364
rect 18696 133952 18748 133958
rect 18696 133894 18748 133900
rect 18604 124160 18656 124166
rect 18604 124102 18656 124108
rect 10324 122800 10376 122806
rect 10324 122742 10376 122748
rect 8944 121440 8996 121446
rect 8944 121382 8996 121388
rect 7564 120080 7616 120086
rect 7564 120022 7616 120028
rect 18708 111790 18736 133894
rect 21376 131102 21404 266358
rect 22744 213988 22796 213994
rect 22744 213930 22796 213936
rect 21456 136740 21508 136746
rect 21456 136682 21508 136688
rect 21364 131096 21416 131102
rect 21364 131038 21416 131044
rect 18696 111784 18748 111790
rect 18696 111726 18748 111732
rect 6918 79248 6974 79257
rect 6918 79183 6974 79192
rect 4894 78568 4950 78577
rect 4894 78503 4950 78512
rect 17222 77888 17278 77897
rect 17222 77823 17278 77832
rect 6920 75200 6972 75206
rect 6920 75142 6972 75148
rect 4804 73840 4856 73846
rect 4804 73782 4856 73788
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3424 70100 3476 70106
rect 3424 70042 3476 70048
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 2778 21312 2834 21321
rect 2778 21247 2834 21256
rect 2792 16574 2820 21247
rect 2792 16546 3372 16574
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 584 480 612 3470
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1688 480 1716 3402
rect 2884 480 2912 3538
rect 3344 490 3372 16546
rect 3436 6497 3464 70042
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 3528 19417 3556 22714
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4816 3534 4844 73782
rect 6932 16574 6960 75142
rect 13820 72548 13872 72554
rect 13820 72490 13872 72496
rect 11060 72480 11112 72486
rect 11060 72422 11112 72428
rect 11072 16574 11100 72422
rect 13832 16574 13860 72490
rect 16580 66904 16632 66910
rect 16580 66846 16632 66852
rect 16592 16574 16620 66846
rect 6932 16546 7696 16574
rect 11072 16546 11928 16574
rect 13832 16546 14320 16574
rect 16592 16546 17080 16574
rect 6460 4956 6512 4962
rect 6460 4898 6512 4904
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3344 462 3648 490
rect 5276 480 5304 4762
rect 6472 480 6500 4898
rect 7668 480 7696 16546
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 8760 4888 8812 4894
rect 8760 4830 8812 4836
rect 8772 480 8800 4830
rect 9968 480 9996 8910
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 480 11192 3402
rect 3620 354 3648 462
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 11900 354 11928 16546
rect 13544 6180 13596 6186
rect 13544 6122 13596 6128
rect 13556 480 13584 6122
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15936 13116 15988 13122
rect 15936 13058 15988 13064
rect 15948 480 15976 13058
rect 17052 480 17080 16546
rect 17236 4962 17264 77823
rect 20718 76528 20774 76537
rect 20718 76463 20774 76472
rect 18604 68672 18656 68678
rect 18604 68614 18656 68620
rect 18616 59362 18644 68614
rect 18604 59356 18656 59362
rect 18604 59298 18656 59304
rect 19338 35184 19394 35193
rect 19338 35119 19394 35128
rect 19352 16574 19380 35119
rect 20732 16574 20760 76463
rect 21468 33114 21496 136682
rect 22756 132462 22784 213930
rect 23492 159390 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 25504 514820 25556 514826
rect 25504 514762 25556 514768
rect 23480 159384 23532 159390
rect 23480 159326 23532 159332
rect 25516 140078 25544 514762
rect 28264 462392 28316 462398
rect 28264 462334 28316 462340
rect 26884 357468 26936 357474
rect 26884 357410 26936 357416
rect 26896 164898 26924 357410
rect 26884 164892 26936 164898
rect 26884 164834 26936 164840
rect 28276 141506 28304 462334
rect 37924 448588 37976 448594
rect 37924 448530 37976 448536
rect 32404 409896 32456 409902
rect 32404 409838 32456 409844
rect 32416 162178 32444 409838
rect 35164 253972 35216 253978
rect 35164 253914 35216 253920
rect 35176 169046 35204 253914
rect 35164 169040 35216 169046
rect 35164 168982 35216 168988
rect 32404 162172 32456 162178
rect 32404 162114 32456 162120
rect 28264 141500 28316 141506
rect 28264 141442 28316 141448
rect 25504 140072 25556 140078
rect 25504 140014 25556 140020
rect 22744 132456 22796 132462
rect 22744 132398 22796 132404
rect 37936 79393 37964 448530
rect 39304 397520 39356 397526
rect 39304 397462 39356 397468
rect 39316 79626 39344 397462
rect 40052 117298 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 43444 501016 43496 501022
rect 43444 500958 43496 500964
rect 40040 117292 40092 117298
rect 40040 117234 40092 117240
rect 39304 79620 39356 79626
rect 39304 79562 39356 79568
rect 43456 79529 43484 500958
rect 65524 484424 65576 484430
rect 65524 484366 65576 484372
rect 65536 452674 65564 484366
rect 62120 452668 62172 452674
rect 62120 452610 62172 452616
rect 65524 452668 65576 452674
rect 65524 452610 65576 452616
rect 62132 449206 62160 452610
rect 49608 449200 49660 449206
rect 49608 449142 49660 449148
rect 62120 449200 62172 449206
rect 62120 449142 62172 449148
rect 49620 446418 49648 449142
rect 45008 446412 45060 446418
rect 45008 446354 45060 446360
rect 49608 446412 49660 446418
rect 49608 446354 49660 446360
rect 43536 345092 43588 345098
rect 43536 345034 43588 345040
rect 43548 79762 43576 345034
rect 44916 240916 44968 240922
rect 44916 240858 44968 240864
rect 44824 238876 44876 238882
rect 44824 238818 44876 238824
rect 44836 227254 44864 238818
rect 44824 227248 44876 227254
rect 44824 227190 44876 227196
rect 43536 79756 43588 79762
rect 43536 79698 43588 79704
rect 43442 79520 43498 79529
rect 43442 79455 43498 79464
rect 37922 79384 37978 79393
rect 37922 79319 37978 79328
rect 44180 76628 44232 76634
rect 44180 76570 44232 76576
rect 30380 76560 30432 76566
rect 30380 76502 30432 76508
rect 26240 72616 26292 72622
rect 26240 72558 26292 72564
rect 21456 33108 21508 33114
rect 21456 33050 21508 33056
rect 19352 16546 20208 16574
rect 20732 16546 21864 16574
rect 18236 7608 18288 7614
rect 18236 7550 18288 7556
rect 19430 7576 19486 7585
rect 17224 4956 17276 4962
rect 17224 4898 17276 4904
rect 18248 480 18276 7550
rect 19430 7511 19486 7520
rect 19444 480 19472 7511
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20180 354 20208 16546
rect 21836 480 21864 16546
rect 25320 10396 25372 10402
rect 25320 10338 25372 10344
rect 24216 9036 24268 9042
rect 24216 8978 24268 8984
rect 23020 7676 23072 7682
rect 23020 7618 23072 7624
rect 23032 480 23060 7618
rect 24228 480 24256 8978
rect 25332 480 25360 10338
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 72558
rect 29000 71052 29052 71058
rect 29000 70994 29052 71000
rect 27620 35216 27672 35222
rect 27620 35158 27672 35164
rect 27632 16574 27660 35158
rect 29012 16574 29040 70994
rect 30392 16574 30420 76502
rect 35900 75268 35952 75274
rect 35900 75210 35952 75216
rect 33140 69692 33192 69698
rect 33140 69634 33192 69640
rect 31760 36576 31812 36582
rect 31760 36518 31812 36524
rect 31772 16574 31800 36518
rect 33152 16574 33180 69634
rect 27632 16546 28488 16574
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 27712 7744 27764 7750
rect 27712 7686 27764 7692
rect 27724 480 27752 7686
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 30116 480 30144 16546
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33612 480 33640 16546
rect 34796 9104 34848 9110
rect 34796 9046 34848 9052
rect 34808 480 34836 9046
rect 35912 6914 35940 75210
rect 37278 74216 37334 74225
rect 37278 74151 37334 74160
rect 35990 71088 36046 71097
rect 35990 71023 36046 71032
rect 36004 16574 36032 71023
rect 37292 16574 37320 74151
rect 40038 71224 40094 71233
rect 40038 71159 40094 71168
rect 38660 21412 38712 21418
rect 38660 21354 38712 21360
rect 38672 16574 38700 21354
rect 40052 16574 40080 71159
rect 36004 16546 36768 16574
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 35912 6886 36032 6914
rect 36004 480 36032 6886
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41878 8936 41934 8945
rect 41878 8871 41934 8880
rect 41892 480 41920 8871
rect 43076 3664 43128 3670
rect 43076 3606 43128 3612
rect 43088 480 43116 3606
rect 44192 3398 44220 76570
rect 44928 75886 44956 240858
rect 45020 224942 45048 446354
rect 69664 396772 69716 396778
rect 69664 396714 69716 396720
rect 69676 385014 69704 396714
rect 68284 385008 68336 385014
rect 68284 384950 68336 384956
rect 69664 385008 69716 385014
rect 69664 384950 69716 384956
rect 68296 358834 68324 384950
rect 71044 369912 71096 369918
rect 71044 369854 71096 369860
rect 71056 362982 71084 369854
rect 69664 362976 69716 362982
rect 69664 362918 69716 362924
rect 71044 362976 71096 362982
rect 71044 362918 71096 362924
rect 65432 358828 65484 358834
rect 65432 358770 65484 358776
rect 68284 358828 68336 358834
rect 68284 358770 68336 358776
rect 65444 358154 65472 358770
rect 64144 358148 64196 358154
rect 64144 358090 64196 358096
rect 65432 358148 65484 358154
rect 65432 358090 65484 358096
rect 64156 318918 64184 358090
rect 69676 343670 69704 362918
rect 66260 343664 66312 343670
rect 66260 343606 66312 343612
rect 69664 343664 69716 343670
rect 69664 343606 69716 343612
rect 66272 338178 66300 343606
rect 66180 338150 66300 338178
rect 66180 336802 66208 338150
rect 64236 336796 64288 336802
rect 64236 336738 64288 336744
rect 66168 336796 66220 336802
rect 66168 336738 66220 336744
rect 62764 318912 62816 318918
rect 62764 318854 62816 318860
rect 64144 318912 64196 318918
rect 64144 318854 64196 318860
rect 61384 303680 61436 303686
rect 61384 303622 61436 303628
rect 61396 297770 61424 303622
rect 62776 299470 62804 318854
rect 64248 303686 64276 336738
rect 68284 320884 68336 320890
rect 68284 320826 68336 320832
rect 64236 303680 64288 303686
rect 64236 303622 64288 303628
rect 61476 299464 61528 299470
rect 61476 299406 61528 299412
rect 62764 299464 62816 299470
rect 62764 299406 62816 299412
rect 60096 297764 60148 297770
rect 60096 297706 60148 297712
rect 61384 297764 61436 297770
rect 61384 297706 61436 297712
rect 60004 294024 60056 294030
rect 60004 293966 60056 293972
rect 58624 290556 58676 290562
rect 58624 290498 58676 290504
rect 50528 286340 50580 286346
rect 50528 286282 50580 286288
rect 50540 279274 50568 286282
rect 58636 285734 58664 290498
rect 56600 285728 56652 285734
rect 56600 285670 56652 285676
rect 58624 285728 58676 285734
rect 58624 285670 58676 285676
rect 56612 282130 56640 285670
rect 60016 282946 60044 293966
rect 60108 290562 60136 297706
rect 61488 294030 61516 299406
rect 61476 294024 61528 294030
rect 61476 293966 61528 293972
rect 68296 292602 68324 320826
rect 65616 292596 65668 292602
rect 65616 292538 65668 292544
rect 68284 292596 68336 292602
rect 68284 292538 68336 292544
rect 60096 290556 60148 290562
rect 60096 290498 60148 290504
rect 65524 290488 65576 290494
rect 65524 290430 65576 290436
rect 57980 282940 58032 282946
rect 57980 282882 58032 282888
rect 60004 282940 60056 282946
rect 60004 282882 60056 282888
rect 55864 282124 55916 282130
rect 55864 282066 55916 282072
rect 56600 282124 56652 282130
rect 56600 282066 56652 282072
rect 45836 279268 45888 279274
rect 45836 279210 45888 279216
rect 50528 279268 50580 279274
rect 50528 279210 50580 279216
rect 45192 264172 45244 264178
rect 45192 264114 45244 264120
rect 45100 238808 45152 238814
rect 45100 238750 45152 238756
rect 45112 229770 45140 238750
rect 45204 233238 45232 264114
rect 45848 248414 45876 279210
rect 54484 278792 54536 278798
rect 54484 278734 54536 278740
rect 53840 275324 53892 275330
rect 53840 275266 53892 275272
rect 53852 271930 53880 275266
rect 50988 271924 51040 271930
rect 50988 271866 51040 271872
rect 53840 271924 53892 271930
rect 53840 271866 53892 271872
rect 51000 268122 51028 271866
rect 46940 268116 46992 268122
rect 46940 268058 46992 268064
rect 50988 268116 51040 268122
rect 50988 268058 51040 268064
rect 46952 267734 46980 268058
rect 46860 267706 46980 267734
rect 46860 264178 46888 267706
rect 54496 266422 54524 278734
rect 55876 275330 55904 282066
rect 57992 280242 58020 282882
rect 57900 280214 58020 280242
rect 57900 278798 57928 280214
rect 57888 278792 57940 278798
rect 57888 278734 57940 278740
rect 62764 278044 62816 278050
rect 62764 277986 62816 277992
rect 55864 275324 55916 275330
rect 55864 275266 55916 275272
rect 58532 268660 58584 268666
rect 58532 268602 58584 268608
rect 58544 266422 58572 268602
rect 53104 266416 53156 266422
rect 53104 266358 53156 266364
rect 54484 266416 54536 266422
rect 54484 266358 54536 266364
rect 56140 266416 56192 266422
rect 56140 266358 56192 266364
rect 58532 266416 58584 266422
rect 58532 266358 58584 266364
rect 46848 264172 46900 264178
rect 46848 264114 46900 264120
rect 53116 253978 53144 266358
rect 56152 262818 56180 266358
rect 62776 262818 62804 277986
rect 65536 276078 65564 290430
rect 65628 286346 65656 292538
rect 65616 286340 65668 286346
rect 65616 286282 65668 286288
rect 63500 276072 63552 276078
rect 63500 276014 63552 276020
rect 65524 276072 65576 276078
rect 65524 276014 65576 276020
rect 63512 270586 63540 276014
rect 63420 270558 63540 270586
rect 63420 268666 63448 270558
rect 63408 268660 63460 268666
rect 63408 268602 63460 268608
rect 54484 262812 54536 262818
rect 54484 262754 54536 262760
rect 56140 262812 56192 262818
rect 56140 262754 56192 262760
rect 60004 262812 60056 262818
rect 60004 262754 60056 262760
rect 62764 262812 62816 262818
rect 62764 262754 62816 262760
rect 49608 253972 49660 253978
rect 49608 253914 49660 253920
rect 53104 253972 53156 253978
rect 53104 253914 53156 253920
rect 49620 249354 49648 253914
rect 54496 251258 54524 262754
rect 60016 255338 60044 262754
rect 57612 255332 57664 255338
rect 57612 255274 57664 255280
rect 60004 255332 60056 255338
rect 60004 255274 60056 255280
rect 54484 251252 54536 251258
rect 54484 251194 54536 251200
rect 50252 251184 50304 251190
rect 50252 251126 50304 251132
rect 46204 249348 46256 249354
rect 46204 249290 46256 249296
rect 49608 249348 49660 249354
rect 49608 249290 49660 249296
rect 45756 248386 45876 248414
rect 45376 244928 45428 244934
rect 45376 244870 45428 244876
rect 45284 240848 45336 240854
rect 45284 240790 45336 240796
rect 45192 233232 45244 233238
rect 45192 233174 45244 233180
rect 45100 229764 45152 229770
rect 45100 229706 45152 229712
rect 45008 224936 45060 224942
rect 45008 224878 45060 224884
rect 45296 141574 45324 240790
rect 45388 231062 45416 244870
rect 45652 240644 45704 240650
rect 45652 240586 45704 240592
rect 45468 240236 45520 240242
rect 45468 240178 45520 240184
rect 45480 232966 45508 240178
rect 45560 239420 45612 239426
rect 45560 239362 45612 239368
rect 45468 232960 45520 232966
rect 45468 232902 45520 232908
rect 45376 231056 45428 231062
rect 45376 230998 45428 231004
rect 45572 230518 45600 239362
rect 45560 230512 45612 230518
rect 45560 230454 45612 230460
rect 45664 205222 45692 240586
rect 45756 238882 45784 248386
rect 45836 240780 45888 240786
rect 45836 240722 45888 240728
rect 45744 238876 45796 238882
rect 45744 238818 45796 238824
rect 45848 238814 45876 240722
rect 46216 240242 46244 249290
rect 50264 243234 50292 251126
rect 57624 248470 57652 255274
rect 57612 248464 57664 248470
rect 57612 248406 57664 248412
rect 51080 248396 51132 248402
rect 51080 248338 51132 248344
rect 51092 245698 51120 248338
rect 51000 245670 51120 245698
rect 51000 244934 51028 245670
rect 50988 244928 51040 244934
rect 50988 244870 51040 244876
rect 47492 243228 47544 243234
rect 47492 243170 47544 243176
rect 50252 243228 50304 243234
rect 50252 243170 50304 243176
rect 47504 240650 47532 243170
rect 71792 240922 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 79324 592680 79376 592686
rect 79324 592622 79376 592628
rect 79336 487830 79364 592622
rect 73160 487824 73212 487830
rect 73160 487766 73212 487772
rect 79324 487824 79376 487830
rect 79324 487766 79376 487772
rect 73172 484430 73200 487766
rect 73160 484424 73212 484430
rect 73160 484366 73212 484372
rect 87696 408468 87748 408474
rect 87696 408410 87748 408416
rect 87708 405754 87736 408410
rect 87696 405748 87748 405754
rect 87696 405690 87748 405696
rect 84200 405680 84252 405686
rect 84200 405622 84252 405628
rect 84212 401674 84240 405622
rect 84200 401668 84252 401674
rect 84200 401610 84252 401616
rect 82452 401600 82504 401606
rect 82452 401542 82504 401548
rect 82464 397526 82492 401542
rect 80704 397520 80756 397526
rect 80704 397462 80756 397468
rect 82452 397520 82504 397526
rect 82452 397462 82504 397468
rect 80716 388482 80744 397462
rect 73804 388476 73856 388482
rect 73804 388418 73856 388424
rect 80704 388476 80756 388482
rect 80704 388418 80756 388424
rect 73816 369918 73844 388418
rect 73804 369912 73856 369918
rect 73804 369854 73856 369860
rect 79324 331900 79376 331906
rect 79324 331842 79376 331848
rect 79336 320890 79364 331842
rect 79324 320884 79376 320890
rect 79324 320826 79376 320832
rect 80060 244928 80112 244934
rect 80060 244870 80112 244876
rect 71780 240916 71832 240922
rect 71780 240858 71832 240864
rect 47492 240644 47544 240650
rect 47492 240586 47544 240592
rect 46204 240236 46256 240242
rect 46204 240178 46256 240184
rect 80072 239834 80100 244870
rect 88352 240854 88380 702406
rect 104164 551540 104216 551546
rect 104164 551482 104216 551488
rect 104176 527202 104204 551482
rect 101404 527196 101456 527202
rect 101404 527138 101456 527144
rect 104164 527196 104216 527202
rect 104164 527138 104216 527144
rect 101416 516186 101444 527138
rect 98644 516180 98696 516186
rect 98644 516122 98696 516128
rect 101404 516180 101456 516186
rect 101404 516122 101456 516128
rect 98656 473074 98684 516122
rect 97264 473068 97316 473074
rect 97264 473010 97316 473016
rect 98644 473068 98696 473074
rect 98644 473010 98696 473016
rect 97276 469266 97304 473010
rect 95884 469260 95936 469266
rect 95884 469202 95936 469208
rect 97264 469260 97316 469266
rect 97264 469202 97316 469208
rect 95896 445738 95924 469202
rect 94504 445732 94556 445738
rect 94504 445674 94556 445680
rect 95884 445732 95936 445738
rect 95884 445674 95936 445680
rect 94516 422346 94544 445674
rect 93124 422340 93176 422346
rect 93124 422282 93176 422288
rect 94504 422340 94556 422346
rect 94504 422282 94556 422288
rect 93136 413982 93164 422282
rect 91100 413976 91152 413982
rect 91100 413918 91152 413924
rect 93124 413976 93176 413982
rect 93124 413918 93176 413924
rect 91112 408542 91140 413918
rect 91100 408536 91152 408542
rect 91100 408478 91152 408484
rect 102784 305652 102836 305658
rect 102784 305594 102836 305600
rect 102796 290426 102824 305594
rect 104912 290494 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 135904 644428 135956 644434
rect 135904 644370 135956 644376
rect 133144 639600 133196 639606
rect 133144 639542 133196 639548
rect 129740 623824 129792 623830
rect 129740 623766 129792 623772
rect 113824 623076 113876 623082
rect 113824 623018 113876 623024
rect 113836 611998 113864 623018
rect 129752 621042 129780 623766
rect 133156 623082 133184 639542
rect 135916 630698 135944 644370
rect 133236 630692 133288 630698
rect 133236 630634 133288 630640
rect 135904 630692 135956 630698
rect 135904 630634 135956 630640
rect 133248 623830 133276 630634
rect 133236 623824 133288 623830
rect 133236 623766 133288 623772
rect 133144 623076 133196 623082
rect 133144 623018 133196 623024
rect 129004 621036 129056 621042
rect 129004 620978 129056 620984
rect 129740 621036 129792 621042
rect 129740 620978 129792 620984
rect 108304 611992 108356 611998
rect 108304 611934 108356 611940
rect 113824 611992 113876 611998
rect 113824 611934 113876 611940
rect 108316 592686 108344 611934
rect 108304 592680 108356 592686
rect 108304 592622 108356 592628
rect 109684 576156 109736 576162
rect 109684 576098 109736 576104
rect 109696 561066 109724 576098
rect 108304 561060 108356 561066
rect 108304 561002 108356 561008
rect 109684 561060 109736 561066
rect 109684 561002 109736 561008
rect 108316 556238 108344 561002
rect 106280 556232 106332 556238
rect 106280 556174 106332 556180
rect 108304 556232 108356 556238
rect 108304 556174 108356 556180
rect 106292 551546 106320 556174
rect 106280 551540 106332 551546
rect 106280 551482 106332 551488
rect 129016 540938 129044 620978
rect 127624 540932 127676 540938
rect 127624 540874 127676 540880
rect 129004 540932 129056 540938
rect 129004 540874 129056 540880
rect 127636 529922 127664 540874
rect 126244 529916 126296 529922
rect 126244 529858 126296 529864
rect 127624 529916 127676 529922
rect 127624 529858 127676 529864
rect 126256 520266 126284 529858
rect 124220 520260 124272 520266
rect 124220 520202 124272 520208
rect 126244 520260 126296 520266
rect 126244 520202 126296 520208
rect 124232 514826 124260 520202
rect 123484 514820 123536 514826
rect 123484 514762 123536 514768
rect 124220 514820 124272 514826
rect 124220 514762 124272 514768
rect 123496 420238 123524 514762
rect 122104 420232 122156 420238
rect 122104 420174 122156 420180
rect 123484 420232 123536 420238
rect 123484 420174 123536 420180
rect 122116 401674 122144 420174
rect 131764 402280 131816 402286
rect 131764 402222 131816 402228
rect 119344 401668 119396 401674
rect 119344 401610 119396 401616
rect 122104 401668 122156 401674
rect 122104 401610 122156 401616
rect 119356 398886 119384 401610
rect 116584 398880 116636 398886
rect 116584 398822 116636 398828
rect 119344 398880 119396 398886
rect 119344 398822 119396 398828
rect 116596 370802 116624 398822
rect 114928 370796 114980 370802
rect 114928 370738 114980 370744
rect 116584 370796 116636 370802
rect 116584 370738 116636 370744
rect 114940 367810 114968 370738
rect 112444 367804 112496 367810
rect 112444 367746 112496 367752
rect 114928 367804 114980 367810
rect 114928 367746 114980 367752
rect 112456 353326 112484 367746
rect 131776 357066 131804 402222
rect 136652 396778 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 153212 678094 153240 702406
rect 169772 695450 169800 702406
rect 169680 695422 169800 695450
rect 169680 692102 169708 695422
rect 201512 694822 201540 702986
rect 182180 694816 182232 694822
rect 182180 694758 182232 694764
rect 201500 694816 201552 694822
rect 201500 694758 201552 694764
rect 160744 692096 160796 692102
rect 160744 692038 160796 692044
rect 169668 692096 169720 692102
rect 169668 692038 169720 692044
rect 147772 678088 147824 678094
rect 147772 678030 147824 678036
rect 153200 678088 153252 678094
rect 153200 678030 153252 678036
rect 147784 675578 147812 678030
rect 147036 675572 147088 675578
rect 147036 675514 147088 675520
rect 147772 675572 147824 675578
rect 147772 675514 147824 675520
rect 147048 667894 147076 675514
rect 160756 674830 160784 692038
rect 182192 690266 182220 694758
rect 180064 690260 180116 690266
rect 180064 690202 180116 690208
rect 182180 690260 182232 690266
rect 182180 690202 182232 690208
rect 159456 674824 159508 674830
rect 159456 674766 159508 674772
rect 160744 674824 160796 674830
rect 160744 674766 160796 674772
rect 159468 668642 159496 674766
rect 157340 668636 157392 668642
rect 157340 668578 157392 668584
rect 159456 668636 159508 668642
rect 159456 668578 159508 668584
rect 145564 667888 145616 667894
rect 145564 667830 145616 667836
rect 147036 667888 147088 667894
rect 147036 667830 147088 667836
rect 145576 658034 145604 667830
rect 157352 665854 157380 668578
rect 150440 665848 150492 665854
rect 150440 665790 150492 665796
rect 157340 665848 157392 665854
rect 157340 665790 157392 665796
rect 150452 662454 150480 665790
rect 180076 662454 180104 690202
rect 146944 662448 146996 662454
rect 146944 662390 146996 662396
rect 150440 662448 150492 662454
rect 150440 662390 150492 662396
rect 173164 662448 173216 662454
rect 173164 662390 173216 662396
rect 180064 662448 180116 662454
rect 180064 662390 180116 662396
rect 142804 658028 142856 658034
rect 142804 657970 142856 657976
rect 145564 658028 145616 658034
rect 145564 657970 145616 657976
rect 142816 652798 142844 657970
rect 142804 652792 142856 652798
rect 142804 652734 142856 652740
rect 138388 652724 138440 652730
rect 138388 652666 138440 652672
rect 138400 644502 138428 652666
rect 138388 644496 138440 644502
rect 138388 644438 138440 644444
rect 146956 618934 146984 662390
rect 173176 652798 173204 662390
rect 218072 658238 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 235184 697610 235212 703520
rect 267660 697610 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 233884 697604 233936 697610
rect 233884 697546 233936 697552
rect 235172 697604 235224 697610
rect 235172 697546 235224 697552
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 233896 684554 233924 697546
rect 233884 684548 233936 684554
rect 233884 684490 233936 684496
rect 230848 684480 230900 684486
rect 230848 684422 230900 684428
rect 230860 681766 230888 684422
rect 229744 681760 229796 681766
rect 229744 681702 229796 681708
rect 230848 681760 230900 681766
rect 230848 681702 230900 681708
rect 229756 663814 229784 681702
rect 266372 674150 266400 697546
rect 279424 687540 279476 687546
rect 279424 687482 279476 687488
rect 279436 674898 279464 687482
rect 272524 674892 272576 674898
rect 272524 674834 272576 674840
rect 279424 674892 279476 674898
rect 279424 674834 279476 674840
rect 266360 674144 266412 674150
rect 266360 674086 266412 674092
rect 228364 663808 228416 663814
rect 228364 663750 228416 663756
rect 229744 663808 229796 663814
rect 229744 663750 229796 663756
rect 215944 658232 215996 658238
rect 215944 658174 215996 658180
rect 218060 658232 218112 658238
rect 218060 658174 218112 658180
rect 167000 652792 167052 652798
rect 167000 652734 167052 652740
rect 173164 652792 173216 652798
rect 173164 652734 173216 652740
rect 167012 650078 167040 652734
rect 215956 650078 215984 658174
rect 228376 652798 228404 663750
rect 272536 658986 272564 674834
rect 275284 674144 275336 674150
rect 275284 674086 275336 674092
rect 275296 661910 275324 674086
rect 275284 661904 275336 661910
rect 275284 661846 275336 661852
rect 278044 661904 278096 661910
rect 278044 661846 278096 661852
rect 260104 658980 260156 658986
rect 260104 658922 260156 658928
rect 272524 658980 272576 658986
rect 272524 658922 272576 658928
rect 222844 652792 222896 652798
rect 222844 652734 222896 652740
rect 228364 652792 228416 652798
rect 228364 652734 228416 652740
rect 165344 650072 165396 650078
rect 165344 650014 165396 650020
rect 167000 650072 167052 650078
rect 167000 650014 167052 650020
rect 213184 650072 213236 650078
rect 213184 650014 213236 650020
rect 215944 650072 215996 650078
rect 215944 650014 215996 650020
rect 165356 646542 165384 650014
rect 159364 646536 159416 646542
rect 159364 646478 159416 646484
rect 165344 646536 165396 646542
rect 165344 646478 165396 646484
rect 159376 639606 159404 646478
rect 159364 639600 159416 639606
rect 159364 639542 159416 639548
rect 213196 638654 213224 650014
rect 222856 640354 222884 652734
rect 221556 640348 221608 640354
rect 221556 640290 221608 640296
rect 222844 640348 222896 640354
rect 222844 640290 222896 640296
rect 210424 638648 210476 638654
rect 210424 638590 210476 638596
rect 213184 638648 213236 638654
rect 213184 638590 213236 638596
rect 145564 618928 145616 618934
rect 145564 618870 145616 618876
rect 146944 618928 146996 618934
rect 146944 618870 146996 618876
rect 145576 608530 145604 618870
rect 143540 608524 143592 608530
rect 143540 608466 143592 608472
rect 145564 608524 145616 608530
rect 145564 608466 145616 608472
rect 143552 604518 143580 608466
rect 142804 604512 142856 604518
rect 142804 604454 142856 604460
rect 143540 604512 143592 604518
rect 143540 604454 143592 604460
rect 142816 586566 142844 604454
rect 141424 586560 141476 586566
rect 141424 586502 141476 586508
rect 142804 586560 142856 586566
rect 142804 586502 142856 586508
rect 141436 576162 141464 586502
rect 141424 576156 141476 576162
rect 141424 576098 141476 576104
rect 210436 573306 210464 638590
rect 221568 638450 221596 640290
rect 220084 638444 220136 638450
rect 220084 638386 220136 638392
rect 221556 638444 221608 638450
rect 221556 638386 221608 638392
rect 220096 580990 220124 638386
rect 260116 626618 260144 658922
rect 278056 652118 278084 661846
rect 282932 653750 282960 702406
rect 300136 700330 300164 703520
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 292580 700324 292632 700330
rect 292580 700266 292632 700272
rect 300124 700324 300176 700330
rect 300124 700266 300176 700272
rect 292592 697610 292620 700266
rect 284944 697604 284996 697610
rect 284944 697546 284996 697552
rect 292580 697604 292632 697610
rect 292580 697546 292632 697552
rect 284956 687546 284984 697546
rect 284944 687540 284996 687546
rect 284944 687482 284996 687488
rect 331232 655790 331260 702986
rect 348804 700330 348832 703520
rect 364996 700398 365024 703520
rect 364984 700392 365036 700398
rect 364984 700334 365036 700340
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 396632 700324 396684 700330
rect 396632 700266 396684 700272
rect 331220 655784 331272 655790
rect 331220 655726 331272 655732
rect 335360 655784 335412 655790
rect 335360 655726 335412 655732
rect 282920 653744 282972 653750
rect 282920 653686 282972 653692
rect 286324 653744 286376 653750
rect 286324 653686 286376 653692
rect 278044 652112 278096 652118
rect 278044 652054 278096 652060
rect 281448 652112 281500 652118
rect 281448 652054 281500 652060
rect 281460 647222 281488 652054
rect 281448 647216 281500 647222
rect 281448 647158 281500 647164
rect 285680 647216 285732 647222
rect 285680 647158 285732 647164
rect 285692 642462 285720 647158
rect 285680 642456 285732 642462
rect 285680 642398 285732 642404
rect 286336 642394 286364 653686
rect 335372 652798 335400 655726
rect 335360 652792 335412 652798
rect 335360 652734 335412 652740
rect 341524 652792 341576 652798
rect 341524 652734 341576 652740
rect 289084 642456 289136 642462
rect 289084 642398 289136 642404
rect 286324 642388 286376 642394
rect 286324 642330 286376 642336
rect 289096 630222 289124 642398
rect 294604 642388 294656 642394
rect 294604 642330 294656 642336
rect 289084 630216 289136 630222
rect 289084 630158 289136 630164
rect 254584 626612 254636 626618
rect 254584 626554 254636 626560
rect 260104 626612 260156 626618
rect 260104 626554 260156 626560
rect 254596 587246 254624 626554
rect 294616 607918 294644 642330
rect 295340 630216 295392 630222
rect 295340 630158 295392 630164
rect 295352 625598 295380 630158
rect 341536 626618 341564 652734
rect 341524 626612 341576 626618
rect 341524 626554 341576 626560
rect 347044 626612 347096 626618
rect 347044 626554 347096 626560
rect 295340 625592 295392 625598
rect 295340 625534 295392 625540
rect 298100 625592 298152 625598
rect 298100 625534 298152 625540
rect 298112 620362 298140 625534
rect 298100 620356 298152 620362
rect 298100 620298 298152 620304
rect 305644 620356 305696 620362
rect 305644 620298 305696 620304
rect 294604 607912 294656 607918
rect 294604 607854 294656 607860
rect 300124 607912 300176 607918
rect 300124 607854 300176 607860
rect 249064 587240 249116 587246
rect 249064 587182 249116 587188
rect 254584 587240 254636 587246
rect 254584 587182 254636 587188
rect 218704 580984 218756 580990
rect 218704 580926 218756 580932
rect 220084 580984 220136 580990
rect 220084 580926 220136 580932
rect 204904 573300 204956 573306
rect 204904 573242 204956 573248
rect 210424 573300 210476 573306
rect 210424 573242 210476 573248
rect 204916 562358 204944 573242
rect 202144 562352 202196 562358
rect 202144 562294 202196 562300
rect 204904 562352 204956 562358
rect 204904 562294 204956 562300
rect 202156 556238 202184 562294
rect 195980 556232 196032 556238
rect 195980 556174 196032 556180
rect 202144 556232 202196 556238
rect 202144 556174 202196 556180
rect 195992 550866 196020 556174
rect 191196 550860 191248 550866
rect 191196 550802 191248 550808
rect 195980 550860 196032 550866
rect 195980 550802 196032 550808
rect 191208 547942 191236 550802
rect 188344 547936 188396 547942
rect 188344 547878 188396 547884
rect 191196 547936 191248 547942
rect 191196 547878 191248 547884
rect 188356 523530 188384 547878
rect 218716 545154 218744 580926
rect 249076 560998 249104 587182
rect 300136 572966 300164 607854
rect 305656 606490 305684 620298
rect 305644 606484 305696 606490
rect 305644 606426 305696 606432
rect 310888 606484 310940 606490
rect 310888 606426 310940 606432
rect 310900 600302 310928 606426
rect 310888 600296 310940 600302
rect 310888 600238 310940 600244
rect 315304 600296 315356 600302
rect 315304 600238 315356 600244
rect 315316 587178 315344 600238
rect 347056 592618 347084 626554
rect 347044 592612 347096 592618
rect 347044 592554 347096 592560
rect 353944 592612 353996 592618
rect 353944 592554 353996 592560
rect 315304 587172 315356 587178
rect 315304 587114 315356 587120
rect 319076 587172 319128 587178
rect 319076 587114 319128 587120
rect 319088 583030 319116 587114
rect 319076 583024 319128 583030
rect 319076 582966 319128 582972
rect 333980 583024 334032 583030
rect 333980 582966 334032 582972
rect 333992 577522 334020 582966
rect 353956 577522 353984 592554
rect 333980 577516 334032 577522
rect 333980 577458 334032 577464
rect 340144 577516 340196 577522
rect 340144 577458 340196 577464
rect 353944 577516 353996 577522
rect 353944 577458 353996 577464
rect 360844 577516 360896 577522
rect 360844 577458 360896 577464
rect 300124 572960 300176 572966
rect 300124 572902 300176 572908
rect 302884 572960 302936 572966
rect 302884 572902 302936 572908
rect 302896 563038 302924 572902
rect 340156 569226 340184 577458
rect 340144 569220 340196 569226
rect 340144 569162 340196 569168
rect 352564 569220 352616 569226
rect 352564 569162 352616 569168
rect 302884 563032 302936 563038
rect 302884 562974 302936 562980
rect 307024 563032 307076 563038
rect 307024 562974 307076 562980
rect 239404 560992 239456 560998
rect 239404 560934 239456 560940
rect 249064 560992 249116 560998
rect 249064 560934 249116 560940
rect 217416 545148 217468 545154
rect 217416 545090 217468 545096
rect 218704 545148 218756 545154
rect 218704 545090 218756 545096
rect 217428 543046 217456 545090
rect 215944 543040 215996 543046
rect 215944 542982 215996 542988
rect 217416 543040 217468 543046
rect 217416 542982 217468 542988
rect 215956 535498 215984 542982
rect 239416 542366 239444 560934
rect 233884 542360 233936 542366
rect 233884 542302 233936 542308
rect 239404 542360 239456 542366
rect 239404 542302 239456 542308
rect 214564 535492 214616 535498
rect 214564 535434 214616 535440
rect 215944 535492 215996 535498
rect 215944 535434 215996 535440
rect 185584 523524 185636 523530
rect 185584 523466 185636 523472
rect 188344 523524 188396 523530
rect 188344 523466 188396 523472
rect 185596 518226 185624 523466
rect 176660 518220 176712 518226
rect 176660 518162 176712 518168
rect 185584 518220 185636 518226
rect 185584 518162 185636 518168
rect 176672 514078 176700 518162
rect 163504 514072 163556 514078
rect 163504 514014 163556 514020
rect 176660 514072 176712 514078
rect 176660 514014 176712 514020
rect 163516 507890 163544 514014
rect 214576 513330 214604 535434
rect 233896 519586 233924 542302
rect 307036 534750 307064 562974
rect 352576 547194 352604 569162
rect 352564 547188 352616 547194
rect 352564 547130 352616 547136
rect 307024 534744 307076 534750
rect 307024 534686 307076 534692
rect 344284 534744 344336 534750
rect 344284 534686 344336 534692
rect 344296 519586 344324 534686
rect 360856 528630 360884 577458
rect 364984 547188 365036 547194
rect 364984 547130 365036 547136
rect 360844 528624 360896 528630
rect 360844 528566 360896 528572
rect 225604 519580 225656 519586
rect 225604 519522 225656 519528
rect 233884 519580 233936 519586
rect 233884 519522 233936 519528
rect 344284 519580 344336 519586
rect 344284 519522 344336 519528
rect 349712 519580 349764 519586
rect 349712 519522 349764 519528
rect 211804 513324 211856 513330
rect 211804 513266 211856 513272
rect 214564 513324 214616 513330
rect 214564 513266 214616 513272
rect 210424 508564 210476 508570
rect 210424 508506 210476 508512
rect 157984 507884 158036 507890
rect 157984 507826 158036 507832
rect 163504 507884 163556 507890
rect 163504 507826 163556 507832
rect 157996 485110 158024 507826
rect 210436 498234 210464 508506
rect 203524 498228 203576 498234
rect 203524 498170 203576 498176
rect 210424 498228 210476 498234
rect 210424 498170 210476 498176
rect 149704 485104 149756 485110
rect 149704 485046 149756 485052
rect 157984 485104 158036 485110
rect 157984 485046 158036 485052
rect 149716 461650 149744 485046
rect 141424 461644 141476 461650
rect 141424 461586 141476 461592
rect 149704 461644 149756 461650
rect 149704 461586 149756 461592
rect 141436 402286 141464 461586
rect 203536 429214 203564 498170
rect 211816 463418 211844 513266
rect 225616 508570 225644 519522
rect 349724 514758 349752 519522
rect 349712 514752 349764 514758
rect 349712 514694 349764 514700
rect 355324 514752 355376 514758
rect 355324 514694 355376 514700
rect 225604 508564 225656 508570
rect 225604 508506 225656 508512
rect 355336 485858 355364 514694
rect 355324 485852 355376 485858
rect 355324 485794 355376 485800
rect 359832 485852 359884 485858
rect 359832 485794 359884 485800
rect 359844 480758 359872 485794
rect 359832 480752 359884 480758
rect 359832 480694 359884 480700
rect 364340 480752 364392 480758
rect 364340 480694 364392 480700
rect 364352 476134 364380 480694
rect 364340 476128 364392 476134
rect 364340 476070 364392 476076
rect 364996 469878 365024 547130
rect 366364 528624 366416 528630
rect 366364 528566 366416 528572
rect 366376 494766 366404 528566
rect 366364 494760 366416 494766
rect 366364 494702 366416 494708
rect 374644 494760 374696 494766
rect 374644 494702 374696 494708
rect 374656 485110 374684 494702
rect 374644 485104 374696 485110
rect 374644 485046 374696 485052
rect 384028 485104 384080 485110
rect 384028 485046 384080 485052
rect 384040 480962 384068 485046
rect 384028 480956 384080 480962
rect 384028 480898 384080 480904
rect 393964 480956 394016 480962
rect 393964 480898 394016 480904
rect 370596 476128 370648 476134
rect 370596 476070 370648 476076
rect 364984 469872 365036 469878
rect 364984 469814 365036 469820
rect 370504 469872 370556 469878
rect 370504 469814 370556 469820
rect 210424 463412 210476 463418
rect 210424 463354 210476 463360
rect 211804 463412 211856 463418
rect 211804 463354 211856 463360
rect 210436 438938 210464 463354
rect 208400 438932 208452 438938
rect 208400 438874 208452 438880
rect 210424 438932 210476 438938
rect 210424 438874 210476 438880
rect 208412 435402 208440 438874
rect 207664 435396 207716 435402
rect 207664 435338 207716 435344
rect 208400 435396 208452 435402
rect 208400 435338 208452 435344
rect 200672 429208 200724 429214
rect 200672 429150 200724 429156
rect 203524 429208 203576 429214
rect 203524 429150 203576 429156
rect 200684 422346 200712 429150
rect 198004 422340 198056 422346
rect 198004 422282 198056 422288
rect 200672 422340 200724 422346
rect 200672 422282 200724 422288
rect 198016 415410 198044 422282
rect 193864 415404 193916 415410
rect 193864 415346 193916 415352
rect 198004 415404 198056 415410
rect 198004 415346 198056 415352
rect 141424 402280 141476 402286
rect 141424 402222 141476 402228
rect 136640 396772 136692 396778
rect 136640 396714 136692 396720
rect 191840 384668 191892 384674
rect 191840 384610 191892 384616
rect 177304 384328 177356 384334
rect 177304 384270 177356 384276
rect 123484 357060 123536 357066
rect 123484 357002 123536 357008
rect 131764 357060 131816 357066
rect 131764 357002 131816 357008
rect 111064 353320 111116 353326
rect 111064 353262 111116 353268
rect 112444 353320 112496 353326
rect 112444 353262 112496 353268
rect 111076 343670 111104 353262
rect 123496 343670 123524 357002
rect 175004 346384 175056 346390
rect 175004 346326 175056 346332
rect 109776 343664 109828 343670
rect 109776 343606 109828 343612
rect 111064 343664 111116 343670
rect 111064 343606 111116 343612
rect 117964 343664 118016 343670
rect 117964 343606 118016 343612
rect 123484 343664 123536 343670
rect 123484 343606 123536 343612
rect 109788 340066 109816 343606
rect 108304 340060 108356 340066
rect 108304 340002 108356 340008
rect 109776 340060 109828 340066
rect 109776 340002 109828 340008
rect 108316 305658 108344 340002
rect 117976 331906 118004 343606
rect 175016 339522 175044 346326
rect 171876 339516 171928 339522
rect 171876 339458 171928 339464
rect 175004 339516 175056 339522
rect 175004 339458 175056 339464
rect 171888 335510 171916 339458
rect 165436 335504 165488 335510
rect 165436 335446 165488 335452
rect 171876 335504 171928 335510
rect 171876 335446 171928 335452
rect 165448 332654 165476 335446
rect 162860 332648 162912 332654
rect 162860 332590 162912 332596
rect 165436 332648 165488 332654
rect 165436 332590 165488 332596
rect 117964 331900 118016 331906
rect 117964 331842 118016 331848
rect 162872 331294 162900 332590
rect 162860 331288 162912 331294
rect 162860 331230 162912 331236
rect 157984 331220 158036 331226
rect 157984 331162 158036 331168
rect 157996 320210 158024 331162
rect 157984 320204 158036 320210
rect 157984 320146 158036 320152
rect 154764 320136 154816 320142
rect 154764 320078 154816 320084
rect 154776 318442 154804 320078
rect 177316 319462 177344 384270
rect 191852 382294 191880 384610
rect 193876 384334 193904 415346
rect 207676 404394 207704 435338
rect 370516 424386 370544 469814
rect 370608 466002 370636 476070
rect 393976 469266 394004 480898
rect 393964 469260 394016 469266
rect 393964 469202 394016 469208
rect 396540 469260 396592 469266
rect 396540 469202 396592 469208
rect 370596 465996 370648 466002
rect 370596 465938 370648 465944
rect 373264 465996 373316 466002
rect 373264 465938 373316 465944
rect 373276 453354 373304 465938
rect 373264 453348 373316 453354
rect 373264 453290 373316 453296
rect 393964 453348 394016 453354
rect 393964 453290 394016 453296
rect 370504 424380 370556 424386
rect 370504 424322 370556 424328
rect 389824 424380 389876 424386
rect 389824 424322 389876 424328
rect 207664 404388 207716 404394
rect 207664 404330 207716 404336
rect 203892 404320 203944 404326
rect 203892 404262 203944 404268
rect 203904 397730 203932 404262
rect 389836 399158 389864 424322
rect 393976 404326 394004 453290
rect 393964 404320 394016 404326
rect 393964 404262 394016 404268
rect 389824 399152 389876 399158
rect 389824 399094 389876 399100
rect 392584 399152 392636 399158
rect 392584 399094 392636 399100
rect 201408 397724 201460 397730
rect 201408 397666 201460 397672
rect 203892 397724 203944 397730
rect 203892 397666 203944 397672
rect 201420 393378 201448 397666
rect 198740 393372 198792 393378
rect 198740 393314 198792 393320
rect 201408 393372 201460 393378
rect 201408 393314 201460 393320
rect 198752 389230 198780 393314
rect 194508 389224 194560 389230
rect 194508 389166 194560 389172
rect 198740 389224 198792 389230
rect 198740 389166 198792 389172
rect 194520 384674 194548 389166
rect 194508 384668 194560 384674
rect 194508 384610 194560 384616
rect 193864 384328 193916 384334
rect 193864 384270 193916 384276
rect 189724 382288 189776 382294
rect 189724 382230 189776 382236
rect 191840 382288 191892 382294
rect 191840 382230 191892 382236
rect 189736 362982 189764 382230
rect 392596 371210 392624 399094
rect 392584 371204 392636 371210
rect 392584 371146 392636 371152
rect 395344 371204 395396 371210
rect 395344 371146 395396 371152
rect 189724 362976 189776 362982
rect 189724 362918 189776 362924
rect 186320 362908 186372 362914
rect 186320 362850 186372 362856
rect 186332 360262 186360 362850
rect 186320 360256 186372 360262
rect 186320 360198 186372 360204
rect 182364 360188 182416 360194
rect 182364 360130 182416 360136
rect 182376 354754 182404 360130
rect 182364 354748 182416 354754
rect 182364 354690 182416 354696
rect 179420 354680 179472 354686
rect 179420 354622 179472 354628
rect 179432 346458 179460 354622
rect 179420 346452 179472 346458
rect 179420 346394 179472 346400
rect 166264 319456 166316 319462
rect 166264 319398 166316 319404
rect 177304 319456 177356 319462
rect 177304 319398 177356 319404
rect 153200 318436 153252 318442
rect 153200 318378 153252 318384
rect 154764 318436 154816 318442
rect 154764 318378 154816 318384
rect 153212 314702 153240 318378
rect 152464 314696 152516 314702
rect 152464 314638 152516 314644
rect 153200 314696 153252 314702
rect 153200 314638 153252 314644
rect 108304 305652 108356 305658
rect 108304 305594 108356 305600
rect 133144 302932 133196 302938
rect 133144 302874 133196 302880
rect 133156 293282 133184 302874
rect 124496 293276 124548 293282
rect 124496 293218 124548 293224
rect 133144 293276 133196 293282
rect 133144 293218 133196 293224
rect 104900 290488 104952 290494
rect 104900 290430 104952 290436
rect 101404 290420 101456 290426
rect 101404 290362 101456 290368
rect 102784 290420 102836 290426
rect 102784 290362 102836 290368
rect 101416 278050 101444 290362
rect 124508 288454 124536 293218
rect 122104 288448 122156 288454
rect 122104 288390 122156 288396
rect 124496 288448 124548 288454
rect 124496 288390 124548 288396
rect 101404 278044 101456 278050
rect 101404 277986 101456 277992
rect 122116 277642 122144 288390
rect 118884 277636 118936 277642
rect 118884 277578 118936 277584
rect 122104 277636 122156 277642
rect 122104 277578 122156 277584
rect 118896 273970 118924 277578
rect 112444 273964 112496 273970
rect 112444 273906 112496 273912
rect 118884 273964 118936 273970
rect 118884 273906 118936 273912
rect 112456 261526 112484 273906
rect 152476 263294 152504 314638
rect 166276 311166 166304 319398
rect 153844 311160 153896 311166
rect 153844 311102 153896 311108
rect 166264 311160 166316 311166
rect 166264 311102 166316 311108
rect 153856 302938 153884 311102
rect 153844 302932 153896 302938
rect 153844 302874 153896 302880
rect 151084 263288 151136 263294
rect 151084 263230 151136 263236
rect 152464 263288 152516 263294
rect 152464 263230 152516 263236
rect 93124 261520 93176 261526
rect 93124 261462 93176 261468
rect 112444 261520 112496 261526
rect 112444 261462 112496 261468
rect 93136 244934 93164 261462
rect 151096 255338 151124 263230
rect 143080 255332 143132 255338
rect 143080 255274 143132 255280
rect 151084 255332 151136 255338
rect 151084 255274 151136 255280
rect 143092 252346 143120 255274
rect 140044 252340 140096 252346
rect 140044 252282 140096 252288
rect 143080 252340 143132 252346
rect 143080 252282 143132 252288
rect 93124 244928 93176 244934
rect 93124 244870 93176 244876
rect 140056 244458 140084 252282
rect 138020 244452 138072 244458
rect 138020 244394 138072 244400
rect 140044 244452 140096 244458
rect 140044 244394 140096 244400
rect 88340 240848 88392 240854
rect 88340 240790 88392 240796
rect 138032 240786 138060 244394
rect 138020 240780 138072 240786
rect 138020 240722 138072 240728
rect 395356 240106 395384 371146
rect 395344 240100 395396 240106
rect 395344 240042 395396 240048
rect 396448 240100 396500 240106
rect 396448 240042 396500 240048
rect 80060 239828 80112 239834
rect 80060 239770 80112 239776
rect 45836 238808 45888 238814
rect 45836 238750 45888 238756
rect 45836 233232 45888 233238
rect 45836 233174 45888 233180
rect 45848 231130 45876 233174
rect 86224 232416 86276 232422
rect 86224 232358 86276 232364
rect 394148 232416 394200 232422
rect 394148 232358 394200 232364
rect 45836 231124 45888 231130
rect 45836 231066 45888 231072
rect 49700 231124 49752 231130
rect 49700 231066 49752 231072
rect 49712 229158 49740 231066
rect 86236 230858 86264 232358
rect 393964 231872 394016 231878
rect 393964 231814 394016 231820
rect 180800 231192 180852 231198
rect 180800 231134 180852 231140
rect 384396 231192 384448 231198
rect 384396 231134 384448 231140
rect 118608 231124 118660 231130
rect 118608 231066 118660 231072
rect 86224 230852 86276 230858
rect 86224 230794 86276 230800
rect 88892 230852 88944 230858
rect 88892 230794 88944 230800
rect 54484 230444 54536 230450
rect 54484 230386 54536 230392
rect 53104 229764 53156 229770
rect 53104 229706 53156 229712
rect 49700 229152 49752 229158
rect 49700 229094 49752 229100
rect 52460 229084 52512 229090
rect 52460 229026 52512 229032
rect 47400 227248 47452 227254
rect 47400 227190 47452 227196
rect 47412 220794 47440 227190
rect 52472 226370 52500 229026
rect 53116 228410 53144 229706
rect 53104 228404 53156 228410
rect 53104 228346 53156 228352
rect 52460 226364 52512 226370
rect 52460 226306 52512 226312
rect 47584 224936 47636 224942
rect 47584 224878 47636 224884
rect 47400 220788 47452 220794
rect 47400 220730 47452 220736
rect 45652 205216 45704 205222
rect 45652 205158 45704 205164
rect 47596 201482 47624 224878
rect 49608 220788 49660 220794
rect 49608 220730 49660 220736
rect 49620 219434 49648 220730
rect 49620 219406 49740 219434
rect 49712 214810 49740 219406
rect 54496 218278 54524 230386
rect 54484 218272 54536 218278
rect 54484 218214 54536 218220
rect 49700 214804 49752 214810
rect 49700 214746 49752 214752
rect 53104 214804 53156 214810
rect 53104 214746 53156 214752
rect 53116 207058 53144 214746
rect 53104 207052 53156 207058
rect 53104 206994 53156 207000
rect 55864 206984 55916 206990
rect 55864 206926 55916 206932
rect 49608 205216 49660 205222
rect 49608 205158 49660 205164
rect 49620 202842 49648 205158
rect 49608 202836 49660 202842
rect 49608 202778 49660 202784
rect 53840 202836 53892 202842
rect 53840 202778 53892 202784
rect 47584 201476 47636 201482
rect 47584 201418 47636 201424
rect 50344 201476 50396 201482
rect 50344 201418 50396 201424
rect 50356 190942 50384 201418
rect 53852 197334 53880 202778
rect 53840 197328 53892 197334
rect 53840 197270 53892 197276
rect 50344 190936 50396 190942
rect 50344 190878 50396 190884
rect 55876 182170 55904 206926
rect 56612 195974 56640 230588
rect 58900 228404 58952 228410
rect 58900 228346 58952 228352
rect 56692 226296 56744 226302
rect 56692 226238 56744 226244
rect 56704 222222 56732 226238
rect 58912 224262 58940 228346
rect 58900 224256 58952 224262
rect 58900 224198 58952 224204
rect 63500 224256 63552 224262
rect 63500 224198 63552 224204
rect 56692 222216 56744 222222
rect 56692 222158 56744 222164
rect 60648 222148 60700 222154
rect 60648 222090 60700 222096
rect 56692 218272 56744 218278
rect 56692 218214 56744 218220
rect 56704 212498 56732 218214
rect 60660 217802 60688 222090
rect 63512 220182 63540 224198
rect 63500 220176 63552 220182
rect 63500 220118 63552 220124
rect 68284 220176 68336 220182
rect 68284 220118 68336 220124
rect 60648 217796 60700 217802
rect 60648 217738 60700 217744
rect 64144 217796 64196 217802
rect 64144 217738 64196 217744
rect 56692 212492 56744 212498
rect 56692 212434 56744 212440
rect 58716 212492 58768 212498
rect 58716 212434 58768 212440
rect 58728 208418 58756 212434
rect 58716 208412 58768 208418
rect 58716 208354 58768 208360
rect 61384 208412 61436 208418
rect 61384 208354 61436 208360
rect 57704 197328 57756 197334
rect 57704 197270 57756 197276
rect 56600 195968 56652 195974
rect 56600 195910 56652 195916
rect 57716 193186 57744 197270
rect 57704 193180 57756 193186
rect 57704 193122 57756 193128
rect 57244 190936 57296 190942
rect 57244 190878 57296 190884
rect 55864 182164 55916 182170
rect 55864 182106 55916 182112
rect 57256 170134 57284 190878
rect 58624 182164 58676 182170
rect 58624 182106 58676 182112
rect 57244 170128 57296 170134
rect 57244 170070 57296 170076
rect 58636 159458 58664 182106
rect 61396 178022 61424 208354
rect 64156 204270 64184 217738
rect 64144 204264 64196 204270
rect 64144 204206 64196 204212
rect 65524 204264 65576 204270
rect 65524 204206 65576 204212
rect 65536 196722 65564 204206
rect 65524 196716 65576 196722
rect 65524 196658 65576 196664
rect 66904 196716 66956 196722
rect 66904 196658 66956 196664
rect 61752 193180 61804 193186
rect 61752 193122 61804 193128
rect 61764 184890 61792 193122
rect 61752 184884 61804 184890
rect 61752 184826 61804 184832
rect 64972 184884 65024 184890
rect 64972 184826 65024 184832
rect 64984 181490 65012 184826
rect 66916 183530 66944 196658
rect 68296 184890 68324 220118
rect 86972 195906 87000 230588
rect 88904 225010 88932 230794
rect 117240 228410 117268 230588
rect 117228 228404 117280 228410
rect 117228 228346 117280 228352
rect 88892 225004 88944 225010
rect 88892 224946 88944 224952
rect 91100 224936 91152 224942
rect 91100 224878 91152 224884
rect 91112 219502 91140 224878
rect 91100 219496 91152 219502
rect 91100 219438 91152 219444
rect 95148 219428 95200 219434
rect 95148 219370 95200 219376
rect 95160 216646 95188 219370
rect 95148 216640 95200 216646
rect 95148 216582 95200 216588
rect 98092 216640 98144 216646
rect 98092 216582 98144 216588
rect 98104 213926 98132 216582
rect 98092 213920 98144 213926
rect 98092 213862 98144 213868
rect 104164 213920 104216 213926
rect 104164 213862 104216 213868
rect 104176 211818 104204 213862
rect 104164 211812 104216 211818
rect 104164 211754 104216 211760
rect 108304 211812 108356 211818
rect 108304 211754 108356 211760
rect 86960 195900 87012 195906
rect 86960 195842 87012 195848
rect 68284 184884 68336 184890
rect 68284 184826 68336 184832
rect 72424 184884 72476 184890
rect 72424 184826 72476 184832
rect 66904 183524 66956 183530
rect 66904 183466 66956 183472
rect 68284 183524 68336 183530
rect 68284 183466 68336 183472
rect 64972 181484 65024 181490
rect 64972 181426 65024 181432
rect 61384 178016 61436 178022
rect 61384 177958 61436 177964
rect 65892 178016 65944 178022
rect 65892 177958 65944 177964
rect 65904 173874 65932 177958
rect 65892 173868 65944 173874
rect 65892 173810 65944 173816
rect 66904 173868 66956 173874
rect 66904 173810 66956 173816
rect 60648 170128 60700 170134
rect 60648 170070 60700 170076
rect 60660 166666 60688 170070
rect 60648 166660 60700 166666
rect 60648 166602 60700 166608
rect 62120 166660 62172 166666
rect 62120 166602 62172 166608
rect 62132 162246 62160 166602
rect 66916 162858 66944 173810
rect 68296 168638 68324 183466
rect 72436 179382 72464 184826
rect 75184 181484 75236 181490
rect 75184 181426 75236 181432
rect 72424 179376 72476 179382
rect 72424 179318 72476 179324
rect 68284 168632 68336 168638
rect 68284 168574 68336 168580
rect 69756 168632 69808 168638
rect 69756 168574 69808 168580
rect 69768 165578 69796 168574
rect 69756 165572 69808 165578
rect 69756 165514 69808 165520
rect 71044 165572 71096 165578
rect 71044 165514 71096 165520
rect 66904 162852 66956 162858
rect 66904 162794 66956 162800
rect 68284 162852 68336 162858
rect 68284 162794 68336 162800
rect 62120 162240 62172 162246
rect 62120 162182 62172 162188
rect 58624 159452 58676 159458
rect 58624 159394 58676 159400
rect 45284 141568 45336 141574
rect 45284 141510 45336 141516
rect 68296 127634 68324 162794
rect 71056 153202 71084 165514
rect 75196 163538 75224 181426
rect 75736 179376 75788 179382
rect 75736 179318 75788 179324
rect 75748 177002 75776 179318
rect 75736 176996 75788 177002
rect 75736 176938 75788 176944
rect 77300 176996 77352 177002
rect 77300 176938 77352 176944
rect 77312 173942 77340 176938
rect 77300 173936 77352 173942
rect 77300 173878 77352 173884
rect 81348 173868 81400 173874
rect 81348 173810 81400 173816
rect 81360 168450 81388 173810
rect 81360 168422 81480 168450
rect 81452 165578 81480 168422
rect 81440 165572 81492 165578
rect 81440 165514 81492 165520
rect 83464 165572 83516 165578
rect 83464 165514 83516 165520
rect 75184 163532 75236 163538
rect 75184 163474 75236 163480
rect 81440 159452 81492 159458
rect 81440 159394 81492 159400
rect 81452 158030 81480 159394
rect 81440 158024 81492 158030
rect 81440 157966 81492 157972
rect 83476 157350 83504 165514
rect 86224 163532 86276 163538
rect 86224 163474 86276 163480
rect 84752 158024 84804 158030
rect 84752 157966 84804 157972
rect 83464 157344 83516 157350
rect 83464 157286 83516 157292
rect 84764 156670 84792 157966
rect 84844 157344 84896 157350
rect 84844 157286 84896 157292
rect 84752 156664 84804 156670
rect 84752 156606 84804 156612
rect 71044 153196 71096 153202
rect 71044 153138 71096 153144
rect 73804 153196 73856 153202
rect 73804 153138 73856 153144
rect 68284 127628 68336 127634
rect 68284 127570 68336 127576
rect 71044 127628 71096 127634
rect 71044 127570 71096 127576
rect 71056 117978 71084 127570
rect 73816 124846 73844 153138
rect 84856 131782 84884 157286
rect 86236 149258 86264 163474
rect 87604 162240 87656 162246
rect 87604 162182 87656 162188
rect 87616 154562 87644 162182
rect 89076 156664 89128 156670
rect 89076 156606 89128 156612
rect 87604 154556 87656 154562
rect 87604 154498 87656 154504
rect 89088 149870 89116 156606
rect 90364 154556 90416 154562
rect 90364 154498 90416 154504
rect 89076 149864 89128 149870
rect 89076 149806 89128 149812
rect 86224 149252 86276 149258
rect 86224 149194 86276 149200
rect 88984 149252 89036 149258
rect 88984 149194 89036 149200
rect 88996 139534 89024 149194
rect 88984 139528 89036 139534
rect 88984 139470 89036 139476
rect 90376 135930 90404 154498
rect 91008 149864 91060 149870
rect 91008 149806 91060 149812
rect 91020 149054 91048 149806
rect 91008 149048 91060 149054
rect 91008 148990 91060 148996
rect 92480 149048 92532 149054
rect 92480 148990 92532 148996
rect 92492 142866 92520 148990
rect 108316 146266 108344 211754
rect 108396 162920 108448 162926
rect 108396 162862 108448 162868
rect 108304 146260 108356 146266
rect 108304 146202 108356 146208
rect 92480 142860 92532 142866
rect 92480 142802 92532 142808
rect 104900 142860 104952 142866
rect 104900 142802 104952 142808
rect 104912 141438 104940 142802
rect 104900 141432 104952 141438
rect 104900 141374 104952 141380
rect 107660 141432 107712 141438
rect 107660 141374 107712 141380
rect 107672 140146 107700 141374
rect 107660 140140 107712 140146
rect 107660 140082 107712 140088
rect 91376 139528 91428 139534
rect 91376 139470 91428 139476
rect 90364 135924 90416 135930
rect 90364 135866 90416 135872
rect 91388 132870 91416 139470
rect 105544 135924 105596 135930
rect 105544 135866 105596 135872
rect 97264 135312 97316 135318
rect 97264 135254 97316 135260
rect 91376 132864 91428 132870
rect 91376 132806 91428 132812
rect 94228 132864 94280 132870
rect 94228 132806 94280 132812
rect 84844 131776 84896 131782
rect 84844 131718 84896 131724
rect 86316 131776 86368 131782
rect 86316 131718 86368 131724
rect 86328 130898 86356 131718
rect 86316 130892 86368 130898
rect 86316 130834 86368 130840
rect 87604 130892 87656 130898
rect 87604 130834 87656 130840
rect 73804 124840 73856 124846
rect 73804 124782 73856 124788
rect 75828 124840 75880 124846
rect 75828 124782 75880 124788
rect 75840 122834 75868 124782
rect 75840 122806 75960 122834
rect 75932 119134 75960 122806
rect 87616 121854 87644 130834
rect 94240 126886 94268 132806
rect 94228 126880 94280 126886
rect 94228 126822 94280 126828
rect 87604 121848 87656 121854
rect 87604 121790 87656 121796
rect 91008 121848 91060 121854
rect 91008 121790 91060 121796
rect 91020 121394 91048 121790
rect 91020 121366 91140 121394
rect 91112 119950 91140 121366
rect 91100 119944 91152 119950
rect 91100 119886 91152 119892
rect 93124 119944 93176 119950
rect 93124 119886 93176 119892
rect 75920 119128 75972 119134
rect 75920 119070 75972 119076
rect 78588 119128 78640 119134
rect 78588 119070 78640 119076
rect 71044 117972 71096 117978
rect 71044 117914 71096 117920
rect 77300 117972 77352 117978
rect 77300 117914 77352 117920
rect 77312 116074 77340 117914
rect 77300 116068 77352 116074
rect 77300 116010 77352 116016
rect 78600 114510 78628 119070
rect 79324 116068 79376 116074
rect 79324 116010 79376 116016
rect 78588 114504 78640 114510
rect 78588 114446 78640 114452
rect 79336 112470 79364 116010
rect 93136 113150 93164 119886
rect 93124 113144 93176 113150
rect 93124 113086 93176 113092
rect 79324 112464 79376 112470
rect 79324 112406 79376 112412
rect 88248 112464 88300 112470
rect 88248 112406 88300 112412
rect 88260 111790 88288 112406
rect 88248 111784 88300 111790
rect 88248 111726 88300 111732
rect 89720 78124 89772 78130
rect 89720 78066 89772 78072
rect 71780 78056 71832 78062
rect 71780 77998 71832 78004
rect 53840 77988 53892 77994
rect 53840 77930 53892 77936
rect 44916 75880 44968 75886
rect 44916 75822 44968 75828
rect 51080 73908 51132 73914
rect 51080 73850 51132 73856
rect 49700 71120 49752 71126
rect 49700 71062 49752 71068
rect 45560 47592 45612 47598
rect 45560 47534 45612 47540
rect 45572 16574 45600 47534
rect 49712 16574 49740 71062
rect 45572 16546 46704 16574
rect 49712 16546 50200 16574
rect 44272 10328 44324 10334
rect 44272 10270 44324 10276
rect 44180 3392 44232 3398
rect 44180 3334 44232 3340
rect 44284 480 44312 10270
rect 45100 3392 45152 3398
rect 45100 3334 45152 3340
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45112 354 45140 3334
rect 46676 480 46704 16546
rect 48964 4956 49016 4962
rect 48964 4898 49016 4904
rect 47860 3732 47912 3738
rect 47860 3674 47912 3680
rect 47872 480 47900 3674
rect 48976 480 49004 4898
rect 50172 480 50200 16546
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 73850
rect 52460 69760 52512 69766
rect 52460 69702 52512 69708
rect 52472 16574 52500 69702
rect 53852 16574 53880 77930
rect 70400 75404 70452 75410
rect 70400 75346 70452 75352
rect 60740 75336 60792 75342
rect 60740 75278 60792 75284
rect 57978 73944 58034 73953
rect 57978 73879 58034 73888
rect 55218 68232 55274 68241
rect 55218 68167 55274 68176
rect 55232 16574 55260 68167
rect 57992 16574 58020 73879
rect 59360 68332 59412 68338
rect 59360 68274 59412 68280
rect 52472 16546 53328 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 57992 16546 58480 16574
rect 52552 5024 52604 5030
rect 52552 4966 52604 4972
rect 52564 480 52592 4966
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 57242 9072 57298 9081
rect 57242 9007 57298 9016
rect 57256 480 57284 9007
rect 58452 480 58480 16546
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59372 354 59400 68274
rect 60752 3398 60780 75278
rect 69020 72684 69072 72690
rect 69020 72626 69072 72632
rect 64880 66972 64932 66978
rect 64880 66914 64932 66920
rect 60832 22840 60884 22846
rect 60832 22782 60884 22788
rect 60740 3392 60792 3398
rect 60740 3334 60792 3340
rect 60844 480 60872 22782
rect 64892 16574 64920 66914
rect 67640 22908 67692 22914
rect 67640 22850 67692 22856
rect 64892 16546 65104 16574
rect 63224 6248 63276 6254
rect 63224 6190 63276 6196
rect 61660 3392 61712 3398
rect 61660 3334 61712 3340
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3334
rect 63236 480 63264 6190
rect 64328 3800 64380 3806
rect 64328 3742 64380 3748
rect 64340 480 64368 3742
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66720 5092 66772 5098
rect 66720 5034 66772 5040
rect 66732 480 66760 5034
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 22850
rect 69032 16574 69060 72626
rect 70412 16574 70440 75346
rect 71792 16574 71820 77998
rect 86960 76696 87012 76702
rect 86960 76638 87012 76644
rect 75918 72448 75974 72457
rect 75918 72383 75974 72392
rect 73158 69592 73214 69601
rect 73158 69527 73214 69536
rect 73172 16574 73200 69527
rect 69032 16546 69152 16574
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 69124 480 69152 16546
rect 70308 6316 70360 6322
rect 70308 6258 70360 6264
rect 70320 480 70348 6258
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 74998 9208 75054 9217
rect 74998 9143 75054 9152
rect 75012 480 75040 9143
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 72383
rect 82820 69896 82872 69902
rect 82820 69838 82872 69844
rect 78680 69828 78732 69834
rect 78680 69770 78732 69776
rect 78692 16574 78720 69770
rect 81440 44872 81492 44878
rect 81440 44814 81492 44820
rect 81452 16574 81480 44814
rect 82832 16574 82860 69838
rect 85580 68400 85632 68406
rect 85580 68342 85632 68348
rect 85592 16574 85620 68342
rect 86972 16574 87000 76638
rect 88340 43444 88392 43450
rect 88340 43386 88392 43392
rect 88352 16574 88380 43386
rect 89732 16574 89760 78066
rect 93858 76664 93914 76673
rect 93858 76599 93914 76608
rect 91098 68368 91154 68377
rect 91098 68303 91154 68312
rect 91112 16574 91140 68303
rect 78692 16546 79272 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 85592 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 78588 6384 78640 6390
rect 78588 6326 78640 6332
rect 77392 3868 77444 3874
rect 77392 3810 77444 3816
rect 77404 480 77432 3810
rect 78600 480 78628 6326
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79244 354 79272 16546
rect 80888 6452 80940 6458
rect 80888 6394 80940 6400
rect 80900 480 80928 6394
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 84476 6520 84528 6526
rect 84476 6462 84528 6468
rect 84488 480 84516 6462
rect 85672 5160 85724 5166
rect 85672 5102 85724 5108
rect 85684 480 85712 5102
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 92478 10296 92534 10305
rect 92478 10231 92534 10240
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 10231
rect 93872 3398 93900 76599
rect 93952 73976 94004 73982
rect 93952 73918 94004 73924
rect 93860 3392 93912 3398
rect 93860 3334 93912 3340
rect 93964 480 93992 73918
rect 97276 71738 97304 135254
rect 105556 126886 105584 135866
rect 108408 133890 108436 162862
rect 118240 156664 118292 156670
rect 118240 156606 118292 156612
rect 109684 146260 109736 146266
rect 109684 146202 109736 146208
rect 108396 133884 108448 133890
rect 108396 133826 108448 133832
rect 109696 129810 109724 146202
rect 118148 142860 118200 142866
rect 118148 142802 118200 142808
rect 117964 141432 118016 141438
rect 117964 141374 118016 141380
rect 117318 137592 117374 137601
rect 117318 137527 117374 137536
rect 117332 136746 117360 137527
rect 117320 136740 117372 136746
rect 117320 136682 117372 136688
rect 117318 136096 117374 136105
rect 117318 136031 117374 136040
rect 117332 135318 117360 136031
rect 117320 135312 117372 135318
rect 117320 135254 117372 135260
rect 117318 134600 117374 134609
rect 117318 134535 117374 134544
rect 117332 133958 117360 134535
rect 117320 133952 117372 133958
rect 117320 133894 117372 133900
rect 117412 133884 117464 133890
rect 117412 133826 117464 133832
rect 117424 133113 117452 133826
rect 117410 133104 117466 133113
rect 117410 133039 117466 133048
rect 117320 132456 117372 132462
rect 117320 132398 117372 132404
rect 117332 131617 117360 132398
rect 117318 131608 117374 131617
rect 117318 131543 117374 131552
rect 117320 131096 117372 131102
rect 117320 131038 117372 131044
rect 117332 130121 117360 131038
rect 117318 130112 117374 130121
rect 117318 130047 117374 130056
rect 109684 129804 109736 129810
rect 109684 129746 109736 129752
rect 111064 129804 111116 129810
rect 111064 129746 111116 129752
rect 100024 126880 100076 126886
rect 100024 126822 100076 126828
rect 105544 126880 105596 126886
rect 105544 126822 105596 126828
rect 109684 126880 109736 126886
rect 109684 126822 109736 126828
rect 100036 115938 100064 126822
rect 109696 122534 109724 126822
rect 109684 122528 109736 122534
rect 109684 122470 109736 122476
rect 100024 115932 100076 115938
rect 100024 115874 100076 115880
rect 111076 109070 111104 129746
rect 117320 129736 117372 129742
rect 117320 129678 117372 129684
rect 117332 128625 117360 129678
rect 117318 128616 117374 128625
rect 117318 128551 117374 128560
rect 117320 128308 117372 128314
rect 117320 128250 117372 128256
rect 117332 127129 117360 128250
rect 117318 127120 117374 127129
rect 117318 127055 117374 127064
rect 117320 126948 117372 126954
rect 117320 126890 117372 126896
rect 117332 125633 117360 126890
rect 117318 125624 117374 125633
rect 117318 125559 117374 125568
rect 117320 124160 117372 124166
rect 117318 124128 117320 124137
rect 117372 124128 117374 124137
rect 117318 124063 117374 124072
rect 117320 122800 117372 122806
rect 117320 122742 117372 122748
rect 117332 122641 117360 122742
rect 117318 122632 117374 122641
rect 117318 122567 117374 122576
rect 113824 122528 113876 122534
rect 113824 122470 113876 122476
rect 113836 109070 113864 122470
rect 117320 121440 117372 121446
rect 117320 121382 117372 121388
rect 117332 121145 117360 121382
rect 117318 121136 117374 121145
rect 117318 121071 117374 121080
rect 117320 120080 117372 120086
rect 117320 120022 117372 120028
rect 117332 119649 117360 120022
rect 117318 119640 117374 119649
rect 117318 119575 117374 119584
rect 117320 118652 117372 118658
rect 117320 118594 117372 118600
rect 117332 118153 117360 118594
rect 117318 118144 117374 118153
rect 117318 118079 117374 118088
rect 117320 117292 117372 117298
rect 117320 117234 117372 117240
rect 117332 116657 117360 117234
rect 117318 116648 117374 116657
rect 117318 116583 117374 116592
rect 117320 115932 117372 115938
rect 117320 115874 117372 115880
rect 117332 115161 117360 115874
rect 117318 115152 117374 115161
rect 117318 115087 117374 115096
rect 117320 114504 117372 114510
rect 117320 114446 117372 114452
rect 117332 113665 117360 114446
rect 117318 113656 117374 113665
rect 117318 113591 117374 113600
rect 117320 113144 117372 113150
rect 117320 113086 117372 113092
rect 117332 112169 117360 113086
rect 117318 112160 117374 112169
rect 117318 112095 117374 112104
rect 117320 111784 117372 111790
rect 117320 111726 117372 111732
rect 117332 110673 117360 111726
rect 117318 110664 117374 110673
rect 117318 110599 117374 110608
rect 111064 109064 111116 109070
rect 111064 109006 111116 109012
rect 112444 109064 112496 109070
rect 112444 109006 112496 109012
rect 113824 109064 113876 109070
rect 113824 109006 113876 109012
rect 112456 103154 112484 109006
rect 117976 103193 118004 141374
rect 118056 139528 118108 139534
rect 118056 139470 118108 139476
rect 117962 103184 118018 103193
rect 112444 103148 112496 103154
rect 112444 103090 112496 103096
rect 115388 103148 115440 103154
rect 117962 103119 118018 103128
rect 115388 103090 115440 103096
rect 115400 100366 115428 103090
rect 115388 100360 115440 100366
rect 115388 100302 115440 100308
rect 117320 100360 117372 100366
rect 117320 100302 117372 100308
rect 117332 97986 117360 100302
rect 117320 97980 117372 97986
rect 117320 97922 117372 97928
rect 118068 89729 118096 139470
rect 118054 89720 118110 89729
rect 118054 89655 118110 89664
rect 118160 88233 118188 142802
rect 118252 95713 118280 156606
rect 118332 155236 118384 155242
rect 118332 155178 118384 155184
rect 118238 95704 118294 95713
rect 118238 95639 118294 95648
rect 118344 94217 118372 155178
rect 118516 153876 118568 153882
rect 118516 153818 118568 153824
rect 118424 152516 118476 152522
rect 118424 152458 118476 152464
rect 118330 94208 118386 94217
rect 118330 94143 118386 94152
rect 118436 91225 118464 152458
rect 118528 92721 118556 153818
rect 118620 109177 118648 231066
rect 150440 231056 150492 231062
rect 150440 230998 150492 231004
rect 120816 229764 120868 229770
rect 120816 229706 120868 229712
rect 120724 227044 120776 227050
rect 120724 226986 120776 226992
rect 118700 224256 118752 224262
rect 118700 224198 118752 224204
rect 118606 109168 118662 109177
rect 118606 109103 118662 109112
rect 118712 98705 118740 224198
rect 119344 187740 119396 187746
rect 119344 187682 119396 187688
rect 118792 151088 118844 151094
rect 118792 151030 118844 151036
rect 118804 100201 118832 151030
rect 118976 145580 119028 145586
rect 118976 145522 119028 145528
rect 118884 144220 118936 144226
rect 118884 144162 118936 144168
rect 118896 104689 118924 144162
rect 118988 106185 119016 145522
rect 118974 106176 119030 106185
rect 118974 106111 119030 106120
rect 118882 104680 118938 104689
rect 118882 104615 118938 104624
rect 118790 100192 118846 100201
rect 118790 100127 118846 100136
rect 118698 98696 118754 98705
rect 118698 98631 118754 98640
rect 118514 92712 118570 92721
rect 118514 92647 118570 92656
rect 118422 91216 118478 91225
rect 118422 91151 118478 91160
rect 118146 88224 118202 88233
rect 118146 88159 118202 88168
rect 118514 86728 118570 86737
rect 118514 86663 118570 86672
rect 118422 83736 118478 83745
rect 118422 83671 118478 83680
rect 118330 82240 118386 82249
rect 118330 82175 118386 82184
rect 116860 79756 116912 79762
rect 116860 79698 116912 79704
rect 116872 79490 116900 79698
rect 116860 79484 116912 79490
rect 116860 79426 116912 79432
rect 106924 78260 106976 78266
rect 106924 78202 106976 78208
rect 102140 76764 102192 76770
rect 102140 76706 102192 76712
rect 97264 71732 97316 71738
rect 97264 71674 97316 71680
rect 100760 71256 100812 71262
rect 100760 71198 100812 71204
rect 96620 71188 96672 71194
rect 96620 71130 96672 71136
rect 95240 55888 95292 55894
rect 95240 55830 95292 55836
rect 95252 16574 95280 55830
rect 96632 16574 96660 71130
rect 99380 19984 99432 19990
rect 99380 19926 99432 19932
rect 99392 16574 99420 19926
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 99392 16546 99880 16574
rect 94780 3392 94832 3398
rect 94780 3334 94832 3340
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 3334
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 98644 7812 98696 7818
rect 98644 7754 98696 7760
rect 98656 480 98684 7754
rect 99852 480 99880 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 100772 354 100800 71198
rect 102152 6914 102180 76706
rect 103520 72752 103572 72758
rect 103520 72694 103572 72700
rect 102232 60036 102284 60042
rect 102232 59978 102284 59984
rect 102244 16574 102272 59978
rect 103532 16574 103560 72694
rect 106280 24132 106332 24138
rect 106280 24074 106332 24080
rect 106292 16574 106320 24074
rect 102244 16546 103376 16574
rect 103532 16546 104112 16574
rect 106292 16546 106504 16574
rect 102152 6886 102272 6914
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105728 7880 105780 7886
rect 105728 7822 105780 7828
rect 105740 480 105768 7822
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 106936 10402 106964 78202
rect 110420 78192 110472 78198
rect 110420 78134 110472 78140
rect 113822 78160 113878 78169
rect 107660 75472 107712 75478
rect 107660 75414 107712 75420
rect 107672 16574 107700 75414
rect 107672 16546 108160 16574
rect 106924 10396 106976 10402
rect 106924 10338 106976 10344
rect 108132 480 108160 16546
rect 109314 7712 109370 7721
rect 109314 7647 109370 7656
rect 109328 480 109356 7647
rect 110432 3398 110460 78134
rect 113822 78095 113878 78104
rect 111798 76800 111854 76809
rect 111798 76735 111854 76744
rect 111812 16574 111840 76735
rect 111812 16546 112392 16574
rect 110512 10464 110564 10470
rect 110512 10406 110564 10412
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 110524 480 110552 10406
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 111628 480 111656 3334
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 113836 13122 113864 78095
rect 114560 72820 114612 72826
rect 114560 72762 114612 72768
rect 114572 16574 114600 72762
rect 115940 68468 115992 68474
rect 115940 68410 115992 68416
rect 115952 16574 115980 68410
rect 118344 61402 118372 82175
rect 118332 61396 118384 61402
rect 118332 61338 118384 61344
rect 118436 46918 118464 83671
rect 118528 80481 118556 86663
rect 118606 85232 118662 85241
rect 118606 85167 118662 85176
rect 118620 80782 118648 85167
rect 118608 80776 118660 80782
rect 118608 80718 118660 80724
rect 118514 80472 118570 80481
rect 118514 80407 118570 80416
rect 119356 79218 119384 187682
rect 120632 109064 120684 109070
rect 120632 109006 120684 109012
rect 120644 108361 120672 109006
rect 120630 108352 120686 108361
rect 120630 108287 120686 108296
rect 120736 97753 120764 226986
rect 120828 102105 120856 229706
rect 143540 228404 143592 228410
rect 143540 228346 143592 228352
rect 140044 227792 140096 227798
rect 140044 227734 140096 227740
rect 122104 205692 122156 205698
rect 122104 205634 122156 205640
rect 121460 178696 121512 178702
rect 121460 178638 121512 178644
rect 121000 149728 121052 149734
rect 121000 149670 121052 149676
rect 120908 136672 120960 136678
rect 120908 136614 120960 136620
rect 120814 102096 120870 102105
rect 120814 102031 120870 102040
rect 120816 97980 120868 97986
rect 120816 97922 120868 97928
rect 120722 97744 120778 97753
rect 120722 97679 120778 97688
rect 120264 84244 120316 84250
rect 120264 84186 120316 84192
rect 120276 79422 120304 84186
rect 120828 80646 120856 97922
rect 120816 80640 120868 80646
rect 120816 80582 120868 80588
rect 120920 79558 120948 136614
rect 121012 107681 121040 149670
rect 121472 139890 121500 178638
rect 121472 139862 121808 139890
rect 122116 139534 122144 205634
rect 140056 199442 140084 227734
rect 143552 200705 143580 228346
rect 146496 227798 146524 230588
rect 150452 229498 150480 230998
rect 176672 229838 176700 230588
rect 163504 229832 163556 229838
rect 163504 229774 163556 229780
rect 176660 229832 176712 229838
rect 176660 229774 176712 229780
rect 150440 229492 150492 229498
rect 150440 229434 150492 229440
rect 153200 229492 153252 229498
rect 153200 229434 153252 229440
rect 144920 227792 144972 227798
rect 144920 227734 144972 227740
rect 146484 227792 146536 227798
rect 146484 227734 146536 227740
rect 143538 200696 143594 200705
rect 143538 200631 143594 200640
rect 140044 199436 140096 199442
rect 140044 199378 140096 199384
rect 144932 196466 144960 227734
rect 153212 226574 153240 229434
rect 161388 228404 161440 228410
rect 161388 228346 161440 228352
rect 153200 226568 153252 226574
rect 153200 226510 153252 226516
rect 155960 226568 156012 226574
rect 155960 226510 156012 226516
rect 155972 223582 156000 226510
rect 155960 223576 156012 223582
rect 155960 223518 156012 223524
rect 157984 223576 158036 223582
rect 157984 223518 158036 223524
rect 157996 208418 158024 223518
rect 157984 208412 158036 208418
rect 157984 208354 158036 208360
rect 155224 203584 155276 203590
rect 155224 203526 155276 203532
rect 153200 202156 153252 202162
rect 153200 202098 153252 202104
rect 148968 198076 149020 198082
rect 148968 198018 149020 198024
rect 147494 196480 147550 196489
rect 144932 196438 145774 196466
rect 147430 196438 147494 196466
rect 148980 196452 149008 198018
rect 147494 196415 147550 196424
rect 138112 195968 138164 195974
rect 153212 195945 153240 202098
rect 153290 196208 153346 196217
rect 153290 196143 153346 196152
rect 138112 195910 138164 195916
rect 139398 195936 139454 195945
rect 138124 195809 138152 195910
rect 139398 195871 139400 195880
rect 139452 195871 139454 195880
rect 142342 195936 142398 195945
rect 153198 195936 153254 195945
rect 142398 195894 142554 195922
rect 142342 195871 142398 195880
rect 153198 195871 153254 195880
rect 139400 195842 139452 195848
rect 138110 195800 138166 195809
rect 138110 195735 138166 195744
rect 140778 195800 140834 195809
rect 140834 195758 140990 195786
rect 140778 195735 140834 195744
rect 150348 195696 150400 195702
rect 150346 195664 150348 195673
rect 150400 195664 150402 195673
rect 150346 195599 150402 195608
rect 153304 193633 153332 196143
rect 153934 195936 153990 195945
rect 153778 195894 153934 195922
rect 153934 195871 153990 195880
rect 155236 194721 155264 203526
rect 155960 200796 156012 200802
rect 155960 200738 156012 200744
rect 155972 195945 156000 200738
rect 159824 198008 159876 198014
rect 159824 197950 159876 197956
rect 158260 196648 158312 196654
rect 158260 196590 158312 196596
rect 158272 195945 158300 196590
rect 155958 195936 156014 195945
rect 155958 195871 156014 195880
rect 158258 195936 158314 195945
rect 158902 195936 158958 195945
rect 158562 195894 158902 195922
rect 158258 195871 158314 195880
rect 158902 195871 158958 195880
rect 159836 195809 159864 197950
rect 161400 195945 161428 228346
rect 162124 208344 162176 208350
rect 162124 208286 162176 208292
rect 162136 196042 162164 208286
rect 163516 199345 163544 229774
rect 166264 228472 166316 228478
rect 166264 228414 166316 228420
rect 166276 200802 166304 228414
rect 179512 220108 179564 220114
rect 179512 220050 179564 220056
rect 166264 200796 166316 200802
rect 166264 200738 166316 200744
rect 164240 199436 164292 199442
rect 164240 199378 164292 199384
rect 163502 199336 163558 199345
rect 163502 199271 163558 199280
rect 162124 196036 162176 196042
rect 162124 195978 162176 195984
rect 161386 195936 161442 195945
rect 161386 195871 161442 195880
rect 159822 195800 159878 195809
rect 159822 195735 159878 195744
rect 153934 194712 153990 194721
rect 153934 194647 153990 194656
rect 155222 194712 155278 194721
rect 155222 194647 155278 194656
rect 153948 194018 153976 194647
rect 153502 193990 153976 194018
rect 151634 193624 151690 193633
rect 151634 193559 151690 193568
rect 153290 193624 153346 193633
rect 153290 193559 153346 193568
rect 151648 191146 151676 193559
rect 151636 191140 151688 191146
rect 151636 191082 151688 191088
rect 149794 190632 149850 190641
rect 149638 190590 149794 190618
rect 149794 190567 149850 190576
rect 164252 189394 164280 199378
rect 166078 196208 166134 196217
rect 166078 196143 166134 196152
rect 165436 195696 165488 195702
rect 165436 195638 165488 195644
rect 165448 190454 165476 195638
rect 165448 190426 165568 190454
rect 164252 189366 164634 189394
rect 144642 186960 144698 186969
rect 144578 186918 144642 186946
rect 144642 186895 144698 186904
rect 162136 184198 162426 184226
rect 136836 182974 137494 183002
rect 136836 180334 136864 182974
rect 137020 182022 137494 182050
rect 136824 180328 136876 180334
rect 136824 180270 136876 180276
rect 136640 180124 136692 180130
rect 136640 180066 136692 180072
rect 136652 178838 136680 180066
rect 122840 178832 122892 178838
rect 122840 178774 122892 178780
rect 136640 178832 136692 178838
rect 136640 178774 136692 178780
rect 122852 151814 122880 178774
rect 137020 178702 137048 182022
rect 141252 180130 141280 181084
rect 162136 180946 162164 184198
rect 162124 180940 162176 180946
rect 162124 180882 162176 180888
rect 144460 180736 144512 180742
rect 146116 180736 146168 180742
rect 144460 180678 144512 180684
rect 146114 180704 146116 180713
rect 146168 180704 146170 180713
rect 144472 180676 144500 180678
rect 146114 180639 146170 180648
rect 161664 180600 161716 180606
rect 161664 180542 161716 180548
rect 141240 180124 141292 180130
rect 141240 180066 141292 180072
rect 137112 179982 137494 180010
rect 137008 178696 137060 178702
rect 137008 178638 137060 178644
rect 137112 177342 137140 179982
rect 143540 179648 143592 179654
rect 143540 179590 143592 179596
rect 143552 179588 143580 179590
rect 137204 179030 137494 179058
rect 124220 177336 124272 177342
rect 124220 177278 124272 177284
rect 137100 177336 137152 177342
rect 137100 177278 137152 177284
rect 124232 151814 124260 177278
rect 137204 176050 137232 179030
rect 140792 177886 140820 179452
rect 148046 179072 148102 179081
rect 147982 179030 148046 179058
rect 148046 179007 148102 179016
rect 142666 178800 142722 178809
rect 142666 178735 142722 178744
rect 144184 178696 144236 178702
rect 144184 178638 144236 178644
rect 140780 177880 140832 177886
rect 140780 177822 140832 177828
rect 141608 177880 141660 177886
rect 141608 177822 141660 177828
rect 137296 176990 137494 177018
rect 125600 176044 125652 176050
rect 125600 175986 125652 175992
rect 137192 176044 137244 176050
rect 137192 175986 137244 175992
rect 125612 151814 125640 175986
rect 137296 175982 137324 176990
rect 137388 176038 137494 176066
rect 128360 175976 128412 175982
rect 128360 175918 128412 175924
rect 137284 175976 137336 175982
rect 137284 175918 137336 175924
rect 126980 173188 127032 173194
rect 126980 173130 127032 173136
rect 126992 151814 127020 173130
rect 128372 151814 128400 175918
rect 135258 174040 135314 174049
rect 135258 173975 135314 173984
rect 135272 173942 135300 173975
rect 133880 173936 133932 173942
rect 133880 173878 133932 173884
rect 135260 173936 135312 173942
rect 135260 173878 135312 173884
rect 131120 173256 131172 173262
rect 131120 173198 131172 173204
rect 130384 165640 130436 165646
rect 130384 165582 130436 165588
rect 122852 151786 122972 151814
rect 124232 151786 124536 151814
rect 125612 151786 126100 151814
rect 126992 151786 127664 151814
rect 128372 151786 129228 151814
rect 122944 139890 122972 151786
rect 124508 139890 124536 151786
rect 126072 139890 126100 151786
rect 127636 139890 127664 151786
rect 129200 139890 129228 151786
rect 130396 142866 130424 165582
rect 130384 142860 130436 142866
rect 130384 142802 130436 142808
rect 131132 139890 131160 173198
rect 132500 172236 132552 172242
rect 132500 172178 132552 172184
rect 132512 139890 132540 172178
rect 133892 139890 133920 173878
rect 137388 173262 137416 176038
rect 137376 173256 137428 173262
rect 137376 173198 137428 173204
rect 135260 172440 135312 172446
rect 135260 172382 135312 172388
rect 135272 151814 135300 172382
rect 137480 172242 137508 174964
rect 137834 174040 137890 174049
rect 137890 173998 137954 174026
rect 137834 173975 137890 173984
rect 141620 173874 141648 177822
rect 142066 176760 142122 176769
rect 142066 176695 142122 176704
rect 140780 173868 140832 173874
rect 140780 173810 140832 173816
rect 141608 173868 141660 173874
rect 141608 173810 141660 173816
rect 138952 172446 138980 173740
rect 139412 173726 139978 173754
rect 138940 172440 138992 172446
rect 138940 172382 138992 172388
rect 137468 172236 137520 172242
rect 137468 172178 137520 172184
rect 138020 171964 138072 171970
rect 138020 171906 138072 171912
rect 138032 151814 138060 171906
rect 135272 151786 135484 151814
rect 138032 151786 138612 151814
rect 135456 139890 135484 151786
rect 137744 143200 137796 143206
rect 137744 143142 137796 143148
rect 137756 139890 137784 143142
rect 122944 139862 123372 139890
rect 124508 139862 124936 139890
rect 126072 139862 126500 139890
rect 127636 139862 128064 139890
rect 129200 139862 129628 139890
rect 131132 139862 131192 139890
rect 132512 139862 132756 139890
rect 133892 139862 134320 139890
rect 135456 139862 135884 139890
rect 137448 139862 137784 139890
rect 138584 139890 138612 151786
rect 139412 143206 139440 173726
rect 140792 173194 140820 173810
rect 140780 173188 140832 173194
rect 140780 173130 140832 173136
rect 140976 171970 141004 173740
rect 141068 173726 142002 173754
rect 140964 171964 141016 171970
rect 140964 171906 141016 171912
rect 141068 161474 141096 173726
rect 142080 171193 142108 176695
rect 144196 174593 144224 178638
rect 161676 178566 161704 180542
rect 159088 178560 159140 178566
rect 159088 178502 159140 178508
rect 161664 178560 161716 178566
rect 161664 178502 161716 178508
rect 159100 176254 159128 178502
rect 159088 176248 159140 176254
rect 159088 176190 159140 176196
rect 159088 175636 159140 175642
rect 159088 175578 159140 175584
rect 144182 174584 144238 174593
rect 144182 174519 144238 174528
rect 156050 174584 156106 174593
rect 156050 174519 156106 174528
rect 145654 173904 145710 173913
rect 145710 173862 145958 173890
rect 145654 173839 145710 173848
rect 142618 173768 142674 173777
rect 148690 173768 148746 173777
rect 142674 173726 142922 173754
rect 142618 173703 142674 173712
rect 142066 171184 142122 171193
rect 142066 171119 142122 171128
rect 142066 171048 142122 171057
rect 142066 170983 142122 170992
rect 142080 161537 142108 170983
rect 140976 161446 141096 161474
rect 142066 161528 142122 161537
rect 142066 161463 142122 161472
rect 139400 143200 139452 143206
rect 139400 143142 139452 143148
rect 140976 142154 141004 161446
rect 143538 142488 143594 142497
rect 143538 142423 143594 142432
rect 140700 142126 141004 142154
rect 142066 142216 142122 142225
rect 142066 142151 142122 142160
rect 140700 139890 140728 142126
rect 138584 139862 139012 139890
rect 140576 139862 140728 139890
rect 142080 139890 142108 142151
rect 143552 139890 143580 142423
rect 144932 139890 144960 173740
rect 146772 173726 146970 173754
rect 146772 173641 146800 173726
rect 148746 173726 148994 173754
rect 149072 173726 149914 173754
rect 150452 173726 150926 173754
rect 152476 173726 152950 173754
rect 148690 173703 148746 173712
rect 146758 173632 146814 173641
rect 146758 173567 146814 173576
rect 146482 143440 146538 143449
rect 146482 143375 146538 143384
rect 146496 139890 146524 143375
rect 148046 143304 148102 143313
rect 148046 143239 148102 143248
rect 148060 139890 148088 143239
rect 149072 142186 149100 173726
rect 149610 143168 149666 143177
rect 149610 143103 149666 143112
rect 149060 142180 149112 142186
rect 149060 142122 149112 142128
rect 149624 139890 149652 143103
rect 150452 142934 150480 173726
rect 152476 161474 152504 173726
rect 151832 161446 152504 161474
rect 151832 143546 151860 161446
rect 151820 143540 151872 143546
rect 151820 143482 151872 143488
rect 151174 143032 151230 143041
rect 151174 142967 151230 142976
rect 151358 143032 151414 143041
rect 151358 142967 151414 142976
rect 150440 142928 150492 142934
rect 150440 142870 150492 142876
rect 151188 139890 151216 142967
rect 151372 142633 151400 142967
rect 154580 142928 154632 142934
rect 154580 142870 154632 142876
rect 151358 142624 151414 142633
rect 151358 142559 151414 142568
rect 152740 142180 152792 142186
rect 152740 142122 152792 142128
rect 152752 139890 152780 142122
rect 154592 139890 154620 142870
rect 156064 139890 156092 174519
rect 157432 143540 157484 143546
rect 157432 143482 157484 143488
rect 157444 139890 157472 143482
rect 159100 139890 159128 175578
rect 165540 175030 165568 190426
rect 165528 175024 165580 175030
rect 165528 174966 165580 174972
rect 163136 174752 163188 174758
rect 163136 174694 163188 174700
rect 165528 174752 165580 174758
rect 165528 174694 165580 174700
rect 160020 171086 160048 173740
rect 160008 171080 160060 171086
rect 160008 171022 160060 171028
rect 162860 164824 162912 164830
rect 162860 164766 162912 164772
rect 162768 143132 162820 143138
rect 162768 143074 162820 143080
rect 160558 143032 160614 143041
rect 160558 142967 160614 142976
rect 160572 139890 160600 142967
rect 162780 139890 162808 143074
rect 162872 143002 162900 164766
rect 162860 142996 162912 143002
rect 162860 142938 162912 142944
rect 163148 142866 163176 174694
rect 163608 173726 163990 173754
rect 164252 173726 165002 173754
rect 163608 164830 163636 173726
rect 163872 171080 163924 171086
rect 163872 171022 163924 171028
rect 163884 165578 163912 171022
rect 163872 165572 163924 165578
rect 163872 165514 163924 165520
rect 163596 164824 163648 164830
rect 163596 164766 163648 164772
rect 164056 143472 164108 143478
rect 164056 143414 164108 143420
rect 163136 142860 163188 142866
rect 163136 142802 163188 142808
rect 164068 140162 164096 143414
rect 164252 142934 164280 173726
rect 164330 166424 164386 166433
rect 164330 166359 164386 166368
rect 164344 151814 164372 166359
rect 165540 161474 165568 174694
rect 165448 161446 165568 161474
rect 164344 151786 165200 151814
rect 164240 142928 164292 142934
rect 164240 142870 164292 142876
rect 142080 139862 142140 139890
rect 143552 139862 143704 139890
rect 144932 139862 145268 139890
rect 146496 139862 146832 139890
rect 148060 139862 148396 139890
rect 149624 139862 149960 139890
rect 151188 139862 151524 139890
rect 152752 139862 153088 139890
rect 154592 139862 154652 139890
rect 156064 139862 156216 139890
rect 157444 139862 157780 139890
rect 159100 139862 159344 139890
rect 160572 139862 160908 139890
rect 162472 139862 162808 139890
rect 164022 140134 164096 140162
rect 164022 139876 164050 140134
rect 165172 139890 165200 151786
rect 165448 150958 165476 161446
rect 165436 150952 165488 150958
rect 165436 150894 165488 150900
rect 166092 143478 166120 196143
rect 166170 196072 166226 196081
rect 166170 196007 166226 196016
rect 166080 143472 166132 143478
rect 166080 143414 166132 143420
rect 166184 143138 166212 196007
rect 166264 195968 166316 195974
rect 166264 195910 166316 195916
rect 166276 178294 166304 195910
rect 166264 178288 166316 178294
rect 166264 178230 166316 178236
rect 167644 178288 167696 178294
rect 167644 178230 167696 178236
rect 166998 166288 167054 166297
rect 166998 166223 167054 166232
rect 166264 165572 166316 165578
rect 166264 165514 166316 165520
rect 166276 147354 166304 165514
rect 166264 147348 166316 147354
rect 166264 147290 166316 147296
rect 166172 143132 166224 143138
rect 166172 143074 166224 143080
rect 167012 139890 167040 166223
rect 167656 165578 167684 178230
rect 179420 174140 179472 174146
rect 179420 174082 179472 174088
rect 167644 165572 167696 165578
rect 167644 165514 167696 165520
rect 169024 165572 169076 165578
rect 169024 165514 169076 165520
rect 167736 150952 167788 150958
rect 167736 150894 167788 150900
rect 167748 143546 167776 150894
rect 168380 147348 168432 147354
rect 168380 147290 168432 147296
rect 167736 143540 167788 143546
rect 167736 143482 167788 143488
rect 168392 139890 168420 147290
rect 169036 146946 169064 165514
rect 178684 149116 178736 149122
rect 178684 149058 178736 149064
rect 169024 146940 169076 146946
rect 169024 146882 169076 146888
rect 175188 146940 175240 146946
rect 175188 146882 175240 146888
rect 175200 146282 175228 146882
rect 175200 146254 175320 146282
rect 175292 143614 175320 146254
rect 175280 143608 175332 143614
rect 175280 143550 175332 143556
rect 169944 143540 169996 143546
rect 169944 143482 169996 143488
rect 178224 143540 178276 143546
rect 178224 143482 178276 143488
rect 169956 139890 169984 143482
rect 174636 142996 174688 143002
rect 174636 142938 174688 142944
rect 171506 142896 171562 142905
rect 171506 142831 171562 142840
rect 171520 139890 171548 142831
rect 173070 142760 173126 142769
rect 173070 142695 173126 142704
rect 173084 139890 173112 142695
rect 174648 139890 174676 142938
rect 176200 142928 176252 142934
rect 176200 142870 176252 142876
rect 176212 139890 176240 142870
rect 178040 142860 178092 142866
rect 178040 142802 178092 142808
rect 178052 139890 178080 142802
rect 165172 139862 165600 139890
rect 167012 139862 167164 139890
rect 168392 139862 168728 139890
rect 169956 139862 170292 139890
rect 171520 139862 171856 139890
rect 173084 139862 173420 139890
rect 174648 139862 174984 139890
rect 176212 139862 176548 139890
rect 178052 139862 178112 139890
rect 122104 139528 122156 139534
rect 122104 139470 122156 139476
rect 178236 139398 178264 143482
rect 178224 139392 178276 139398
rect 178224 139334 178276 139340
rect 178696 139330 178724 149058
rect 178684 139324 178736 139330
rect 178684 139266 178736 139272
rect 179432 126177 179460 174082
rect 179418 126168 179474 126177
rect 179418 126103 179474 126112
rect 179524 116657 179552 220050
rect 179604 160744 179656 160750
rect 179604 160686 179656 160692
rect 179510 116648 179566 116657
rect 179510 116583 179566 116592
rect 179616 113937 179644 160686
rect 180156 139392 180208 139398
rect 180156 139334 180208 139340
rect 179694 130520 179750 130529
rect 179694 130455 179750 130464
rect 179602 113928 179658 113937
rect 179602 113863 179658 113872
rect 121090 108352 121146 108361
rect 121090 108287 121146 108296
rect 120998 107672 121054 107681
rect 120998 107607 121054 107616
rect 120908 79552 120960 79558
rect 120908 79494 120960 79500
rect 120264 79416 120316 79422
rect 120264 79358 120316 79364
rect 119344 79212 119396 79218
rect 119344 79154 119396 79160
rect 120906 77616 120962 77625
rect 120906 77551 120962 77560
rect 120920 76634 120948 77551
rect 120908 76628 120960 76634
rect 120908 76570 120960 76576
rect 120908 76152 120960 76158
rect 120908 76094 120960 76100
rect 120724 75540 120776 75546
rect 120724 75482 120776 75488
rect 120080 64932 120132 64938
rect 120080 64874 120132 64880
rect 118424 46912 118476 46918
rect 118424 46854 118476 46860
rect 120092 16574 120120 64874
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 120092 16546 120672 16574
rect 113824 13116 113876 13122
rect 113824 13058 113876 13064
rect 114006 10432 114062 10441
rect 114006 10367 114062 10376
rect 114020 480 114048 10367
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 117320 10396 117372 10402
rect 117320 10338 117372 10344
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 10338
rect 117688 3936 117740 3942
rect 117688 3878 117740 3884
rect 117700 3602 117728 3878
rect 117688 3596 117740 3602
rect 117688 3538 117740 3544
rect 119896 3596 119948 3602
rect 119896 3538 119948 3544
rect 118792 3188 118844 3194
rect 118792 3130 118844 3136
rect 118804 480 118832 3130
rect 119908 480 119936 3538
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 120736 3194 120764 75482
rect 120816 74996 120868 75002
rect 120816 74938 120868 74944
rect 120828 21418 120856 74938
rect 120920 47598 120948 76094
rect 121104 75274 121132 108287
rect 178960 82136 179012 82142
rect 178960 82078 179012 82084
rect 121828 80640 121880 80646
rect 121828 80582 121880 80588
rect 174452 80640 174504 80646
rect 174452 80582 174504 80588
rect 174544 80640 174596 80646
rect 178040 80640 178092 80646
rect 174544 80582 174596 80588
rect 174910 80608 174966 80617
rect 121840 77246 121868 80582
rect 125140 80368 125192 80374
rect 125140 80310 125192 80316
rect 124772 80300 124824 80306
rect 124772 80242 124824 80248
rect 123482 80200 123538 80209
rect 123482 80135 123538 80144
rect 123576 80164 123628 80170
rect 123300 80096 123352 80102
rect 123300 80038 123352 80044
rect 123208 80028 123260 80034
rect 123208 79970 123260 79976
rect 122196 79960 122248 79966
rect 122196 79902 122248 79908
rect 121828 77240 121880 77246
rect 121828 77182 121880 77188
rect 122104 76900 122156 76906
rect 122104 76842 122156 76848
rect 121092 75268 121144 75274
rect 121092 75210 121144 75216
rect 121460 71324 121512 71330
rect 121460 71266 121512 71272
rect 120908 47592 120960 47598
rect 120908 47534 120960 47540
rect 120816 21412 120868 21418
rect 120816 21354 120868 21360
rect 121472 16574 121500 71266
rect 121472 16546 122052 16574
rect 122024 3482 122052 16546
rect 122116 3602 122144 76842
rect 122208 3942 122236 79902
rect 122378 79792 122434 79801
rect 122378 79727 122434 79736
rect 123024 79756 123076 79762
rect 122288 76084 122340 76090
rect 122288 76026 122340 76032
rect 122300 9042 122328 76026
rect 122392 36582 122420 79727
rect 123024 79698 123076 79704
rect 122932 77444 122984 77450
rect 122932 77386 122984 77392
rect 122840 74044 122892 74050
rect 122840 73986 122892 73992
rect 122380 36576 122432 36582
rect 122380 36518 122432 36524
rect 122852 16574 122880 73986
rect 122944 73953 122972 77386
rect 123036 75070 123064 79698
rect 123116 78192 123168 78198
rect 123116 78134 123168 78140
rect 123128 77586 123156 78134
rect 123116 77580 123168 77586
rect 123116 77522 123168 77528
rect 123024 75064 123076 75070
rect 123024 75006 123076 75012
rect 122930 73944 122986 73953
rect 122930 73879 122986 73888
rect 123220 72554 123248 79970
rect 123312 78169 123340 80038
rect 123298 78160 123354 78169
rect 123298 78095 123354 78104
rect 123208 72548 123260 72554
rect 123208 72490 123260 72496
rect 122852 16546 123064 16574
rect 122288 9036 122340 9042
rect 122288 8978 122340 8984
rect 122196 3936 122248 3942
rect 122196 3878 122248 3884
rect 122104 3596 122156 3602
rect 122104 3538 122156 3544
rect 122024 3454 122328 3482
rect 120724 3188 120776 3194
rect 120724 3130 120776 3136
rect 122300 480 122328 3454
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 123496 3874 123524 80135
rect 123576 80106 123628 80112
rect 123484 3868 123536 3874
rect 123484 3810 123536 3816
rect 123588 3738 123616 80106
rect 124126 78024 124182 78033
rect 124126 77959 124182 77968
rect 123668 77920 123720 77926
rect 123668 77862 123720 77868
rect 123680 64938 123708 77862
rect 123944 77240 123996 77246
rect 123944 77182 123996 77188
rect 123956 75750 123984 77182
rect 123944 75744 123996 75750
rect 123944 75686 123996 75692
rect 123668 64932 123720 64938
rect 123668 64874 123720 64880
rect 124140 14618 124168 77959
rect 124784 73710 124812 80242
rect 124956 80232 125008 80238
rect 124956 80174 125008 80180
rect 124864 79824 124916 79830
rect 124864 79766 124916 79772
rect 124772 73704 124824 73710
rect 124772 73646 124824 73652
rect 124220 20052 124272 20058
rect 124220 19994 124272 20000
rect 124232 16574 124260 19994
rect 124232 16546 124720 16574
rect 124128 14612 124180 14618
rect 124128 14554 124180 14560
rect 123576 3732 123628 3738
rect 123576 3674 123628 3680
rect 124692 480 124720 16546
rect 124876 3534 124904 79766
rect 124968 75342 124996 80174
rect 125152 79626 125180 80310
rect 174464 80170 174492 80582
rect 174556 80345 174584 80582
rect 174728 80572 174780 80578
rect 178040 80582 178092 80588
rect 174910 80543 174966 80552
rect 174728 80514 174780 80520
rect 174636 80436 174688 80442
rect 174636 80378 174688 80384
rect 174542 80336 174598 80345
rect 174542 80271 174598 80280
rect 174452 80164 174504 80170
rect 174452 80106 174504 80112
rect 125244 80022 125580 80050
rect 125140 79620 125192 79626
rect 125140 79562 125192 79568
rect 125048 78600 125100 78606
rect 125048 78542 125100 78548
rect 125060 75818 125088 78542
rect 125140 77716 125192 77722
rect 125140 77658 125192 77664
rect 125048 75812 125100 75818
rect 125048 75754 125100 75760
rect 124956 75336 125008 75342
rect 124956 75278 125008 75284
rect 125048 73364 125100 73370
rect 125048 73306 125100 73312
rect 124956 72276 125008 72282
rect 124956 72218 125008 72224
rect 124864 3528 124916 3534
rect 124864 3470 124916 3476
rect 124968 3466 124996 72218
rect 125060 3670 125088 73306
rect 125152 10470 125180 77658
rect 125244 73846 125272 80022
rect 125658 79830 125686 80036
rect 125750 79966 125778 80036
rect 125842 79971 125870 80036
rect 125738 79960 125790 79966
rect 125738 79902 125790 79908
rect 125828 79962 125884 79971
rect 125828 79897 125884 79906
rect 125646 79824 125698 79830
rect 125934 79778 125962 80036
rect 125646 79766 125698 79772
rect 125888 79750 125962 79778
rect 125600 79552 125652 79558
rect 125600 79494 125652 79500
rect 125692 79552 125744 79558
rect 125692 79494 125744 79500
rect 125612 78946 125640 79494
rect 125600 78940 125652 78946
rect 125600 78882 125652 78888
rect 125416 78464 125468 78470
rect 125416 78406 125468 78412
rect 125232 73840 125284 73846
rect 125232 73782 125284 73788
rect 125232 73704 125284 73710
rect 125232 73646 125284 73652
rect 125244 43450 125272 73646
rect 125428 73522 125456 78406
rect 125508 75812 125560 75818
rect 125508 75754 125560 75760
rect 125600 75812 125652 75818
rect 125600 75754 125652 75760
rect 125336 73494 125456 73522
rect 125336 55894 125364 73494
rect 125520 70394 125548 75754
rect 125612 75274 125640 75754
rect 125600 75268 125652 75274
rect 125600 75210 125652 75216
rect 125704 72282 125732 79494
rect 125888 75954 125916 79750
rect 126026 79642 126054 80036
rect 126118 79966 126146 80036
rect 126106 79960 126158 79966
rect 126106 79902 126158 79908
rect 126210 79898 126238 80036
rect 126302 79966 126330 80036
rect 126290 79960 126342 79966
rect 126290 79902 126342 79908
rect 126198 79892 126250 79898
rect 126198 79834 126250 79840
rect 126394 79812 126422 80036
rect 126486 79966 126514 80036
rect 126474 79960 126526 79966
rect 126474 79902 126526 79908
rect 126578 79898 126606 80036
rect 126670 79898 126698 80036
rect 126762 79966 126790 80036
rect 126750 79960 126802 79966
rect 126750 79902 126802 79908
rect 126566 79892 126618 79898
rect 126566 79834 126618 79840
rect 126658 79892 126710 79898
rect 126658 79834 126710 79840
rect 126348 79784 126422 79812
rect 126244 79756 126296 79762
rect 126244 79698 126296 79704
rect 126026 79614 126100 79642
rect 125968 79144 126020 79150
rect 125968 79086 126020 79092
rect 125876 75948 125928 75954
rect 125876 75890 125928 75896
rect 125876 75676 125928 75682
rect 125876 75618 125928 75624
rect 125692 72276 125744 72282
rect 125692 72218 125744 72224
rect 125428 70366 125548 70394
rect 125428 60042 125456 70366
rect 125416 60036 125468 60042
rect 125416 59978 125468 59984
rect 125324 55888 125376 55894
rect 125324 55830 125376 55836
rect 125232 43444 125284 43450
rect 125232 43386 125284 43392
rect 125140 10464 125192 10470
rect 125140 10406 125192 10412
rect 125888 7614 125916 75618
rect 125980 8974 126008 79086
rect 126072 77897 126100 79614
rect 126152 79620 126204 79626
rect 126152 79562 126204 79568
rect 126164 78674 126192 79562
rect 126256 79150 126284 79698
rect 126348 79626 126376 79784
rect 126520 79756 126572 79762
rect 126520 79698 126572 79704
rect 126336 79620 126388 79626
rect 126336 79562 126388 79568
rect 126336 79484 126388 79490
rect 126336 79426 126388 79432
rect 126244 79144 126296 79150
rect 126244 79086 126296 79092
rect 126164 78646 126284 78674
rect 126150 78296 126206 78305
rect 126150 78231 126206 78240
rect 126164 78062 126192 78231
rect 126152 78056 126204 78062
rect 126152 77998 126204 78004
rect 126058 77888 126114 77897
rect 126058 77823 126114 77832
rect 126256 75970 126284 78646
rect 126348 76498 126376 79426
rect 126336 76492 126388 76498
rect 126336 76434 126388 76440
rect 126060 75948 126112 75954
rect 126256 75942 126376 75970
rect 126060 75890 126112 75896
rect 125968 8968 126020 8974
rect 125968 8910 126020 8916
rect 125876 7608 125928 7614
rect 125876 7550 125928 7556
rect 126072 4826 126100 75890
rect 126244 74316 126296 74322
rect 126244 74258 126296 74264
rect 126152 73092 126204 73098
rect 126152 73034 126204 73040
rect 126164 66910 126192 73034
rect 126152 66904 126204 66910
rect 126152 66846 126204 66852
rect 126060 4820 126112 4826
rect 126060 4762 126112 4768
rect 125876 4140 125928 4146
rect 125876 4082 125928 4088
rect 125048 3664 125100 3670
rect 125048 3606 125100 3612
rect 124956 3460 125008 3466
rect 124956 3402 125008 3408
rect 125888 480 125916 4082
rect 126256 3806 126284 74258
rect 126348 4894 126376 75942
rect 126532 6186 126560 79698
rect 126612 79688 126664 79694
rect 126854 79676 126882 80036
rect 126808 79648 126882 79676
rect 126808 79642 126836 79648
rect 126612 79630 126664 79636
rect 126624 72486 126652 79630
rect 126716 79614 126836 79642
rect 126716 73098 126744 79614
rect 126946 79608 126974 80036
rect 127038 79801 127066 80036
rect 127130 79830 127158 80036
rect 127222 79966 127250 80036
rect 127210 79960 127262 79966
rect 127210 79902 127262 79908
rect 127314 79898 127342 80036
rect 127406 79898 127434 80036
rect 127498 79966 127526 80036
rect 127486 79960 127538 79966
rect 127486 79902 127538 79908
rect 127302 79892 127354 79898
rect 127302 79834 127354 79840
rect 127394 79892 127446 79898
rect 127394 79834 127446 79840
rect 127118 79824 127170 79830
rect 127024 79792 127080 79801
rect 127118 79766 127170 79772
rect 127024 79727 127080 79736
rect 127440 79756 127492 79762
rect 127590 79744 127618 80036
rect 127682 79778 127710 80036
rect 127774 79898 127802 80036
rect 127762 79892 127814 79898
rect 127762 79834 127814 79840
rect 127866 79812 127894 80036
rect 127958 79966 127986 80036
rect 127946 79960 127998 79966
rect 128050 79937 128078 80036
rect 128142 79966 128170 80036
rect 128130 79960 128182 79966
rect 127946 79902 127998 79908
rect 128036 79928 128092 79937
rect 128130 79902 128182 79908
rect 128036 79863 128092 79872
rect 127866 79784 127940 79812
rect 127682 79750 127756 79778
rect 127440 79698 127492 79704
rect 127544 79716 127618 79744
rect 127728 79744 127756 79750
rect 127728 79716 127848 79744
rect 127072 79688 127124 79694
rect 127072 79630 127124 79636
rect 127348 79688 127400 79694
rect 127348 79630 127400 79636
rect 126900 79580 126974 79608
rect 126796 79552 126848 79558
rect 126796 79494 126848 79500
rect 126808 76537 126836 79494
rect 126794 76528 126850 76537
rect 126794 76463 126850 76472
rect 126900 75682 126928 79580
rect 126980 79280 127032 79286
rect 126980 79222 127032 79228
rect 126992 79082 127020 79222
rect 126980 79076 127032 79082
rect 126980 79018 127032 79024
rect 126980 77104 127032 77110
rect 126980 77046 127032 77052
rect 126888 75676 126940 75682
rect 126888 75618 126940 75624
rect 126704 73092 126756 73098
rect 126704 73034 126756 73040
rect 126612 72480 126664 72486
rect 126612 72422 126664 72428
rect 126992 71126 127020 77046
rect 127084 75993 127112 79630
rect 127256 79144 127308 79150
rect 127256 79086 127308 79092
rect 127268 78946 127296 79086
rect 127256 78940 127308 78946
rect 127256 78882 127308 78888
rect 127360 76090 127388 79630
rect 127452 78266 127480 79698
rect 127440 78260 127492 78266
rect 127440 78202 127492 78208
rect 127544 76106 127572 79716
rect 127624 79620 127676 79626
rect 127624 79562 127676 79568
rect 127716 79620 127768 79626
rect 127716 79562 127768 79568
rect 127348 76084 127400 76090
rect 127348 76026 127400 76032
rect 127452 76078 127572 76106
rect 127070 75984 127126 75993
rect 127070 75919 127126 75928
rect 127256 75948 127308 75954
rect 127256 75890 127308 75896
rect 126980 71120 127032 71126
rect 126980 71062 127032 71068
rect 127268 35222 127296 75890
rect 127348 75676 127400 75682
rect 127348 75618 127400 75624
rect 127256 35216 127308 35222
rect 127256 35158 127308 35164
rect 127360 7750 127388 75618
rect 127452 72622 127480 76078
rect 127440 72616 127492 72622
rect 127440 72558 127492 72564
rect 127440 72480 127492 72486
rect 127440 72422 127492 72428
rect 127452 69698 127480 72422
rect 127636 71774 127664 79562
rect 127728 75954 127756 79562
rect 127716 75948 127768 75954
rect 127716 75890 127768 75896
rect 127820 75682 127848 79716
rect 127912 75954 127940 79784
rect 128084 79756 128136 79762
rect 128234 79744 128262 80036
rect 128326 79898 128354 80036
rect 128418 79937 128446 80036
rect 128510 79966 128538 80036
rect 128498 79960 128550 79966
rect 128404 79928 128460 79937
rect 128314 79892 128366 79898
rect 128498 79902 128550 79908
rect 128404 79863 128460 79872
rect 128314 79834 128366 79840
rect 128084 79698 128136 79704
rect 128188 79716 128262 79744
rect 128360 79756 128412 79762
rect 127992 79688 128044 79694
rect 127992 79630 128044 79636
rect 127900 75948 127952 75954
rect 127900 75890 127952 75896
rect 127808 75676 127860 75682
rect 127808 75618 127860 75624
rect 128004 73370 128032 79630
rect 127992 73364 128044 73370
rect 127992 73306 128044 73312
rect 128096 72486 128124 79698
rect 128084 72480 128136 72486
rect 128084 72422 128136 72428
rect 127544 71746 127664 71774
rect 127440 69692 127492 69698
rect 127440 69634 127492 69640
rect 127348 7744 127400 7750
rect 127348 7686 127400 7692
rect 127544 7682 127572 71746
rect 128188 70394 128216 79716
rect 128360 79698 128412 79704
rect 128452 79756 128504 79762
rect 128602 79744 128630 80036
rect 128694 79937 128722 80036
rect 128786 79966 128814 80036
rect 128774 79960 128826 79966
rect 128680 79928 128736 79937
rect 128774 79902 128826 79908
rect 128878 79898 128906 80036
rect 128680 79863 128736 79872
rect 128866 79892 128918 79898
rect 128866 79834 128918 79840
rect 128452 79698 128504 79704
rect 128556 79716 128630 79744
rect 128728 79756 128780 79762
rect 128268 79620 128320 79626
rect 128268 79562 128320 79568
rect 128280 76158 128308 79562
rect 128268 76152 128320 76158
rect 128268 76094 128320 76100
rect 128268 75948 128320 75954
rect 128268 75890 128320 75896
rect 128280 71058 128308 75890
rect 128372 75206 128400 79698
rect 128360 75200 128412 75206
rect 128360 75142 128412 75148
rect 128464 74225 128492 79698
rect 128556 75002 128584 79716
rect 128970 79744 128998 80036
rect 129062 79937 129090 80036
rect 129048 79928 129104 79937
rect 129154 79898 129182 80036
rect 129246 79966 129274 80036
rect 129234 79960 129286 79966
rect 129234 79902 129286 79908
rect 129048 79863 129104 79872
rect 129142 79892 129194 79898
rect 129142 79834 129194 79840
rect 129338 79778 129366 80036
rect 129430 79898 129458 80036
rect 129522 79971 129550 80036
rect 129508 79962 129564 79971
rect 129418 79892 129470 79898
rect 129508 79897 129564 79906
rect 129614 79898 129642 80036
rect 129706 79898 129734 80036
rect 129418 79834 129470 79840
rect 129602 79892 129654 79898
rect 129602 79834 129654 79840
rect 129694 79892 129746 79898
rect 129694 79834 129746 79840
rect 128728 79698 128780 79704
rect 128924 79716 128998 79744
rect 129188 79756 129240 79762
rect 128636 79212 128688 79218
rect 128636 79154 128688 79160
rect 128544 74996 128596 75002
rect 128544 74938 128596 74944
rect 128450 74216 128506 74225
rect 128450 74151 128506 74160
rect 128268 71052 128320 71058
rect 128268 70994 128320 71000
rect 128648 70394 128676 79154
rect 128740 78169 128768 79698
rect 128820 79552 128872 79558
rect 128820 79494 128872 79500
rect 128726 78160 128782 78169
rect 128726 78095 128782 78104
rect 128832 76242 128860 79494
rect 128924 79218 128952 79716
rect 129188 79698 129240 79704
rect 129292 79750 129366 79778
rect 129462 79792 129518 79801
rect 129096 79688 129148 79694
rect 129096 79630 129148 79636
rect 129004 79416 129056 79422
rect 129004 79358 129056 79364
rect 129016 79218 129044 79358
rect 128912 79212 128964 79218
rect 128912 79154 128964 79160
rect 129004 79212 129056 79218
rect 129004 79154 129056 79160
rect 129108 77432 129136 79630
rect 127820 70366 128216 70394
rect 128556 70366 128676 70394
rect 128740 76214 128860 76242
rect 128924 77404 129136 77432
rect 127820 9110 127848 70366
rect 128556 10334 128584 70366
rect 128544 10328 128596 10334
rect 128544 10270 128596 10276
rect 127808 9104 127860 9110
rect 127808 9046 127860 9052
rect 127532 7676 127584 7682
rect 127532 7618 127584 7624
rect 126520 6180 126572 6186
rect 126520 6122 126572 6128
rect 128740 5030 128768 76214
rect 128924 76106 128952 77404
rect 129004 77308 129056 77314
rect 129004 77250 129056 77256
rect 128832 76078 128952 76106
rect 128832 69766 128860 76078
rect 128912 75948 128964 75954
rect 128912 75890 128964 75896
rect 128820 69760 128872 69766
rect 128820 69702 128872 69708
rect 128728 5024 128780 5030
rect 128728 4966 128780 4972
rect 128924 4962 128952 75890
rect 129016 6390 129044 77250
rect 129200 77110 129228 79698
rect 129188 77104 129240 77110
rect 129188 77046 129240 77052
rect 129188 76968 129240 76974
rect 129188 76910 129240 76916
rect 129094 74488 129150 74497
rect 129094 74423 129150 74432
rect 129004 6384 129056 6390
rect 129004 6326 129056 6332
rect 128912 4956 128964 4962
rect 128912 4898 128964 4904
rect 126336 4888 126388 4894
rect 126336 4830 126388 4836
rect 128176 3868 128228 3874
rect 128176 3810 128228 3816
rect 126244 3800 126296 3806
rect 126244 3742 126296 3748
rect 126980 3528 127032 3534
rect 126980 3470 127032 3476
rect 126992 480 127020 3470
rect 128188 480 128216 3810
rect 129108 3534 129136 74423
rect 129200 22846 129228 76910
rect 129292 75954 129320 79750
rect 129462 79727 129518 79736
rect 129556 79756 129608 79762
rect 129280 75948 129332 75954
rect 129280 75890 129332 75896
rect 129476 73914 129504 79727
rect 129798 79744 129826 80036
rect 129890 79830 129918 80036
rect 129982 79937 130010 80036
rect 129968 79928 130024 79937
rect 129968 79863 130024 79872
rect 129878 79824 129930 79830
rect 129878 79766 129930 79772
rect 129556 79698 129608 79704
rect 129752 79716 129826 79744
rect 129568 79558 129596 79698
rect 129556 79552 129608 79558
rect 129556 79494 129608 79500
rect 129648 79552 129700 79558
rect 129648 79494 129700 79500
rect 129556 79416 129608 79422
rect 129556 79358 129608 79364
rect 129568 74322 129596 79358
rect 129660 77353 129688 79494
rect 129752 77994 129780 79716
rect 130074 79676 130102 80036
rect 130166 79744 130194 80036
rect 130258 79812 130286 80036
rect 130350 79966 130378 80036
rect 130338 79960 130390 79966
rect 130338 79902 130390 79908
rect 130258 79801 130332 79812
rect 130258 79792 130346 79801
rect 130258 79784 130290 79792
rect 130166 79716 130240 79744
rect 130290 79727 130346 79736
rect 129922 79656 129978 79665
rect 130074 79648 130148 79676
rect 129922 79591 129978 79600
rect 129740 77988 129792 77994
rect 129740 77930 129792 77936
rect 129646 77344 129702 77353
rect 129646 77279 129702 77288
rect 129936 76974 129964 79591
rect 130016 79552 130068 79558
rect 130016 79494 130068 79500
rect 129924 76968 129976 76974
rect 129924 76910 129976 76916
rect 130028 76888 130056 79494
rect 130120 77450 130148 79648
rect 130108 77444 130160 77450
rect 130108 77386 130160 77392
rect 130028 76860 130148 76888
rect 129924 76832 129976 76838
rect 129924 76774 129976 76780
rect 129740 75608 129792 75614
rect 129740 75550 129792 75556
rect 129556 74316 129608 74322
rect 129556 74258 129608 74264
rect 129464 73908 129516 73914
rect 129464 73850 129516 73856
rect 129188 22840 129240 22846
rect 129188 22782 129240 22788
rect 129752 16574 129780 75550
rect 129936 70394 129964 76774
rect 130120 76616 130148 76860
rect 130212 76838 130240 79716
rect 130442 79676 130470 80036
rect 130534 79966 130562 80036
rect 130626 79966 130654 80036
rect 130522 79960 130574 79966
rect 130522 79902 130574 79908
rect 130614 79960 130666 79966
rect 130718 79937 130746 80036
rect 130614 79902 130666 79908
rect 130704 79928 130760 79937
rect 130704 79863 130760 79872
rect 130810 79744 130838 80036
rect 130902 79830 130930 80036
rect 130994 79966 131022 80036
rect 130982 79960 131034 79966
rect 130982 79902 131034 79908
rect 130890 79824 130942 79830
rect 131086 79778 131114 80036
rect 131178 79971 131206 80036
rect 131164 79962 131220 79971
rect 131270 79966 131298 80036
rect 131362 79966 131390 80036
rect 131454 79966 131482 80036
rect 131164 79897 131220 79906
rect 131258 79960 131310 79966
rect 131258 79902 131310 79908
rect 131350 79960 131402 79966
rect 131350 79902 131402 79908
rect 131442 79960 131494 79966
rect 131546 79937 131574 80036
rect 131442 79902 131494 79908
rect 131532 79928 131588 79937
rect 131532 79863 131588 79872
rect 131258 79824 131310 79830
rect 130890 79766 130942 79772
rect 131040 79750 131114 79778
rect 131256 79792 131258 79801
rect 131310 79792 131312 79801
rect 131040 79744 131068 79750
rect 130718 79716 130838 79744
rect 130994 79716 131068 79744
rect 131256 79727 131312 79736
rect 131638 79744 131666 80036
rect 131730 79971 131758 80036
rect 131716 79962 131772 79971
rect 131716 79897 131772 79906
rect 131822 79744 131850 80036
rect 131638 79716 131712 79744
rect 130290 79656 130346 79665
rect 130442 79648 130516 79676
rect 130290 79591 130346 79600
rect 130200 76832 130252 76838
rect 130200 76774 130252 76780
rect 129844 70366 129964 70394
rect 130028 76588 130148 76616
rect 130200 76628 130252 76634
rect 129844 68338 129872 70366
rect 129832 68332 129884 68338
rect 129832 68274 129884 68280
rect 129752 16546 129964 16574
rect 129096 3528 129148 3534
rect 129096 3470 129148 3476
rect 129936 3482 129964 16546
rect 130028 6322 130056 76588
rect 130200 76570 130252 76576
rect 130108 76492 130160 76498
rect 130108 76434 130160 76440
rect 130120 22914 130148 76434
rect 130212 66978 130240 76570
rect 130200 66972 130252 66978
rect 130200 66914 130252 66920
rect 130108 22908 130160 22914
rect 130108 22850 130160 22856
rect 130016 6316 130068 6322
rect 130016 6258 130068 6264
rect 130304 5098 130332 79591
rect 130488 6254 130516 79648
rect 130718 79642 130746 79716
rect 130994 79676 131022 79716
rect 130672 79614 130746 79642
rect 130948 79648 131022 79676
rect 131304 79688 131356 79694
rect 131210 79656 131266 79665
rect 130568 79416 130620 79422
rect 130568 79358 130620 79364
rect 130580 76634 130608 79358
rect 130568 76628 130620 76634
rect 130568 76570 130620 76576
rect 130672 76498 130700 79614
rect 130752 79552 130804 79558
rect 130752 79494 130804 79500
rect 130660 76492 130712 76498
rect 130660 76434 130712 76440
rect 130764 73154 130792 79494
rect 130844 79484 130896 79490
rect 130844 79426 130896 79432
rect 130856 79218 130884 79426
rect 130844 79212 130896 79218
rect 130844 79154 130896 79160
rect 130948 75410 130976 79648
rect 131304 79630 131356 79636
rect 131578 79656 131634 79665
rect 131210 79591 131266 79600
rect 131028 79212 131080 79218
rect 131028 79154 131080 79160
rect 131040 77586 131068 79154
rect 131120 77852 131172 77858
rect 131120 77794 131172 77800
rect 131028 77580 131080 77586
rect 131028 77522 131080 77528
rect 131132 75546 131160 77794
rect 131120 75540 131172 75546
rect 131120 75482 131172 75488
rect 130936 75404 130988 75410
rect 130936 75346 130988 75352
rect 130672 73126 130792 73154
rect 130672 72690 130700 73126
rect 130660 72684 130712 72690
rect 130660 72626 130712 72632
rect 131224 69834 131252 79591
rect 131316 77217 131344 79630
rect 131396 79620 131448 79626
rect 131578 79591 131634 79600
rect 131396 79562 131448 79568
rect 131408 77353 131436 79562
rect 131488 79552 131540 79558
rect 131488 79494 131540 79500
rect 131394 77344 131450 77353
rect 131394 77279 131450 77288
rect 131396 77240 131448 77246
rect 131302 77208 131358 77217
rect 131396 77182 131448 77188
rect 131302 77143 131358 77152
rect 131304 77104 131356 77110
rect 131304 77046 131356 77052
rect 131212 69828 131264 69834
rect 131212 69770 131264 69776
rect 131316 6526 131344 77046
rect 131408 44878 131436 77182
rect 131500 69902 131528 79494
rect 131488 69896 131540 69902
rect 131488 69838 131540 69844
rect 131396 44872 131448 44878
rect 131396 44814 131448 44820
rect 131304 6520 131356 6526
rect 131304 6462 131356 6468
rect 130476 6248 130528 6254
rect 130476 6190 130528 6196
rect 131592 5166 131620 79591
rect 131684 77314 131712 79716
rect 131776 79716 131850 79744
rect 131914 79744 131942 80036
rect 132006 79966 132034 80036
rect 131994 79960 132046 79966
rect 131994 79902 132046 79908
rect 132098 79898 132126 80036
rect 132190 79903 132218 80036
rect 132086 79892 132138 79898
rect 132086 79834 132138 79840
rect 132176 79894 132232 79903
rect 132176 79829 132232 79838
rect 132282 79830 132310 80036
rect 132374 79898 132402 80036
rect 132466 79966 132494 80036
rect 132454 79960 132506 79966
rect 132558 79937 132586 80036
rect 132650 79966 132678 80036
rect 132742 79966 132770 80036
rect 132834 79971 132862 80036
rect 132638 79960 132690 79966
rect 132454 79902 132506 79908
rect 132544 79928 132600 79937
rect 132362 79892 132414 79898
rect 132638 79902 132690 79908
rect 132730 79960 132782 79966
rect 132730 79902 132782 79908
rect 132820 79962 132876 79971
rect 132820 79897 132876 79906
rect 132544 79863 132600 79872
rect 132362 79834 132414 79840
rect 132270 79824 132322 79830
rect 132500 79824 132552 79830
rect 132270 79766 132322 79772
rect 132420 79772 132500 79778
rect 132420 79766 132552 79772
rect 132420 79750 132540 79766
rect 132592 79756 132644 79762
rect 131914 79716 131988 79744
rect 131672 77308 131724 77314
rect 131672 77250 131724 77256
rect 131776 70394 131804 79716
rect 131960 77246 131988 79716
rect 132224 79620 132276 79626
rect 132224 79562 132276 79568
rect 132132 79552 132184 79558
rect 132132 79494 132184 79500
rect 131948 77240 132000 77246
rect 131948 77182 132000 77188
rect 132144 77110 132172 79494
rect 132132 77104 132184 77110
rect 132132 77046 132184 77052
rect 132236 70394 132264 79562
rect 132316 79552 132368 79558
rect 132316 79494 132368 79500
rect 132328 76702 132356 79494
rect 132420 76770 132448 79750
rect 132592 79698 132644 79704
rect 132498 79656 132554 79665
rect 132498 79591 132554 79600
rect 132512 78130 132540 79591
rect 132604 78441 132632 79698
rect 132776 79688 132828 79694
rect 132926 79676 132954 80036
rect 133018 79830 133046 80036
rect 133110 79898 133138 80036
rect 133202 79966 133230 80036
rect 133190 79960 133242 79966
rect 133190 79902 133242 79908
rect 133098 79892 133150 79898
rect 133098 79834 133150 79840
rect 133006 79824 133058 79830
rect 133006 79766 133058 79772
rect 133052 79688 133104 79694
rect 132926 79648 133000 79676
rect 132776 79630 132828 79636
rect 132684 79416 132736 79422
rect 132684 79358 132736 79364
rect 132696 78946 132724 79358
rect 132684 78940 132736 78946
rect 132684 78882 132736 78888
rect 132684 78736 132736 78742
rect 132684 78678 132736 78684
rect 132590 78432 132646 78441
rect 132590 78367 132646 78376
rect 132500 78124 132552 78130
rect 132500 78066 132552 78072
rect 132408 76764 132460 76770
rect 132408 76706 132460 76712
rect 132316 76696 132368 76702
rect 132696 76673 132724 78678
rect 132788 78169 132816 79630
rect 132868 79552 132920 79558
rect 132868 79494 132920 79500
rect 132774 78160 132830 78169
rect 132774 78095 132830 78104
rect 132776 78056 132828 78062
rect 132776 77998 132828 78004
rect 132316 76638 132368 76644
rect 132682 76664 132738 76673
rect 132682 76599 132738 76608
rect 132684 71732 132736 71738
rect 132684 71674 132736 71680
rect 131684 70366 131804 70394
rect 132144 70366 132264 70394
rect 131684 6458 131712 70366
rect 131762 69592 131818 69601
rect 131762 69527 131818 69536
rect 131672 6452 131724 6458
rect 131672 6394 131724 6400
rect 131580 5160 131632 5166
rect 131580 5102 131632 5108
rect 130292 5092 130344 5098
rect 130292 5034 130344 5040
rect 131776 3874 131804 69527
rect 132144 68406 132172 70366
rect 132132 68400 132184 68406
rect 132132 68342 132184 68348
rect 132696 6914 132724 71674
rect 132788 19990 132816 77998
rect 132880 77926 132908 79494
rect 132972 78742 133000 79648
rect 133052 79630 133104 79636
rect 133294 79642 133322 80036
rect 133386 79778 133414 80036
rect 133478 79966 133506 80036
rect 133570 79966 133598 80036
rect 133662 79971 133690 80036
rect 133466 79960 133518 79966
rect 133466 79902 133518 79908
rect 133558 79960 133610 79966
rect 133558 79902 133610 79908
rect 133648 79962 133704 79971
rect 133754 79966 133782 80036
rect 133846 79966 133874 80036
rect 133938 79966 133966 80036
rect 134030 79971 134058 80036
rect 133648 79897 133704 79906
rect 133742 79960 133794 79966
rect 133742 79902 133794 79908
rect 133834 79960 133886 79966
rect 133834 79902 133886 79908
rect 133926 79960 133978 79966
rect 133926 79902 133978 79908
rect 134016 79962 134072 79971
rect 134122 79966 134150 80036
rect 134214 79971 134242 80036
rect 134016 79897 134072 79906
rect 134110 79960 134162 79966
rect 134110 79902 134162 79908
rect 134200 79962 134256 79971
rect 134306 79966 134334 80036
rect 134398 79966 134426 80036
rect 134490 79966 134518 80036
rect 134200 79897 134256 79906
rect 134294 79960 134346 79966
rect 134294 79902 134346 79908
rect 134386 79960 134438 79966
rect 134386 79902 134438 79908
rect 134478 79960 134530 79966
rect 134478 79902 134530 79908
rect 133880 79824 133932 79830
rect 133386 79750 133644 79778
rect 133880 79766 133932 79772
rect 134064 79824 134116 79830
rect 134064 79766 134116 79772
rect 134156 79824 134208 79830
rect 134582 79812 134610 80036
rect 134674 79971 134702 80036
rect 134660 79962 134716 79971
rect 134766 79966 134794 80036
rect 134858 79966 134886 80036
rect 134950 79966 134978 80036
rect 134660 79897 134716 79906
rect 134754 79960 134806 79966
rect 134754 79902 134806 79908
rect 134846 79960 134898 79966
rect 134846 79902 134898 79908
rect 134938 79960 134990 79966
rect 134938 79902 134990 79908
rect 134156 79766 134208 79772
rect 134338 79792 134394 79801
rect 133420 79688 133472 79694
rect 132960 78736 133012 78742
rect 132960 78678 133012 78684
rect 133064 78470 133092 79630
rect 133144 79620 133196 79626
rect 133294 79614 133368 79642
rect 133420 79630 133472 79636
rect 133512 79688 133564 79694
rect 133512 79630 133564 79636
rect 133144 79562 133196 79568
rect 133052 78464 133104 78470
rect 133052 78406 133104 78412
rect 132960 78328 133012 78334
rect 132960 78270 133012 78276
rect 132868 77920 132920 77926
rect 132868 77862 132920 77868
rect 132866 77208 132922 77217
rect 132866 77143 132922 77152
rect 132880 24138 132908 77143
rect 132868 24132 132920 24138
rect 132868 24074 132920 24080
rect 132776 19984 132828 19990
rect 132776 19926 132828 19932
rect 132972 7886 133000 78270
rect 132960 7880 133012 7886
rect 132960 7822 133012 7828
rect 133156 7818 133184 79562
rect 133234 78296 133290 78305
rect 133234 78231 133290 78240
rect 133248 73982 133276 78231
rect 133340 78062 133368 79614
rect 133432 78674 133460 79630
rect 133420 78668 133472 78674
rect 133420 78610 133472 78616
rect 133524 78554 133552 79630
rect 133616 78810 133644 79750
rect 133696 79756 133748 79762
rect 133696 79698 133748 79704
rect 133604 78804 133656 78810
rect 133604 78746 133656 78752
rect 133602 78704 133658 78713
rect 133602 78639 133658 78648
rect 133432 78526 133552 78554
rect 133328 78056 133380 78062
rect 133328 77998 133380 78004
rect 133328 77920 133380 77926
rect 133328 77862 133380 77868
rect 133236 73976 133288 73982
rect 133236 73918 133288 73924
rect 133340 71194 133368 77862
rect 133432 72826 133460 78526
rect 133512 78464 133564 78470
rect 133512 78406 133564 78412
rect 133420 72820 133472 72826
rect 133420 72762 133472 72768
rect 133524 71262 133552 78406
rect 133616 72758 133644 78639
rect 133708 78402 133736 79698
rect 133788 79552 133840 79558
rect 133788 79494 133840 79500
rect 133696 78396 133748 78402
rect 133696 78338 133748 78344
rect 133696 78260 133748 78266
rect 133696 78202 133748 78208
rect 133604 72752 133656 72758
rect 133604 72694 133656 72700
rect 133512 71256 133564 71262
rect 133512 71198 133564 71204
rect 133328 71188 133380 71194
rect 133328 71130 133380 71136
rect 133708 70394 133736 78202
rect 133800 75682 133828 79494
rect 133892 77858 133920 79766
rect 133972 79756 134024 79762
rect 133972 79698 134024 79704
rect 133984 79665 134012 79698
rect 133970 79656 134026 79665
rect 133970 79591 134026 79600
rect 133972 79484 134024 79490
rect 133972 79426 134024 79432
rect 133880 77852 133932 77858
rect 133880 77794 133932 77800
rect 133880 77444 133932 77450
rect 133880 77386 133932 77392
rect 133788 75676 133840 75682
rect 133788 75618 133840 75624
rect 133708 70366 133828 70394
rect 133144 7812 133196 7818
rect 133144 7754 133196 7760
rect 132696 6886 133000 6914
rect 131764 3868 131816 3874
rect 131764 3810 131816 3816
rect 131764 3732 131816 3738
rect 131764 3674 131816 3680
rect 129936 3454 130608 3482
rect 129372 3188 129424 3194
rect 129372 3130 129424 3136
rect 129384 480 129412 3130
rect 130580 480 130608 3454
rect 131776 480 131804 3674
rect 132972 480 133000 6886
rect 133800 3670 133828 70366
rect 133788 3664 133840 3670
rect 133788 3606 133840 3612
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133892 354 133920 77386
rect 133984 70394 134012 79426
rect 134076 77722 134104 79766
rect 134064 77716 134116 77722
rect 134064 77658 134116 77664
rect 134168 76809 134196 79766
rect 134248 79756 134300 79762
rect 134338 79727 134394 79736
rect 134444 79784 134610 79812
rect 134800 79824 134852 79830
rect 134660 79792 134716 79801
rect 134248 79698 134300 79704
rect 134260 78713 134288 79698
rect 134352 79218 134380 79727
rect 134340 79212 134392 79218
rect 134340 79154 134392 79160
rect 134444 79064 134472 79784
rect 134352 79036 134472 79064
rect 134628 79736 134660 79744
rect 135042 79812 135070 80036
rect 135134 79835 135162 80036
rect 134996 79784 135070 79812
rect 135120 79826 135176 79835
rect 134996 79778 135024 79784
rect 134800 79766 134852 79772
rect 134628 79727 134716 79736
rect 134628 79716 134702 79727
rect 134246 78704 134302 78713
rect 134246 78639 134302 78648
rect 134154 76800 134210 76809
rect 134154 76735 134210 76744
rect 134352 70394 134380 79036
rect 134628 78962 134656 79716
rect 134708 79552 134760 79558
rect 134708 79494 134760 79500
rect 133984 70366 134104 70394
rect 134076 20058 134104 70366
rect 134260 70366 134380 70394
rect 134444 78934 134656 78962
rect 134260 68474 134288 70366
rect 134248 68468 134300 68474
rect 134248 68410 134300 68416
rect 134064 20052 134116 20058
rect 134064 19994 134116 20000
rect 134444 10402 134472 78934
rect 134720 77994 134748 79494
rect 134708 77988 134760 77994
rect 134708 77930 134760 77936
rect 134524 77716 134576 77722
rect 134524 77658 134576 77664
rect 134432 10396 134484 10402
rect 134432 10338 134484 10344
rect 134536 4146 134564 77658
rect 134812 76906 134840 79766
rect 134950 79750 135024 79778
rect 135120 79761 135176 79770
rect 134950 79642 134978 79750
rect 135226 79676 135254 80036
rect 135318 79744 135346 80036
rect 135410 79966 135438 80036
rect 135502 79971 135530 80036
rect 135398 79960 135450 79966
rect 135398 79902 135450 79908
rect 135488 79962 135544 79971
rect 135594 79966 135622 80036
rect 135488 79897 135544 79906
rect 135582 79960 135634 79966
rect 135582 79902 135634 79908
rect 135444 79824 135496 79830
rect 135686 79778 135714 80036
rect 135778 79966 135806 80036
rect 135766 79960 135818 79966
rect 135766 79902 135818 79908
rect 135870 79812 135898 80036
rect 135962 79937 135990 80036
rect 135948 79928 136004 79937
rect 136054 79898 136082 80036
rect 136146 79966 136174 80036
rect 136238 79966 136266 80036
rect 136134 79960 136186 79966
rect 136134 79902 136186 79908
rect 136226 79960 136278 79966
rect 136226 79902 136278 79908
rect 135948 79863 136004 79872
rect 136042 79892 136094 79898
rect 136042 79834 136094 79840
rect 136330 79812 136358 80036
rect 135444 79766 135496 79772
rect 135318 79716 135392 79744
rect 134904 79614 134978 79642
rect 135074 79656 135130 79665
rect 134800 76900 134852 76906
rect 134800 76842 134852 76848
rect 134616 74520 134668 74526
rect 134616 74462 134668 74468
rect 134524 4140 134576 4146
rect 134524 4082 134576 4088
rect 134628 3194 134656 74462
rect 134904 71330 134932 79614
rect 135074 79591 135130 79600
rect 135180 79648 135254 79676
rect 135088 74050 135116 79591
rect 135180 79490 135208 79648
rect 135260 79552 135312 79558
rect 135260 79494 135312 79500
rect 135168 79484 135220 79490
rect 135168 79426 135220 79432
rect 135168 79212 135220 79218
rect 135168 79154 135220 79160
rect 135180 79014 135208 79154
rect 135168 79008 135220 79014
rect 135168 78950 135220 78956
rect 135272 77353 135300 79494
rect 135364 77722 135392 79716
rect 135352 77716 135404 77722
rect 135352 77658 135404 77664
rect 135258 77344 135314 77353
rect 135456 77294 135484 79766
rect 135594 79750 135714 79778
rect 135824 79784 135898 79812
rect 136284 79784 136358 79812
rect 135594 79676 135622 79750
rect 135824 79676 135852 79784
rect 135258 77279 135314 77288
rect 135364 77266 135484 77294
rect 135548 79648 135622 79676
rect 135732 79648 135852 79676
rect 135904 79688 135956 79694
rect 135364 74526 135392 77266
rect 135444 75676 135496 75682
rect 135444 75618 135496 75624
rect 135352 74520 135404 74526
rect 135352 74462 135404 74468
rect 135076 74044 135128 74050
rect 135076 73986 135128 73992
rect 134892 71324 134944 71330
rect 134892 71266 134944 71272
rect 135260 3596 135312 3602
rect 135260 3538 135312 3544
rect 134616 3188 134668 3194
rect 134616 3130 134668 3136
rect 135272 480 135300 3538
rect 135456 3126 135484 75618
rect 135548 75614 135576 79648
rect 135628 79552 135680 79558
rect 135628 79494 135680 79500
rect 135536 75608 135588 75614
rect 135536 75550 135588 75556
rect 135536 75472 135588 75478
rect 135536 75414 135588 75420
rect 135548 3194 135576 75414
rect 135640 3738 135668 79494
rect 135732 77314 135760 79648
rect 136180 79688 136232 79694
rect 135904 79630 135956 79636
rect 135994 79656 136050 79665
rect 135720 77308 135772 77314
rect 135720 77250 135772 77256
rect 135812 75268 135864 75274
rect 135812 75210 135864 75216
rect 135720 75200 135772 75206
rect 135720 75142 135772 75148
rect 135732 21690 135760 75142
rect 135824 53038 135852 75210
rect 135812 53032 135864 53038
rect 135812 52974 135864 52980
rect 135720 21684 135772 21690
rect 135720 21626 135772 21632
rect 135916 16574 135944 79630
rect 136180 79630 136232 79636
rect 135994 79591 136050 79600
rect 136088 79620 136140 79626
rect 136008 77450 136036 79591
rect 136088 79562 136140 79568
rect 135996 77444 136048 77450
rect 135996 77386 136048 77392
rect 135996 77308 136048 77314
rect 135996 77250 136048 77256
rect 136008 71738 136036 77250
rect 135996 71732 136048 71738
rect 135996 71674 136048 71680
rect 135916 16546 136036 16574
rect 135628 3732 135680 3738
rect 135628 3674 135680 3680
rect 136008 3482 136036 16546
rect 136100 3602 136128 79562
rect 136192 75478 136220 79630
rect 136284 75682 136312 79784
rect 136422 79744 136450 80036
rect 136376 79716 136450 79744
rect 136272 75676 136324 75682
rect 136272 75618 136324 75624
rect 136180 75472 136232 75478
rect 136180 75414 136232 75420
rect 136376 75206 136404 79716
rect 136514 79506 136542 80036
rect 136606 79971 136634 80036
rect 136592 79962 136648 79971
rect 136592 79897 136648 79906
rect 136698 79744 136726 80036
rect 136468 79478 136542 79506
rect 136652 79716 136726 79744
rect 136468 75274 136496 79478
rect 136548 78600 136600 78606
rect 136548 78542 136600 78548
rect 136560 77897 136588 78542
rect 136546 77888 136602 77897
rect 136546 77823 136602 77832
rect 136652 77654 136680 79716
rect 136790 79676 136818 80036
rect 136744 79648 136818 79676
rect 136882 79676 136910 80036
rect 136974 79744 137002 80036
rect 137066 79937 137094 80036
rect 137052 79928 137108 79937
rect 137158 79898 137186 80036
rect 137052 79863 137108 79872
rect 137146 79892 137198 79898
rect 137146 79834 137198 79840
rect 137250 79778 137278 80036
rect 137204 79750 137278 79778
rect 136974 79716 137048 79744
rect 136882 79648 136956 79676
rect 136640 77648 136692 77654
rect 136640 77590 136692 77596
rect 136456 75268 136508 75274
rect 136456 75210 136508 75216
rect 136744 75206 136772 79648
rect 136928 78826 136956 79648
rect 136836 78798 136956 78826
rect 136836 75274 136864 78798
rect 136914 78704 136970 78713
rect 136914 78639 136970 78648
rect 136824 75268 136876 75274
rect 136824 75210 136876 75216
rect 136364 75200 136416 75206
rect 136364 75142 136416 75148
rect 136732 75200 136784 75206
rect 136732 75142 136784 75148
rect 136824 75132 136876 75138
rect 136824 75074 136876 75080
rect 136732 75064 136784 75070
rect 136732 75006 136784 75012
rect 136744 4826 136772 75006
rect 136836 11762 136864 75074
rect 136928 21486 136956 78639
rect 137020 78266 137048 79716
rect 137100 79688 137152 79694
rect 137100 79630 137152 79636
rect 137008 78260 137060 78266
rect 137008 78202 137060 78208
rect 137112 75342 137140 79630
rect 137100 75336 137152 75342
rect 137100 75278 137152 75284
rect 137008 75268 137060 75274
rect 137008 75210 137060 75216
rect 137020 46850 137048 75210
rect 137100 75200 137152 75206
rect 137100 75142 137152 75148
rect 137112 59362 137140 75142
rect 137204 69018 137232 79750
rect 137342 79676 137370 80036
rect 137434 79898 137462 80036
rect 137422 79892 137474 79898
rect 137422 79834 137474 79840
rect 137526 79778 137554 80036
rect 137618 79898 137646 80036
rect 137606 79892 137658 79898
rect 137606 79834 137658 79840
rect 137710 79778 137738 80036
rect 137480 79750 137554 79778
rect 137664 79750 137738 79778
rect 137802 79778 137830 80036
rect 137894 79966 137922 80036
rect 137986 79971 138014 80036
rect 137882 79960 137934 79966
rect 137882 79902 137934 79908
rect 137972 79962 138028 79971
rect 137972 79897 138028 79906
rect 137928 79824 137980 79830
rect 137926 79792 137928 79801
rect 137980 79792 137982 79801
rect 137802 79750 137876 79778
rect 137342 79648 137416 79676
rect 137284 79348 137336 79354
rect 137284 79290 137336 79296
rect 137296 79150 137324 79290
rect 137284 79144 137336 79150
rect 137284 79086 137336 79092
rect 137282 77888 137338 77897
rect 137282 77823 137338 77832
rect 137296 77625 137324 77823
rect 137282 77616 137338 77625
rect 137282 77551 137338 77560
rect 137284 75336 137336 75342
rect 137284 75278 137336 75284
rect 137296 70446 137324 75278
rect 137284 70440 137336 70446
rect 137284 70382 137336 70388
rect 137388 70394 137416 79648
rect 137480 75138 137508 79750
rect 137560 79688 137612 79694
rect 137560 79630 137612 79636
rect 137572 76566 137600 79630
rect 137664 77926 137692 79750
rect 137652 77920 137704 77926
rect 137652 77862 137704 77868
rect 137848 77294 137876 79750
rect 138078 79744 138106 80036
rect 138170 79937 138198 80036
rect 138156 79928 138212 79937
rect 138262 79898 138290 80036
rect 138156 79863 138212 79872
rect 138250 79892 138302 79898
rect 138250 79834 138302 79840
rect 138354 79778 138382 80036
rect 137926 79727 137982 79736
rect 138032 79716 138106 79744
rect 138204 79756 138256 79762
rect 137928 79688 137980 79694
rect 137928 79630 137980 79636
rect 137756 77266 137876 77294
rect 137560 76560 137612 76566
rect 137560 76502 137612 76508
rect 137468 75132 137520 75138
rect 137468 75074 137520 75080
rect 137756 75070 137784 77266
rect 137744 75064 137796 75070
rect 137744 75006 137796 75012
rect 137940 74322 137968 79630
rect 138032 78810 138060 79716
rect 138204 79698 138256 79704
rect 138308 79750 138382 79778
rect 138020 78804 138072 78810
rect 138020 78746 138072 78752
rect 138112 78804 138164 78810
rect 138112 78746 138164 78752
rect 138018 78704 138074 78713
rect 138018 78639 138074 78648
rect 138032 75342 138060 78639
rect 138020 75336 138072 75342
rect 138020 75278 138072 75284
rect 138020 75200 138072 75206
rect 138020 75142 138072 75148
rect 137928 74316 137980 74322
rect 137928 74258 137980 74264
rect 137388 70366 137968 70394
rect 137192 69012 137244 69018
rect 137192 68954 137244 68960
rect 137100 59356 137152 59362
rect 137100 59298 137152 59304
rect 137008 46844 137060 46850
rect 137008 46786 137060 46792
rect 136916 21480 136968 21486
rect 136916 21422 136968 21428
rect 136824 11756 136876 11762
rect 136824 11698 136876 11704
rect 137940 4894 137968 70366
rect 138032 5030 138060 75142
rect 138124 10334 138152 78746
rect 138216 75138 138244 79698
rect 138308 78305 138336 79750
rect 138446 79676 138474 80036
rect 138538 79966 138566 80036
rect 138526 79960 138578 79966
rect 138630 79937 138658 80036
rect 138526 79902 138578 79908
rect 138616 79928 138672 79937
rect 138616 79863 138672 79872
rect 138722 79830 138750 80036
rect 138814 79971 138842 80036
rect 138800 79962 138856 79971
rect 138906 79966 138934 80036
rect 138998 79966 139026 80036
rect 139090 79966 139118 80036
rect 138800 79897 138856 79906
rect 138894 79960 138946 79966
rect 138894 79902 138946 79908
rect 138986 79960 139038 79966
rect 138986 79902 139038 79908
rect 139078 79960 139130 79966
rect 139078 79902 139130 79908
rect 138710 79824 138762 79830
rect 138570 79792 138626 79801
rect 138710 79766 138762 79772
rect 138848 79824 138900 79830
rect 139182 79801 139210 80036
rect 139274 79812 139302 80036
rect 139366 79937 139394 80036
rect 139352 79928 139408 79937
rect 139352 79863 139408 79872
rect 138848 79766 138900 79772
rect 139168 79792 139224 79801
rect 138570 79727 138626 79736
rect 138400 79648 138474 79676
rect 138400 78810 138428 79648
rect 138388 78804 138440 78810
rect 138388 78746 138440 78752
rect 138388 78668 138440 78674
rect 138388 78610 138440 78616
rect 138294 78296 138350 78305
rect 138294 78231 138350 78240
rect 138296 76900 138348 76906
rect 138296 76842 138348 76848
rect 138204 75132 138256 75138
rect 138204 75074 138256 75080
rect 138204 74996 138256 75002
rect 138204 74938 138256 74944
rect 138216 21622 138244 74938
rect 138308 46238 138336 76842
rect 138400 47598 138428 78610
rect 138584 76906 138612 79727
rect 138756 79688 138808 79694
rect 138756 79630 138808 79636
rect 138664 79620 138716 79626
rect 138664 79562 138716 79568
rect 138572 76900 138624 76906
rect 138572 76842 138624 76848
rect 138480 75336 138532 75342
rect 138480 75278 138532 75284
rect 138492 60722 138520 75278
rect 138676 75206 138704 79562
rect 138664 75200 138716 75206
rect 138664 75142 138716 75148
rect 138572 75132 138624 75138
rect 138572 75074 138624 75080
rect 138584 66230 138612 75074
rect 138768 75002 138796 79630
rect 138756 74996 138808 75002
rect 138756 74938 138808 74944
rect 138860 74534 138888 79766
rect 139274 79784 139348 79812
rect 139168 79727 139224 79736
rect 139216 79688 139268 79694
rect 139216 79630 139268 79636
rect 139032 79620 139084 79626
rect 139032 79562 139084 79568
rect 139044 78010 139072 79562
rect 139124 79416 139176 79422
rect 139124 79358 139176 79364
rect 139136 79082 139164 79358
rect 139124 79076 139176 79082
rect 139124 79018 139176 79024
rect 139228 78305 139256 79630
rect 139214 78296 139270 78305
rect 139214 78231 139270 78240
rect 139044 77982 139256 78010
rect 139124 77648 139176 77654
rect 139124 77590 139176 77596
rect 138676 74506 138888 74534
rect 138676 68882 138704 74506
rect 138756 70440 138808 70446
rect 139136 70394 139164 77590
rect 139228 74118 139256 77982
rect 139320 77178 139348 79784
rect 139458 79744 139486 80036
rect 139550 79903 139578 80036
rect 139536 79894 139592 79903
rect 139536 79829 139592 79838
rect 139642 79778 139670 80036
rect 139734 79898 139762 80036
rect 139722 79892 139774 79898
rect 139722 79834 139774 79840
rect 139826 79778 139854 80036
rect 139918 79966 139946 80036
rect 139906 79960 139958 79966
rect 139906 79902 139958 79908
rect 140010 79778 140038 80036
rect 140102 79898 140130 80036
rect 140194 79898 140222 80036
rect 140090 79892 140142 79898
rect 140090 79834 140142 79840
rect 140182 79892 140234 79898
rect 140182 79834 140234 79840
rect 140286 79778 140314 80036
rect 140378 79966 140406 80036
rect 140470 79966 140498 80036
rect 140366 79960 140418 79966
rect 140366 79902 140418 79908
rect 140458 79960 140510 79966
rect 140458 79902 140510 79908
rect 140562 79898 140590 80036
rect 140654 79898 140682 80036
rect 140550 79892 140602 79898
rect 140550 79834 140602 79840
rect 140642 79892 140694 79898
rect 140642 79834 140694 79840
rect 140746 79830 140774 80036
rect 140838 79971 140866 80036
rect 140824 79962 140880 79971
rect 140824 79897 140880 79906
rect 139642 79750 139716 79778
rect 139826 79750 139900 79778
rect 140010 79750 140084 79778
rect 139458 79716 139532 79744
rect 139398 79656 139454 79665
rect 139398 79591 139454 79600
rect 139308 77172 139360 77178
rect 139308 77114 139360 77120
rect 139412 75274 139440 79591
rect 139504 78538 139532 79716
rect 139584 79688 139636 79694
rect 139584 79630 139636 79636
rect 139492 78532 139544 78538
rect 139492 78474 139544 78480
rect 139492 77240 139544 77246
rect 139492 77182 139544 77188
rect 139400 75268 139452 75274
rect 139400 75210 139452 75216
rect 139400 75132 139452 75138
rect 139400 75074 139452 75080
rect 139216 74112 139268 74118
rect 139216 74054 139268 74060
rect 138756 70382 138808 70388
rect 138664 68876 138716 68882
rect 138664 68818 138716 68824
rect 138572 66224 138624 66230
rect 138572 66166 138624 66172
rect 138480 60716 138532 60722
rect 138480 60658 138532 60664
rect 138388 47592 138440 47598
rect 138388 47534 138440 47540
rect 138664 46844 138716 46850
rect 138664 46786 138716 46792
rect 138296 46232 138348 46238
rect 138296 46174 138348 46180
rect 138204 21616 138256 21622
rect 138204 21558 138256 21564
rect 138112 10328 138164 10334
rect 138112 10270 138164 10276
rect 138020 5024 138072 5030
rect 138020 4966 138072 4972
rect 137928 4888 137980 4894
rect 137928 4830 137980 4836
rect 136732 4820 136784 4826
rect 136732 4762 136784 4768
rect 138676 3806 138704 46786
rect 138664 3800 138716 3806
rect 138664 3742 138716 3748
rect 136088 3596 136140 3602
rect 136088 3538 136140 3544
rect 136008 3454 136496 3482
rect 135536 3188 135588 3194
rect 135536 3130 135588 3136
rect 135444 3120 135496 3126
rect 135444 3062 135496 3068
rect 136468 480 136496 3454
rect 138768 3262 138796 70382
rect 138952 70366 139164 70394
rect 138848 69012 138900 69018
rect 138848 68954 138900 68960
rect 138860 3330 138888 68954
rect 138952 4418 138980 70366
rect 139412 23050 139440 75074
rect 139504 42226 139532 77182
rect 139596 53310 139624 79630
rect 139688 59022 139716 79750
rect 139768 79688 139820 79694
rect 139768 79630 139820 79636
rect 139780 77994 139808 79630
rect 139768 77988 139820 77994
rect 139768 77930 139820 77936
rect 139768 75268 139820 75274
rect 139768 75210 139820 75216
rect 139780 60314 139808 75210
rect 139768 60308 139820 60314
rect 139768 60250 139820 60256
rect 139872 60246 139900 79750
rect 139952 79688 140004 79694
rect 139952 79630 140004 79636
rect 139964 78674 139992 79630
rect 139952 78668 140004 78674
rect 139952 78610 140004 78616
rect 139952 77308 140004 77314
rect 139952 77250 140004 77256
rect 139964 67182 139992 77250
rect 140056 70242 140084 79750
rect 140240 79750 140314 79778
rect 140412 79824 140464 79830
rect 140412 79766 140464 79772
rect 140734 79824 140786 79830
rect 140734 79766 140786 79772
rect 140930 79778 140958 80036
rect 141022 79898 141050 80036
rect 141114 79898 141142 80036
rect 141010 79892 141062 79898
rect 141010 79834 141062 79840
rect 141102 79892 141154 79898
rect 141102 79834 141154 79840
rect 140240 79744 140268 79750
rect 140194 79716 140268 79744
rect 140194 79642 140222 79716
rect 140318 79656 140374 79665
rect 140194 79614 140268 79642
rect 140136 79552 140188 79558
rect 140136 79494 140188 79500
rect 140148 77246 140176 79494
rect 140240 77314 140268 79614
rect 140318 79591 140320 79600
rect 140372 79591 140374 79600
rect 140320 79562 140372 79568
rect 140320 79484 140372 79490
rect 140320 79426 140372 79432
rect 140332 78810 140360 79426
rect 140320 78804 140372 78810
rect 140320 78746 140372 78752
rect 140320 78668 140372 78674
rect 140320 78610 140372 78616
rect 140228 77308 140280 77314
rect 140228 77250 140280 77256
rect 140136 77240 140188 77246
rect 140136 77182 140188 77188
rect 140332 75138 140360 78610
rect 140424 78130 140452 79766
rect 140504 79756 140556 79762
rect 140930 79750 141096 79778
rect 140504 79698 140556 79704
rect 140412 78124 140464 78130
rect 140412 78066 140464 78072
rect 140412 77920 140464 77926
rect 140412 77862 140464 77868
rect 140320 75132 140372 75138
rect 140320 75074 140372 75080
rect 140044 70236 140096 70242
rect 140044 70178 140096 70184
rect 140042 67552 140098 67561
rect 140042 67487 140098 67496
rect 139952 67176 140004 67182
rect 139952 67118 140004 67124
rect 139860 60240 139912 60246
rect 139860 60182 139912 60188
rect 139676 59016 139728 59022
rect 139676 58958 139728 58964
rect 139584 53304 139636 53310
rect 139584 53246 139636 53252
rect 139492 42220 139544 42226
rect 139492 42162 139544 42168
rect 139400 23044 139452 23050
rect 139400 22986 139452 22992
rect 139400 21684 139452 21690
rect 139400 21626 139452 21632
rect 139412 16574 139440 21626
rect 139412 16546 139624 16574
rect 138940 4412 138992 4418
rect 138940 4354 138992 4360
rect 138848 3324 138900 3330
rect 138848 3266 138900 3272
rect 138756 3256 138808 3262
rect 138756 3198 138808 3204
rect 137652 3188 137704 3194
rect 137652 3130 137704 3136
rect 137664 480 137692 3130
rect 138848 3120 138900 3126
rect 138848 3062 138900 3068
rect 138860 480 138888 3062
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 140056 3466 140084 67487
rect 140136 66224 140188 66230
rect 140136 66166 140188 66172
rect 140148 3602 140176 66166
rect 140228 59356 140280 59362
rect 140228 59298 140280 59304
rect 140240 3874 140268 59298
rect 140320 53032 140372 53038
rect 140320 52974 140372 52980
rect 140228 3868 140280 3874
rect 140228 3810 140280 3816
rect 140136 3596 140188 3602
rect 140136 3538 140188 3544
rect 140332 3534 140360 52974
rect 140424 11830 140452 77862
rect 140516 77761 140544 79698
rect 140596 79688 140648 79694
rect 140872 79688 140924 79694
rect 140596 79630 140648 79636
rect 140686 79656 140742 79665
rect 140502 77752 140558 77761
rect 140502 77687 140558 77696
rect 140608 77489 140636 79630
rect 140872 79630 140924 79636
rect 140686 79591 140742 79600
rect 140700 78470 140728 79591
rect 140780 79280 140832 79286
rect 140780 79222 140832 79228
rect 140792 79150 140820 79222
rect 140780 79144 140832 79150
rect 140780 79086 140832 79092
rect 140780 78804 140832 78810
rect 140780 78746 140832 78752
rect 140792 78713 140820 78746
rect 140778 78704 140834 78713
rect 140778 78639 140834 78648
rect 140688 78464 140740 78470
rect 140688 78406 140740 78412
rect 140780 78396 140832 78402
rect 140780 78338 140832 78344
rect 140594 77480 140650 77489
rect 140594 77415 140650 77424
rect 140596 77172 140648 77178
rect 140596 77114 140648 77120
rect 140608 71398 140636 77114
rect 140596 71392 140648 71398
rect 140596 71334 140648 71340
rect 140792 12374 140820 78338
rect 140884 78266 140912 79630
rect 140964 79620 141016 79626
rect 140964 79562 141016 79568
rect 140872 78260 140924 78266
rect 140872 78202 140924 78208
rect 140976 77976 141004 79562
rect 141068 78198 141096 79750
rect 141206 79744 141234 80036
rect 141298 79812 141326 80036
rect 141390 79966 141418 80036
rect 141378 79960 141430 79966
rect 141482 79937 141510 80036
rect 141378 79902 141430 79908
rect 141468 79928 141524 79937
rect 141574 79898 141602 80036
rect 141666 79966 141694 80036
rect 141758 79966 141786 80036
rect 141850 79966 141878 80036
rect 141654 79960 141706 79966
rect 141654 79902 141706 79908
rect 141746 79960 141798 79966
rect 141746 79902 141798 79908
rect 141838 79960 141890 79966
rect 141838 79902 141890 79908
rect 141468 79863 141524 79872
rect 141562 79892 141614 79898
rect 141562 79834 141614 79840
rect 141298 79784 141372 79812
rect 141206 79716 141280 79744
rect 141148 79416 141200 79422
rect 141148 79358 141200 79364
rect 141056 78192 141108 78198
rect 141056 78134 141108 78140
rect 141160 77976 141188 79358
rect 140884 77948 141004 77976
rect 141068 77948 141188 77976
rect 140884 18834 140912 77948
rect 140964 77852 141016 77858
rect 140964 77794 141016 77800
rect 140976 31414 141004 77794
rect 141068 46442 141096 77948
rect 141148 76492 141200 76498
rect 141148 76434 141200 76440
rect 141160 51882 141188 76434
rect 141252 57322 141280 79716
rect 141344 78402 141372 79784
rect 141514 79792 141570 79801
rect 141942 79778 141970 80036
rect 142034 79971 142062 80036
rect 142020 79962 142076 79971
rect 142020 79897 142076 79906
rect 142126 79812 142154 80036
rect 142218 79966 142246 80036
rect 142310 79966 142338 80036
rect 142402 79966 142430 80036
rect 142494 79971 142522 80036
rect 142206 79960 142258 79966
rect 142206 79902 142258 79908
rect 142298 79960 142350 79966
rect 142298 79902 142350 79908
rect 142390 79960 142442 79966
rect 142390 79902 142442 79908
rect 142480 79962 142536 79971
rect 142586 79966 142614 80036
rect 142678 79966 142706 80036
rect 142770 79971 142798 80036
rect 142480 79897 142536 79906
rect 142574 79960 142626 79966
rect 142574 79902 142626 79908
rect 142666 79960 142718 79966
rect 142666 79902 142718 79908
rect 142756 79962 142812 79971
rect 142756 79897 142812 79906
rect 142080 79801 142154 79812
rect 141514 79727 141570 79736
rect 141850 79750 141970 79778
rect 142066 79792 142154 79801
rect 141424 79688 141476 79694
rect 141424 79630 141476 79636
rect 141332 78396 141384 78402
rect 141332 78338 141384 78344
rect 141332 78260 141384 78266
rect 141332 78202 141384 78208
rect 141344 67114 141372 78202
rect 141436 68814 141464 79630
rect 141528 76498 141556 79727
rect 141850 79676 141878 79750
rect 142122 79784 142154 79792
rect 142436 79824 142488 79830
rect 142436 79766 142488 79772
rect 142528 79824 142580 79830
rect 142528 79766 142580 79772
rect 142620 79824 142672 79830
rect 142620 79766 142672 79772
rect 142710 79792 142766 79801
rect 142066 79727 142122 79736
rect 141976 79688 142028 79694
rect 141850 79648 141924 79676
rect 141700 79552 141752 79558
rect 141700 79494 141752 79500
rect 141712 77858 141740 79494
rect 141792 79484 141844 79490
rect 141792 79426 141844 79432
rect 141700 77852 141752 77858
rect 141700 77794 141752 77800
rect 141804 77586 141832 79426
rect 141792 77580 141844 77586
rect 141792 77522 141844 77528
rect 141516 76492 141568 76498
rect 141516 76434 141568 76440
rect 141896 70394 141924 79648
rect 142160 79688 142212 79694
rect 141976 79630 142028 79636
rect 142066 79656 142122 79665
rect 141988 74050 142016 79630
rect 142160 79630 142212 79636
rect 142066 79591 142122 79600
rect 142080 75914 142108 79591
rect 142172 76498 142200 79630
rect 142252 79620 142304 79626
rect 142252 79562 142304 79568
rect 142344 79620 142396 79626
rect 142344 79562 142396 79568
rect 142264 77178 142292 79562
rect 142252 77172 142304 77178
rect 142252 77114 142304 77120
rect 142356 76809 142384 79562
rect 142342 76800 142398 76809
rect 142252 76764 142304 76770
rect 142342 76735 142398 76744
rect 142252 76706 142304 76712
rect 142160 76492 142212 76498
rect 142160 76434 142212 76440
rect 142080 75886 142200 75914
rect 141976 74044 142028 74050
rect 141976 73986 142028 73992
rect 141528 70366 141924 70394
rect 141528 70174 141556 70366
rect 141516 70168 141568 70174
rect 141516 70110 141568 70116
rect 141424 68808 141476 68814
rect 141424 68750 141476 68756
rect 141332 67108 141384 67114
rect 141332 67050 141384 67056
rect 141240 57316 141292 57322
rect 141240 57258 141292 57264
rect 141148 51876 141200 51882
rect 141148 51818 141200 51824
rect 141056 46436 141108 46442
rect 141056 46378 141108 46384
rect 140964 31408 141016 31414
rect 140964 31350 141016 31356
rect 140872 18828 140924 18834
rect 140872 18770 140924 18776
rect 140780 12368 140832 12374
rect 140780 12310 140832 12316
rect 140412 11824 140464 11830
rect 140412 11766 140464 11772
rect 140320 3528 140372 3534
rect 140320 3470 140372 3476
rect 141240 3528 141292 3534
rect 141240 3470 141292 3476
rect 140044 3460 140096 3466
rect 140044 3402 140096 3408
rect 141252 480 141280 3470
rect 142172 3398 142200 75886
rect 142264 4146 142292 76706
rect 142344 76628 142396 76634
rect 142344 76570 142396 76576
rect 142356 24274 142384 76570
rect 142448 31346 142476 79766
rect 142540 45082 142568 79766
rect 142632 76650 142660 79766
rect 142862 79778 142890 80036
rect 142710 79727 142766 79736
rect 142816 79750 142890 79778
rect 142724 76770 142752 79727
rect 142712 76764 142764 76770
rect 142712 76706 142764 76712
rect 142632 76622 142752 76650
rect 142816 76634 142844 79750
rect 142954 79676 142982 80036
rect 143046 79812 143074 80036
rect 143138 79966 143166 80036
rect 143230 79966 143258 80036
rect 143126 79960 143178 79966
rect 143126 79902 143178 79908
rect 143218 79960 143270 79966
rect 143218 79902 143270 79908
rect 143172 79824 143224 79830
rect 143046 79784 143120 79812
rect 142954 79648 143028 79676
rect 142896 79348 142948 79354
rect 142896 79290 142948 79296
rect 142908 79150 142936 79290
rect 142896 79144 142948 79150
rect 142896 79086 142948 79092
rect 142620 76492 142672 76498
rect 142620 76434 142672 76440
rect 142632 47870 142660 76434
rect 142724 54738 142752 76622
rect 142804 76628 142856 76634
rect 142804 76570 142856 76576
rect 142896 74316 142948 74322
rect 142896 74258 142948 74264
rect 142712 54732 142764 54738
rect 142712 54674 142764 54680
rect 142620 47864 142672 47870
rect 142620 47806 142672 47812
rect 142528 45076 142580 45082
rect 142528 45018 142580 45024
rect 142436 31340 142488 31346
rect 142436 31282 142488 31288
rect 142344 24268 142396 24274
rect 142344 24210 142396 24216
rect 142434 10976 142490 10985
rect 142434 10911 142490 10920
rect 142252 4140 142304 4146
rect 142252 4082 142304 4088
rect 142160 3392 142212 3398
rect 142160 3334 142212 3340
rect 142448 480 142476 10911
rect 142908 3738 142936 74258
rect 143000 73982 143028 79648
rect 143092 78169 143120 79784
rect 143322 79812 143350 80036
rect 143414 79937 143442 80036
rect 143400 79928 143456 79937
rect 143400 79863 143456 79872
rect 143506 79812 143534 80036
rect 143598 79937 143626 80036
rect 143690 79966 143718 80036
rect 143782 79971 143810 80036
rect 143678 79960 143730 79966
rect 143584 79928 143640 79937
rect 143678 79902 143730 79908
rect 143768 79962 143824 79971
rect 143874 79966 143902 80036
rect 143768 79897 143824 79906
rect 143862 79960 143914 79966
rect 143862 79902 143914 79908
rect 143584 79863 143640 79872
rect 143966 79830 143994 80036
rect 144058 79937 144086 80036
rect 144044 79928 144100 79937
rect 144150 79898 144178 80036
rect 144242 79966 144270 80036
rect 144334 79971 144362 80036
rect 144230 79960 144282 79966
rect 144230 79902 144282 79908
rect 144320 79962 144376 79971
rect 144426 79966 144454 80036
rect 144044 79863 144100 79872
rect 144138 79892 144190 79898
rect 144320 79897 144376 79906
rect 144414 79960 144466 79966
rect 144414 79902 144466 79908
rect 144138 79834 144190 79840
rect 143172 79766 143224 79772
rect 143276 79784 143350 79812
rect 143460 79784 143534 79812
rect 143954 79824 144006 79830
rect 143078 78160 143134 78169
rect 143078 78095 143134 78104
rect 143184 77110 143212 79766
rect 143276 78305 143304 79784
rect 143460 79778 143488 79784
rect 143414 79750 143488 79778
rect 144518 79801 144546 80036
rect 144610 79830 144638 80036
rect 144702 79966 144730 80036
rect 144690 79960 144742 79966
rect 144690 79902 144742 79908
rect 144794 79898 144822 80036
rect 144886 79971 144914 80036
rect 144872 79962 144928 79971
rect 144782 79892 144834 79898
rect 144872 79897 144928 79906
rect 144782 79834 144834 79840
rect 144598 79824 144650 79830
rect 143954 79766 144006 79772
rect 144274 79792 144330 79801
rect 143632 79756 143684 79762
rect 143414 79744 143442 79750
rect 143368 79716 143442 79744
rect 143368 78713 143396 79716
rect 143632 79698 143684 79704
rect 144184 79756 144236 79762
rect 144504 79792 144560 79801
rect 144274 79727 144330 79736
rect 144368 79756 144420 79762
rect 144184 79698 144236 79704
rect 143460 79665 143580 79676
rect 143460 79656 143594 79665
rect 143460 79648 143538 79656
rect 143354 78704 143410 78713
rect 143354 78639 143410 78648
rect 143262 78296 143318 78305
rect 143262 78231 143318 78240
rect 143172 77104 143224 77110
rect 143172 77046 143224 77052
rect 143460 77042 143488 79648
rect 143538 79591 143594 79600
rect 143540 79416 143592 79422
rect 143540 79358 143592 79364
rect 143552 79082 143580 79358
rect 143540 79076 143592 79082
rect 143540 79018 143592 79024
rect 143540 77852 143592 77858
rect 143540 77794 143592 77800
rect 143448 77036 143500 77042
rect 143448 76978 143500 76984
rect 142988 73976 143040 73982
rect 142988 73918 143040 73924
rect 143552 70394 143580 77794
rect 143644 75274 143672 79698
rect 143724 79688 143776 79694
rect 144000 79688 144052 79694
rect 143724 79630 143776 79636
rect 143814 79656 143870 79665
rect 143632 75268 143684 75274
rect 143632 75210 143684 75216
rect 143552 70366 143672 70394
rect 143540 4412 143592 4418
rect 143540 4354 143592 4360
rect 142896 3732 142948 3738
rect 142896 3674 142948 3680
rect 143552 480 143580 4354
rect 143644 3942 143672 70366
rect 143736 4078 143764 79630
rect 144000 79630 144052 79636
rect 143814 79591 143870 79600
rect 143828 4962 143856 79591
rect 143906 78704 143962 78713
rect 143906 78639 143962 78648
rect 143920 20262 143948 78639
rect 144012 25702 144040 79630
rect 144092 79484 144144 79490
rect 144092 79426 144144 79432
rect 144104 79014 144132 79426
rect 144092 79008 144144 79014
rect 144092 78950 144144 78956
rect 144196 76974 144224 79698
rect 144184 76968 144236 76974
rect 144184 76910 144236 76916
rect 144288 75914 144316 79727
rect 144598 79766 144650 79772
rect 144872 79792 144928 79801
rect 144504 79727 144560 79736
rect 144736 79756 144788 79762
rect 144368 79698 144420 79704
rect 144736 79698 144788 79704
rect 144840 79736 144872 79744
rect 144840 79727 144928 79736
rect 144840 79716 144914 79727
rect 144380 77858 144408 79698
rect 144460 79688 144512 79694
rect 144460 79630 144512 79636
rect 144644 79688 144696 79694
rect 144644 79630 144696 79636
rect 144472 78606 144500 79630
rect 144552 79620 144604 79626
rect 144552 79562 144604 79568
rect 144460 78600 144512 78606
rect 144460 78542 144512 78548
rect 144368 77852 144420 77858
rect 144368 77794 144420 77800
rect 144460 76560 144512 76566
rect 144460 76502 144512 76508
rect 144104 75886 144316 75914
rect 144104 31278 144132 75886
rect 144184 75268 144236 75274
rect 144184 75210 144236 75216
rect 144196 46374 144224 75210
rect 144276 60716 144328 60722
rect 144276 60658 144328 60664
rect 144184 46368 144236 46374
rect 144184 46310 144236 46316
rect 144092 31272 144144 31278
rect 144092 31214 144144 31220
rect 144000 25696 144052 25702
rect 144000 25638 144052 25644
rect 143908 20256 143960 20262
rect 143908 20198 143960 20204
rect 143816 4956 143868 4962
rect 143816 4898 143868 4904
rect 143724 4072 143776 4078
rect 143724 4014 143776 4020
rect 143632 3936 143684 3942
rect 143632 3878 143684 3884
rect 144288 3602 144316 60658
rect 144276 3596 144328 3602
rect 144276 3538 144328 3544
rect 144472 3194 144500 76502
rect 144564 4010 144592 79562
rect 144656 74089 144684 79630
rect 144748 76945 144776 79698
rect 144734 76936 144790 76945
rect 144734 76871 144790 76880
rect 144642 74080 144698 74089
rect 144642 74015 144698 74024
rect 144840 73681 144868 79716
rect 144978 79676 145006 80036
rect 145070 79971 145098 80036
rect 145056 79962 145112 79971
rect 145162 79966 145190 80036
rect 145254 79966 145282 80036
rect 145346 79966 145374 80036
rect 145438 79966 145466 80036
rect 145056 79897 145112 79906
rect 145150 79960 145202 79966
rect 145150 79902 145202 79908
rect 145242 79960 145294 79966
rect 145242 79902 145294 79908
rect 145334 79960 145386 79966
rect 145334 79902 145386 79908
rect 145426 79960 145478 79966
rect 145426 79902 145478 79908
rect 145288 79824 145340 79830
rect 145288 79766 145340 79772
rect 145196 79756 145248 79762
rect 145196 79698 145248 79704
rect 144932 79648 145006 79676
rect 145104 79688 145156 79694
rect 144932 77654 144960 79648
rect 145104 79630 145156 79636
rect 145116 78792 145144 79630
rect 145024 78764 145144 78792
rect 144920 77648 144972 77654
rect 144920 77590 144972 77596
rect 145024 77500 145052 78764
rect 145102 78704 145158 78713
rect 145102 78639 145158 78648
rect 144932 77472 145052 77500
rect 144826 73672 144882 73681
rect 144826 73607 144882 73616
rect 144932 14822 144960 77472
rect 145012 77376 145064 77382
rect 145012 77318 145064 77324
rect 145024 20058 145052 77318
rect 145116 76702 145144 78639
rect 145208 78402 145236 79698
rect 145300 78606 145328 79766
rect 145530 79676 145558 80036
rect 145622 79966 145650 80036
rect 145610 79960 145662 79966
rect 145610 79902 145662 79908
rect 145714 79744 145742 80036
rect 145806 79937 145834 80036
rect 145792 79928 145848 79937
rect 145792 79863 145848 79872
rect 145668 79716 145742 79744
rect 145898 79744 145926 80036
rect 145990 79898 146018 80036
rect 145978 79892 146030 79898
rect 145978 79834 146030 79840
rect 146082 79778 146110 80036
rect 146174 79966 146202 80036
rect 146162 79960 146214 79966
rect 146162 79902 146214 79908
rect 146266 79812 146294 80036
rect 146036 79750 146110 79778
rect 146220 79784 146294 79812
rect 145898 79716 145972 79744
rect 145530 79648 145604 79676
rect 145380 79620 145432 79626
rect 145380 79562 145432 79568
rect 145288 78600 145340 78606
rect 145288 78542 145340 78548
rect 145196 78396 145248 78402
rect 145196 78338 145248 78344
rect 145392 77976 145420 79562
rect 145300 77948 145420 77976
rect 145104 76696 145156 76702
rect 145104 76638 145156 76644
rect 145194 76392 145250 76401
rect 145194 76327 145250 76336
rect 145104 76084 145156 76090
rect 145104 76026 145156 76032
rect 145116 20194 145144 76026
rect 145208 25634 145236 76327
rect 145300 26994 145328 77948
rect 145380 76696 145432 76702
rect 145380 76638 145432 76644
rect 145392 76548 145420 76638
rect 145392 76520 145512 76548
rect 145380 76356 145432 76362
rect 145380 76298 145432 76304
rect 145392 49298 145420 76298
rect 145484 61606 145512 76520
rect 145576 64394 145604 79648
rect 145668 76362 145696 79716
rect 145944 79642 145972 79716
rect 146036 79665 146064 79750
rect 146116 79688 146168 79694
rect 145748 79620 145800 79626
rect 145748 79562 145800 79568
rect 145852 79614 145972 79642
rect 146022 79656 146078 79665
rect 145760 77382 145788 79562
rect 145852 78334 145880 79614
rect 146116 79630 146168 79636
rect 146022 79591 146078 79600
rect 145932 79552 145984 79558
rect 145932 79494 145984 79500
rect 145840 78328 145892 78334
rect 145840 78270 145892 78276
rect 145748 77376 145800 77382
rect 145748 77318 145800 77324
rect 145656 76356 145708 76362
rect 145656 76298 145708 76304
rect 145944 76090 145972 79494
rect 146022 78704 146078 78713
rect 146022 78639 146078 78648
rect 146036 76634 146064 78639
rect 146128 78169 146156 79630
rect 146114 78160 146170 78169
rect 146114 78095 146170 78104
rect 146024 76628 146076 76634
rect 146024 76570 146076 76576
rect 146220 76537 146248 79784
rect 146358 79744 146386 80036
rect 146450 79937 146478 80036
rect 146542 79966 146570 80036
rect 146530 79960 146582 79966
rect 146436 79928 146492 79937
rect 146530 79902 146582 79908
rect 146436 79863 146492 79872
rect 146312 79716 146386 79744
rect 146484 79756 146536 79762
rect 146312 76838 146340 79716
rect 146634 79744 146662 80036
rect 146726 79971 146754 80036
rect 146712 79962 146768 79971
rect 146818 79966 146846 80036
rect 146910 79966 146938 80036
rect 146712 79897 146768 79906
rect 146806 79960 146858 79966
rect 146806 79902 146858 79908
rect 146898 79960 146950 79966
rect 146898 79902 146950 79908
rect 147002 79812 147030 80036
rect 147094 79966 147122 80036
rect 147082 79960 147134 79966
rect 147082 79902 147134 79908
rect 147186 79812 147214 80036
rect 147278 79937 147306 80036
rect 147264 79928 147320 79937
rect 147264 79863 147320 79872
rect 146758 79792 146814 79801
rect 146634 79716 146708 79744
rect 147002 79784 147076 79812
rect 147186 79784 147260 79812
rect 146758 79727 146814 79736
rect 146484 79698 146536 79704
rect 146496 78792 146524 79698
rect 146680 79665 146708 79716
rect 146666 79656 146722 79665
rect 146576 79620 146628 79626
rect 146666 79591 146722 79600
rect 146576 79562 146628 79568
rect 146404 78764 146524 78792
rect 146300 76832 146352 76838
rect 146300 76774 146352 76780
rect 146298 76664 146354 76673
rect 146298 76599 146354 76608
rect 146206 76528 146262 76537
rect 146206 76463 146262 76472
rect 145932 76084 145984 76090
rect 145932 76026 145984 76032
rect 145564 64388 145616 64394
rect 145564 64330 145616 64336
rect 145472 61600 145524 61606
rect 145472 61542 145524 61548
rect 145380 49292 145432 49298
rect 145380 49234 145432 49240
rect 145288 26988 145340 26994
rect 145288 26930 145340 26936
rect 145196 25628 145248 25634
rect 145196 25570 145248 25576
rect 145104 20188 145156 20194
rect 145104 20130 145156 20136
rect 145012 20052 145064 20058
rect 145012 19994 145064 20000
rect 144920 14816 144972 14822
rect 144920 14758 144972 14764
rect 144552 4004 144604 4010
rect 144552 3946 144604 3952
rect 146312 3874 146340 76599
rect 146404 6050 146432 78764
rect 146484 78668 146536 78674
rect 146484 78610 146536 78616
rect 146496 6866 146524 78610
rect 146484 6860 146536 6866
rect 146484 6802 146536 6808
rect 146588 6118 146616 79562
rect 146668 79280 146720 79286
rect 146668 79222 146720 79228
rect 146680 79150 146708 79222
rect 146668 79144 146720 79150
rect 146668 79086 146720 79092
rect 146668 78736 146720 78742
rect 146668 78678 146720 78684
rect 146680 9586 146708 78678
rect 146772 77294 146800 79727
rect 146944 79688 146996 79694
rect 146944 79630 146996 79636
rect 146852 79620 146904 79626
rect 146852 79562 146904 79568
rect 146864 77897 146892 79562
rect 146850 77888 146906 77897
rect 146850 77823 146906 77832
rect 146772 77266 146892 77294
rect 146760 76628 146812 76634
rect 146760 76570 146812 76576
rect 146668 9580 146720 9586
rect 146668 9522 146720 9528
rect 146772 8906 146800 76570
rect 146864 9654 146892 77266
rect 146956 12238 146984 79630
rect 147048 78742 147076 79784
rect 147128 79688 147180 79694
rect 147128 79630 147180 79636
rect 147036 78736 147088 78742
rect 147036 78678 147088 78684
rect 147140 77294 147168 79630
rect 147232 78674 147260 79784
rect 147370 79744 147398 80036
rect 147462 79971 147490 80036
rect 147448 79962 147504 79971
rect 147448 79897 147504 79906
rect 147554 79898 147582 80036
rect 147542 79892 147594 79898
rect 147542 79834 147594 79840
rect 147646 79830 147674 80036
rect 147634 79824 147686 79830
rect 147634 79766 147686 79772
rect 147738 79744 147766 80036
rect 147830 79966 147858 80036
rect 147818 79960 147870 79966
rect 147818 79902 147870 79908
rect 147922 79778 147950 80036
rect 148014 79966 148042 80036
rect 148002 79960 148054 79966
rect 148002 79902 148054 79908
rect 147876 79750 147950 79778
rect 147370 79716 147444 79744
rect 147738 79716 147812 79744
rect 147220 78668 147272 78674
rect 147220 78610 147272 78616
rect 147312 78396 147364 78402
rect 147312 78338 147364 78344
rect 147048 77266 147168 77294
rect 147048 12306 147076 77266
rect 147324 73914 147352 78338
rect 147416 76673 147444 79716
rect 147588 79688 147640 79694
rect 147494 79656 147550 79665
rect 147588 79630 147640 79636
rect 147494 79591 147550 79600
rect 147402 76664 147458 76673
rect 147402 76599 147458 76608
rect 147508 76537 147536 79591
rect 147600 76809 147628 79630
rect 147680 79552 147732 79558
rect 147680 79494 147732 79500
rect 147692 79286 147720 79494
rect 147680 79280 147732 79286
rect 147680 79222 147732 79228
rect 147680 78668 147732 78674
rect 147680 78610 147732 78616
rect 147586 76800 147642 76809
rect 147586 76735 147642 76744
rect 147494 76528 147550 76537
rect 147494 76463 147550 76472
rect 147312 73908 147364 73914
rect 147312 73850 147364 73856
rect 147036 12300 147088 12306
rect 147036 12242 147088 12248
rect 146944 12232 146996 12238
rect 146944 12174 146996 12180
rect 147692 12170 147720 78610
rect 147784 76770 147812 79716
rect 147876 78674 147904 79750
rect 148106 79744 148134 80036
rect 148198 79812 148226 80036
rect 148290 79937 148318 80036
rect 148276 79928 148332 79937
rect 148382 79898 148410 80036
rect 148474 79898 148502 80036
rect 148566 79966 148594 80036
rect 148658 79966 148686 80036
rect 148554 79960 148606 79966
rect 148554 79902 148606 79908
rect 148646 79960 148698 79966
rect 148646 79902 148698 79908
rect 148276 79863 148332 79872
rect 148370 79892 148422 79898
rect 148370 79834 148422 79840
rect 148462 79892 148514 79898
rect 148462 79834 148514 79840
rect 148750 79830 148778 80036
rect 148738 79824 148790 79830
rect 148198 79801 148272 79812
rect 148198 79792 148286 79801
rect 148198 79784 148230 79792
rect 148106 79716 148180 79744
rect 148738 79766 148790 79772
rect 148230 79727 148286 79736
rect 147956 79688 148008 79694
rect 147956 79630 148008 79636
rect 147864 78668 147916 78674
rect 147864 78610 147916 78616
rect 147968 77518 147996 79630
rect 148048 79620 148100 79626
rect 148048 79562 148100 79568
rect 147956 77512 148008 77518
rect 147956 77454 148008 77460
rect 147772 76764 147824 76770
rect 147772 76706 147824 76712
rect 147956 76628 148008 76634
rect 147956 76570 148008 76576
rect 147862 76528 147918 76537
rect 147772 76492 147824 76498
rect 147862 76463 147918 76472
rect 147772 76434 147824 76440
rect 147784 24206 147812 76434
rect 147876 32502 147904 76463
rect 147864 32496 147916 32502
rect 147864 32438 147916 32444
rect 147968 32434 147996 76570
rect 148060 43586 148088 79562
rect 148152 45014 148180 79716
rect 148232 79688 148284 79694
rect 148416 79688 148468 79694
rect 148232 79630 148284 79636
rect 148322 79656 148378 79665
rect 148244 60178 148272 79630
rect 148416 79630 148468 79636
rect 148692 79688 148744 79694
rect 148842 79676 148870 80036
rect 148934 79801 148962 80036
rect 149026 79966 149054 80036
rect 149014 79960 149066 79966
rect 149014 79902 149066 79908
rect 148920 79792 148976 79801
rect 149118 79778 149146 80036
rect 148920 79727 148976 79736
rect 149072 79750 149146 79778
rect 149210 79778 149238 80036
rect 149302 79898 149330 80036
rect 149394 79966 149422 80036
rect 149382 79960 149434 79966
rect 149382 79902 149434 79908
rect 149290 79892 149342 79898
rect 149290 79834 149342 79840
rect 149486 79812 149514 80036
rect 149578 79937 149606 80036
rect 149670 79966 149698 80036
rect 149658 79960 149710 79966
rect 149564 79928 149620 79937
rect 149658 79902 149710 79908
rect 149564 79863 149620 79872
rect 149486 79784 149560 79812
rect 149210 79750 149376 79778
rect 148692 79630 148744 79636
rect 148796 79648 148870 79676
rect 148968 79688 149020 79694
rect 148322 79591 148378 79600
rect 148336 65754 148364 79591
rect 148428 76634 148456 79630
rect 148600 79552 148652 79558
rect 148600 79494 148652 79500
rect 148416 76628 148468 76634
rect 148416 76570 148468 76576
rect 148612 76498 148640 79494
rect 148600 76492 148652 76498
rect 148600 76434 148652 76440
rect 148704 73953 148732 79630
rect 148796 78305 148824 79648
rect 148968 79630 149020 79636
rect 148782 78296 148838 78305
rect 148782 78231 148838 78240
rect 148784 78124 148836 78130
rect 148784 78066 148836 78072
rect 148690 73944 148746 73953
rect 148690 73879 148746 73888
rect 148796 70394 148824 78066
rect 148980 77897 149008 79630
rect 149072 78198 149100 79750
rect 149152 79688 149204 79694
rect 149152 79630 149204 79636
rect 149060 78192 149112 78198
rect 149060 78134 149112 78140
rect 149164 77976 149192 79630
rect 149244 79620 149296 79626
rect 149244 79562 149296 79568
rect 149256 78033 149284 79562
rect 149072 77948 149192 77976
rect 149242 78024 149298 78033
rect 149242 77959 149298 77968
rect 148966 77888 149022 77897
rect 148966 77823 149022 77832
rect 148704 70366 148824 70394
rect 148324 65748 148376 65754
rect 148324 65690 148376 65696
rect 148704 62966 148732 70366
rect 148692 62960 148744 62966
rect 148692 62902 148744 62908
rect 148232 60172 148284 60178
rect 148232 60114 148284 60120
rect 148140 45008 148192 45014
rect 148140 44950 148192 44956
rect 148048 43580 148100 43586
rect 148048 43522 148100 43528
rect 147956 32428 148008 32434
rect 147956 32370 148008 32376
rect 147772 24200 147824 24206
rect 147772 24142 147824 24148
rect 147772 21480 147824 21486
rect 147772 21422 147824 21428
rect 147784 16574 147812 21422
rect 147784 16546 147904 16574
rect 147680 12164 147732 12170
rect 147680 12106 147732 12112
rect 146852 9648 146904 9654
rect 146852 9590 146904 9596
rect 146760 8900 146812 8906
rect 146760 8842 146812 8848
rect 146576 6112 146628 6118
rect 146576 6054 146628 6060
rect 146392 6044 146444 6050
rect 146392 5986 146444 5992
rect 144736 3868 144788 3874
rect 144736 3810 144788 3816
rect 146300 3868 146352 3874
rect 146300 3810 146352 3816
rect 144460 3188 144512 3194
rect 144460 3130 144512 3136
rect 144748 480 144776 3810
rect 145932 3800 145984 3806
rect 145932 3742 145984 3748
rect 145944 480 145972 3742
rect 147128 3664 147180 3670
rect 147128 3606 147180 3612
rect 147140 480 147168 3606
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149072 3806 149100 77948
rect 149152 77852 149204 77858
rect 149152 77794 149204 77800
rect 149164 6730 149192 77794
rect 149348 76480 149376 79750
rect 149428 79688 149480 79694
rect 149428 79630 149480 79636
rect 149440 77722 149468 79630
rect 149428 77716 149480 77722
rect 149428 77658 149480 77664
rect 149256 76452 149376 76480
rect 149256 75274 149284 76452
rect 149532 75914 149560 79784
rect 149762 79778 149790 80036
rect 149854 79966 149882 80036
rect 149842 79960 149894 79966
rect 149842 79902 149894 79908
rect 149946 79898 149974 80036
rect 149934 79892 149986 79898
rect 149934 79834 149986 79840
rect 150038 79830 150066 80036
rect 150130 79937 150158 80036
rect 150116 79928 150172 79937
rect 150116 79863 150172 79872
rect 149612 79756 149664 79762
rect 149612 79698 149664 79704
rect 149716 79750 149790 79778
rect 150026 79824 150078 79830
rect 150222 79812 150250 80036
rect 150314 79898 150342 80036
rect 150302 79892 150354 79898
rect 150302 79834 150354 79840
rect 150026 79766 150078 79772
rect 150176 79784 150250 79812
rect 149348 75886 149560 75914
rect 149244 75268 149296 75274
rect 149244 75210 149296 75216
rect 149244 75132 149296 75138
rect 149244 75074 149296 75080
rect 149256 6798 149284 75074
rect 149348 9450 149376 75886
rect 149428 75268 149480 75274
rect 149428 75210 149480 75216
rect 149520 75268 149572 75274
rect 149520 75210 149572 75216
rect 149440 9518 149468 75210
rect 149532 12102 149560 75210
rect 149624 75138 149652 79698
rect 149716 79472 149744 79750
rect 149888 79688 149940 79694
rect 149888 79630 149940 79636
rect 149716 79444 149836 79472
rect 149702 78160 149758 78169
rect 149702 78095 149758 78104
rect 149612 75132 149664 75138
rect 149612 75074 149664 75080
rect 149612 74996 149664 75002
rect 149612 74938 149664 74944
rect 149520 12096 149572 12102
rect 149520 12038 149572 12044
rect 149624 12034 149652 74938
rect 149716 14686 149744 78095
rect 149808 75274 149836 79444
rect 149900 77858 149928 79630
rect 149980 79620 150032 79626
rect 149980 79562 150032 79568
rect 149888 77852 149940 77858
rect 149888 77794 149940 77800
rect 149888 77716 149940 77722
rect 149888 77658 149940 77664
rect 149796 75268 149848 75274
rect 149796 75210 149848 75216
rect 149900 64874 149928 77658
rect 149992 75002 150020 79562
rect 150176 78169 150204 79784
rect 150256 79688 150308 79694
rect 150406 79676 150434 80036
rect 150498 79966 150526 80036
rect 150486 79960 150538 79966
rect 150486 79902 150538 79908
rect 150590 79778 150618 80036
rect 150682 79971 150710 80036
rect 150668 79962 150724 79971
rect 150774 79966 150802 80036
rect 150866 79966 150894 80036
rect 150958 79966 150986 80036
rect 151050 79966 151078 80036
rect 150668 79897 150724 79906
rect 150762 79960 150814 79966
rect 150762 79902 150814 79908
rect 150854 79960 150906 79966
rect 150854 79902 150906 79908
rect 150946 79960 150998 79966
rect 150946 79902 150998 79908
rect 151038 79960 151090 79966
rect 151038 79902 151090 79908
rect 150898 79792 150954 79801
rect 150590 79750 150664 79778
rect 150256 79630 150308 79636
rect 150360 79648 150434 79676
rect 150162 78160 150218 78169
rect 150162 78095 150218 78104
rect 150268 77897 150296 79630
rect 150254 77888 150310 77897
rect 150254 77823 150310 77832
rect 150360 76673 150388 79648
rect 150532 79620 150584 79626
rect 150532 79562 150584 79568
rect 150440 79008 150492 79014
rect 150440 78950 150492 78956
rect 150346 76664 150402 76673
rect 150346 76599 150402 76608
rect 149980 74996 150032 75002
rect 149980 74938 150032 74944
rect 149808 64846 149928 64874
rect 149808 14754 149836 64846
rect 149796 14748 149848 14754
rect 149796 14690 149848 14696
rect 149704 14680 149756 14686
rect 149704 14622 149756 14628
rect 149612 12028 149664 12034
rect 149612 11970 149664 11976
rect 149428 9512 149480 9518
rect 149428 9454 149480 9460
rect 149336 9444 149388 9450
rect 149336 9386 149388 9392
rect 150452 7682 150480 78950
rect 150544 77450 150572 79562
rect 150532 77444 150584 77450
rect 150532 77386 150584 77392
rect 150532 75200 150584 75206
rect 150532 75142 150584 75148
rect 150544 22982 150572 75142
rect 150636 28422 150664 79750
rect 150898 79727 150954 79736
rect 151142 79744 151170 80036
rect 151234 79937 151262 80036
rect 151326 79966 151354 80036
rect 151314 79960 151366 79966
rect 151220 79928 151276 79937
rect 151314 79902 151366 79908
rect 151418 79898 151446 80036
rect 151220 79863 151276 79872
rect 151406 79892 151458 79898
rect 151406 79834 151458 79840
rect 151510 79778 151538 80036
rect 151268 79756 151320 79762
rect 150808 79620 150860 79626
rect 150808 79562 150860 79568
rect 150820 78860 150848 79562
rect 150912 79014 150940 79727
rect 151142 79716 151216 79744
rect 151084 79620 151136 79626
rect 151084 79562 151136 79568
rect 150992 79552 151044 79558
rect 150992 79494 151044 79500
rect 150900 79008 150952 79014
rect 150900 78950 150952 78956
rect 151004 78946 151032 79494
rect 150992 78940 151044 78946
rect 150992 78882 151044 78888
rect 150820 78832 150940 78860
rect 150912 78402 150940 78832
rect 151096 78792 151124 79562
rect 151004 78764 151124 78792
rect 150716 78396 150768 78402
rect 150716 78338 150768 78344
rect 150900 78396 150952 78402
rect 150900 78338 150952 78344
rect 150728 29850 150756 78338
rect 150808 78328 150860 78334
rect 151004 78282 151032 78764
rect 151084 78668 151136 78674
rect 151084 78610 151136 78616
rect 150808 78270 150860 78276
rect 150820 76906 150848 78270
rect 150912 78254 151032 78282
rect 150808 76900 150860 76906
rect 150808 76842 150860 76848
rect 150808 75268 150860 75274
rect 150808 75210 150860 75216
rect 150820 55962 150848 75210
rect 150912 58954 150940 78254
rect 150990 78160 151046 78169
rect 150990 78095 151046 78104
rect 151004 75546 151032 78095
rect 150992 75540 151044 75546
rect 150992 75482 151044 75488
rect 151096 72826 151124 78610
rect 151188 75206 151216 79716
rect 151268 79698 151320 79704
rect 151360 79756 151412 79762
rect 151360 79698 151412 79704
rect 151464 79750 151538 79778
rect 151280 75274 151308 79698
rect 151268 75268 151320 75274
rect 151268 75210 151320 75216
rect 151176 75200 151228 75206
rect 151176 75142 151228 75148
rect 151084 72820 151136 72826
rect 151084 72762 151136 72768
rect 151372 70394 151400 79698
rect 151464 72758 151492 79750
rect 151602 79676 151630 80036
rect 151694 79971 151722 80036
rect 151680 79962 151736 79971
rect 151680 79897 151736 79906
rect 151786 79812 151814 80036
rect 151740 79784 151814 79812
rect 151602 79648 151676 79676
rect 151648 78713 151676 79648
rect 151634 78704 151690 78713
rect 151634 78639 151690 78648
rect 151740 78441 151768 79784
rect 151878 79744 151906 80036
rect 151970 79937 151998 80036
rect 152062 79966 152090 80036
rect 152154 79966 152182 80036
rect 152050 79960 152102 79966
rect 151956 79928 152012 79937
rect 152050 79902 152102 79908
rect 152142 79960 152194 79966
rect 152142 79902 152194 79908
rect 151956 79863 152012 79872
rect 152050 79824 152102 79830
rect 151832 79716 151906 79744
rect 152016 79772 152050 79778
rect 152246 79812 152274 80036
rect 152338 79971 152366 80036
rect 152324 79962 152380 79971
rect 152430 79966 152458 80036
rect 152324 79897 152380 79906
rect 152418 79960 152470 79966
rect 152418 79902 152470 79908
rect 152522 79898 152550 80036
rect 152614 79971 152642 80036
rect 152600 79962 152656 79971
rect 152510 79892 152562 79898
rect 152600 79897 152656 79906
rect 152706 79898 152734 80036
rect 152798 79966 152826 80036
rect 152890 79966 152918 80036
rect 152982 79966 153010 80036
rect 152786 79960 152838 79966
rect 152786 79902 152838 79908
rect 152878 79960 152930 79966
rect 152878 79902 152930 79908
rect 152970 79960 153022 79966
rect 152970 79902 153022 79908
rect 153074 79898 153102 80036
rect 153166 79966 153194 80036
rect 153258 79966 153286 80036
rect 153350 79966 153378 80036
rect 153442 79971 153470 80036
rect 153154 79960 153206 79966
rect 153154 79902 153206 79908
rect 153246 79960 153298 79966
rect 153246 79902 153298 79908
rect 153338 79960 153390 79966
rect 153338 79902 153390 79908
rect 153428 79962 153484 79971
rect 152510 79834 152562 79840
rect 152694 79892 152746 79898
rect 152694 79834 152746 79840
rect 153062 79892 153114 79898
rect 153428 79897 153484 79906
rect 153062 79834 153114 79840
rect 152016 79766 152102 79772
rect 152200 79784 152274 79812
rect 152878 79824 152930 79830
rect 152738 79792 152794 79801
rect 152016 79750 152090 79766
rect 151726 78432 151782 78441
rect 151726 78367 151782 78376
rect 151544 78192 151596 78198
rect 151544 78134 151596 78140
rect 151556 76634 151584 78134
rect 151544 76628 151596 76634
rect 151544 76570 151596 76576
rect 151452 72752 151504 72758
rect 151452 72694 151504 72700
rect 151004 70366 151400 70394
rect 151004 68610 151032 70366
rect 150992 68604 151044 68610
rect 150992 68546 151044 68552
rect 150900 58948 150952 58954
rect 150900 58890 150952 58896
rect 150808 55956 150860 55962
rect 150808 55898 150860 55904
rect 150716 29844 150768 29850
rect 150716 29786 150768 29792
rect 150624 28416 150676 28422
rect 150624 28358 150676 28364
rect 150532 22976 150584 22982
rect 150532 22918 150584 22924
rect 150440 7676 150492 7682
rect 150440 7618 150492 7624
rect 149244 6792 149296 6798
rect 149244 6734 149296 6740
rect 149152 6724 149204 6730
rect 149152 6666 149204 6672
rect 151832 6594 151860 79716
rect 151912 79620 151964 79626
rect 151912 79562 151964 79568
rect 151924 78742 151952 79562
rect 151912 78736 151964 78742
rect 151912 78678 151964 78684
rect 151912 77308 151964 77314
rect 151912 77250 151964 77256
rect 151924 16182 151952 77250
rect 152016 72690 152044 79750
rect 152094 79656 152150 79665
rect 152094 79591 152150 79600
rect 152004 72684 152056 72690
rect 152004 72626 152056 72632
rect 152108 70394 152136 79591
rect 152200 77314 152228 79784
rect 152556 79756 152608 79762
rect 152794 79772 152878 79778
rect 152794 79766 152930 79772
rect 152794 79750 152918 79766
rect 153384 79756 153436 79762
rect 152738 79727 152794 79736
rect 152556 79698 152608 79704
rect 153534 79744 153562 80036
rect 153626 79966 153654 80036
rect 153614 79960 153666 79966
rect 153614 79902 153666 79908
rect 153718 79830 153746 80036
rect 153706 79824 153758 79830
rect 153810 79801 153838 80036
rect 153902 79898 153930 80036
rect 153994 79937 154022 80036
rect 154086 79966 154114 80036
rect 154178 79966 154206 80036
rect 154270 79966 154298 80036
rect 154362 79966 154390 80036
rect 154074 79960 154126 79966
rect 153980 79928 154036 79937
rect 153890 79892 153942 79898
rect 154074 79902 154126 79908
rect 154166 79960 154218 79966
rect 154166 79902 154218 79908
rect 154258 79960 154310 79966
rect 154258 79902 154310 79908
rect 154350 79960 154402 79966
rect 154454 79937 154482 80036
rect 154546 79966 154574 80036
rect 154534 79960 154586 79966
rect 154350 79902 154402 79908
rect 154440 79928 154496 79937
rect 153980 79863 154036 79872
rect 154638 79937 154666 80036
rect 154534 79902 154586 79908
rect 154624 79928 154680 79937
rect 154440 79863 154496 79872
rect 154624 79863 154680 79872
rect 153890 79834 153942 79840
rect 154730 79830 154758 80036
rect 154822 79966 154850 80036
rect 154914 79966 154942 80036
rect 155006 79971 155034 80036
rect 154810 79960 154862 79966
rect 154810 79902 154862 79908
rect 154902 79960 154954 79966
rect 154902 79902 154954 79908
rect 154992 79962 155048 79971
rect 154992 79897 155048 79906
rect 155098 79898 155126 80036
rect 155190 79971 155218 80036
rect 155176 79962 155232 79971
rect 155282 79966 155310 80036
rect 155086 79892 155138 79898
rect 155176 79897 155232 79906
rect 155270 79960 155322 79966
rect 155374 79937 155402 80036
rect 155466 79966 155494 80036
rect 155558 79966 155586 80036
rect 155650 79971 155678 80036
rect 155454 79960 155506 79966
rect 155270 79902 155322 79908
rect 155360 79928 155416 79937
rect 155454 79902 155506 79908
rect 155546 79960 155598 79966
rect 155546 79902 155598 79908
rect 155636 79962 155692 79971
rect 155636 79897 155692 79906
rect 155742 79898 155770 80036
rect 155834 79971 155862 80036
rect 155820 79962 155876 79971
rect 155926 79966 155954 80036
rect 156018 79966 156046 80036
rect 156110 79971 156138 80036
rect 155360 79863 155416 79872
rect 155730 79892 155782 79898
rect 155820 79897 155876 79906
rect 155914 79960 155966 79966
rect 155914 79902 155966 79908
rect 156006 79960 156058 79966
rect 156006 79902 156058 79908
rect 156096 79962 156152 79971
rect 156096 79897 156152 79906
rect 155086 79834 155138 79840
rect 155730 79834 155782 79840
rect 154212 79824 154264 79830
rect 153706 79766 153758 79772
rect 153796 79792 153852 79801
rect 153384 79698 153436 79704
rect 153488 79716 153562 79744
rect 154212 79766 154264 79772
rect 154580 79824 154632 79830
rect 154580 79766 154632 79772
rect 154718 79824 154770 79830
rect 155224 79824 155276 79830
rect 154718 79766 154770 79772
rect 155130 79792 155186 79801
rect 153796 79727 153852 79736
rect 154028 79756 154080 79762
rect 152280 79688 152332 79694
rect 152280 79630 152332 79636
rect 152188 77308 152240 77314
rect 152188 77250 152240 77256
rect 152186 77208 152242 77217
rect 152186 77143 152242 77152
rect 152016 70366 152136 70394
rect 152016 20126 152044 70366
rect 152200 29782 152228 77143
rect 152292 40798 152320 79630
rect 152464 79552 152516 79558
rect 152464 79494 152516 79500
rect 152476 78198 152504 79494
rect 152464 78192 152516 78198
rect 152464 78134 152516 78140
rect 152464 78056 152516 78062
rect 152464 77998 152516 78004
rect 152476 76498 152504 77998
rect 152568 76702 152596 79698
rect 152832 79688 152884 79694
rect 152832 79630 152884 79636
rect 153016 79688 153068 79694
rect 153016 79630 153068 79636
rect 152648 79620 152700 79626
rect 152648 79562 152700 79568
rect 152556 76696 152608 76702
rect 152556 76638 152608 76644
rect 152464 76492 152516 76498
rect 152464 76434 152516 76440
rect 152660 70394 152688 79562
rect 152740 79552 152792 79558
rect 152740 79494 152792 79500
rect 152752 78441 152780 79494
rect 152844 78713 152872 79630
rect 152924 79552 152976 79558
rect 152924 79494 152976 79500
rect 152830 78704 152886 78713
rect 152830 78639 152886 78648
rect 152738 78432 152794 78441
rect 152738 78367 152794 78376
rect 152738 77480 152794 77489
rect 152738 77415 152794 77424
rect 152752 72622 152780 77415
rect 152936 77217 152964 79494
rect 152922 77208 152978 77217
rect 152922 77143 152978 77152
rect 153028 75138 153056 79630
rect 153108 78736 153160 78742
rect 153108 78678 153160 78684
rect 153120 77194 153148 78678
rect 153292 77852 153344 77858
rect 153292 77794 153344 77800
rect 153120 77166 153240 77194
rect 153108 76696 153160 76702
rect 153108 76638 153160 76644
rect 153016 75132 153068 75138
rect 153016 75074 153068 75080
rect 152740 72616 152792 72622
rect 152740 72558 152792 72564
rect 152384 70366 152688 70394
rect 152384 54670 152412 70366
rect 152372 54664 152424 54670
rect 152372 54606 152424 54612
rect 152280 40792 152332 40798
rect 152280 40734 152332 40740
rect 152188 29776 152240 29782
rect 152188 29718 152240 29724
rect 153120 29714 153148 76638
rect 153212 76430 153240 77166
rect 153200 76424 153252 76430
rect 153200 76366 153252 76372
rect 153200 76288 153252 76294
rect 153200 76230 153252 76236
rect 153108 29708 153160 29714
rect 153108 29650 153160 29656
rect 152004 20120 152056 20126
rect 152004 20062 152056 20068
rect 151912 16176 151964 16182
rect 151912 16118 151964 16124
rect 151820 6588 151872 6594
rect 151820 6530 151872 6536
rect 153212 6526 153240 76230
rect 153304 28354 153332 77794
rect 153396 39506 153424 79698
rect 153488 78062 153516 79716
rect 154028 79698 154080 79704
rect 153660 79688 153712 79694
rect 153566 79656 153622 79665
rect 153660 79630 153712 79636
rect 153936 79688 153988 79694
rect 153936 79630 153988 79636
rect 153566 79591 153622 79600
rect 153476 78056 153528 78062
rect 153476 77998 153528 78004
rect 153476 77240 153528 77246
rect 153476 77182 153528 77188
rect 153488 51814 153516 77182
rect 153580 54602 153608 79591
rect 153672 78334 153700 79630
rect 153752 79620 153804 79626
rect 153752 79562 153804 79568
rect 153660 78328 153712 78334
rect 153660 78270 153712 78276
rect 153660 78056 153712 78062
rect 153660 77998 153712 78004
rect 153672 58886 153700 77998
rect 153764 77858 153792 79562
rect 153844 79552 153896 79558
rect 153844 79494 153896 79500
rect 153752 77852 153804 77858
rect 153752 77794 153804 77800
rect 153856 70394 153884 79494
rect 153948 76294 153976 79630
rect 154040 77246 154068 79698
rect 154224 77314 154252 79766
rect 154304 79756 154356 79762
rect 154304 79698 154356 79704
rect 154316 78033 154344 79698
rect 154488 79620 154540 79626
rect 154488 79562 154540 79568
rect 154500 78062 154528 79562
rect 154592 78169 154620 79766
rect 154856 79756 154908 79762
rect 154856 79698 154908 79704
rect 155040 79756 155092 79762
rect 155224 79766 155276 79772
rect 155316 79824 155368 79830
rect 155868 79824 155920 79830
rect 155316 79766 155368 79772
rect 155774 79792 155830 79801
rect 155130 79727 155132 79736
rect 155040 79698 155092 79704
rect 155184 79727 155186 79736
rect 155132 79698 155184 79704
rect 154762 79656 154818 79665
rect 154762 79591 154818 79600
rect 154578 78160 154634 78169
rect 154578 78095 154634 78104
rect 154488 78056 154540 78062
rect 154302 78024 154358 78033
rect 154488 77998 154540 78004
rect 154302 77959 154358 77968
rect 154580 77988 154632 77994
rect 154580 77930 154632 77936
rect 154212 77308 154264 77314
rect 154212 77250 154264 77256
rect 154028 77240 154080 77246
rect 154028 77182 154080 77188
rect 153936 76288 153988 76294
rect 153936 76230 153988 76236
rect 154028 75132 154080 75138
rect 154028 75074 154080 75080
rect 153764 70366 153884 70394
rect 153764 67046 153792 70366
rect 153752 67040 153804 67046
rect 153752 66982 153804 66988
rect 153660 58880 153712 58886
rect 153660 58822 153712 58828
rect 153568 54596 153620 54602
rect 153568 54538 153620 54544
rect 153476 51808 153528 51814
rect 153476 51750 153528 51756
rect 154040 50726 154068 75074
rect 154028 50720 154080 50726
rect 154028 50662 154080 50668
rect 153844 47592 153896 47598
rect 153844 47534 153896 47540
rect 153384 39500 153436 39506
rect 153384 39442 153436 39448
rect 153292 28348 153344 28354
rect 153292 28290 153344 28296
rect 153752 11756 153804 11762
rect 153752 11698 153804 11704
rect 153200 6520 153252 6526
rect 153200 6462 153252 6468
rect 151820 4888 151872 4894
rect 151820 4830 151872 4836
rect 149060 3800 149112 3806
rect 149060 3742 149112 3748
rect 150624 3324 150676 3330
rect 150624 3266 150676 3272
rect 149520 3256 149572 3262
rect 149520 3198 149572 3204
rect 149532 480 149560 3198
rect 150636 480 150664 3266
rect 151832 480 151860 4830
rect 153016 3188 153068 3194
rect 153016 3130 153068 3136
rect 153028 480 153056 3130
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 11698
rect 153856 3126 153884 47534
rect 154592 21554 154620 77930
rect 154672 74724 154724 74730
rect 154672 74666 154724 74672
rect 154684 25566 154712 74666
rect 154776 26926 154804 79591
rect 154868 78742 154896 79698
rect 154948 79620 155000 79626
rect 154948 79562 155000 79568
rect 154856 78736 154908 78742
rect 154856 78678 154908 78684
rect 154856 78192 154908 78198
rect 154856 78134 154908 78140
rect 154868 55894 154896 78134
rect 154960 60110 154988 79562
rect 155052 77994 155080 79698
rect 155132 78056 155184 78062
rect 155132 77998 155184 78004
rect 155040 77988 155092 77994
rect 155040 77930 155092 77936
rect 155040 77784 155092 77790
rect 155040 77726 155092 77732
rect 155052 61538 155080 77726
rect 155144 66978 155172 77998
rect 155236 71262 155264 79766
rect 155328 78198 155356 79766
rect 156202 79812 156230 80036
rect 155868 79766 155920 79772
rect 156064 79784 156230 79812
rect 156294 79801 156322 80036
rect 156386 79966 156414 80036
rect 156478 79966 156506 80036
rect 156570 79971 156598 80036
rect 156374 79960 156426 79966
rect 156374 79902 156426 79908
rect 156466 79960 156518 79966
rect 156466 79902 156518 79908
rect 156556 79962 156612 79971
rect 156662 79966 156690 80036
rect 156754 79966 156782 80036
rect 156846 79966 156874 80036
rect 156556 79897 156612 79906
rect 156650 79960 156702 79966
rect 156650 79902 156702 79908
rect 156742 79960 156794 79966
rect 156742 79902 156794 79908
rect 156834 79960 156886 79966
rect 156834 79902 156886 79908
rect 156938 79898 156966 80036
rect 157030 79898 157058 80036
rect 157122 79903 157150 80036
rect 157214 79966 157242 80036
rect 157202 79960 157254 79966
rect 156926 79892 156978 79898
rect 156926 79834 156978 79840
rect 157018 79892 157070 79898
rect 157018 79834 157070 79840
rect 157108 79894 157164 79903
rect 157202 79902 157254 79908
rect 157306 79898 157334 80036
rect 157398 79971 157426 80036
rect 157384 79962 157440 79971
rect 157490 79966 157518 80036
rect 157108 79829 157164 79838
rect 157294 79892 157346 79898
rect 157384 79897 157440 79906
rect 157478 79960 157530 79966
rect 157478 79902 157530 79908
rect 157294 79834 157346 79840
rect 157432 79824 157484 79830
rect 156280 79792 156336 79801
rect 155774 79727 155830 79736
rect 155500 79688 155552 79694
rect 155500 79630 155552 79636
rect 155684 79688 155736 79694
rect 155684 79630 155736 79636
rect 155408 79620 155460 79626
rect 155408 79562 155460 79568
rect 155316 78192 155368 78198
rect 155316 78134 155368 78140
rect 155314 77888 155370 77897
rect 155314 77823 155370 77832
rect 155328 73846 155356 77823
rect 155420 77790 155448 79562
rect 155408 77784 155460 77790
rect 155408 77726 155460 77732
rect 155512 74730 155540 79630
rect 155592 79552 155644 79558
rect 155592 79494 155644 79500
rect 155500 74724 155552 74730
rect 155500 74666 155552 74672
rect 155316 73840 155368 73846
rect 155316 73782 155368 73788
rect 155604 71330 155632 79494
rect 155696 77897 155724 79630
rect 155682 77888 155738 77897
rect 155682 77823 155738 77832
rect 155788 76022 155816 79727
rect 155880 78878 155908 79766
rect 155960 79620 156012 79626
rect 155960 79562 156012 79568
rect 155868 78872 155920 78878
rect 155868 78814 155920 78820
rect 155972 78724 156000 79562
rect 155880 78696 156000 78724
rect 155880 77382 155908 78696
rect 156064 78656 156092 79784
rect 156786 79792 156842 79801
rect 156280 79727 156336 79736
rect 156604 79756 156656 79762
rect 156604 79698 156656 79704
rect 156708 79750 156786 79778
rect 156142 79656 156198 79665
rect 156142 79591 156198 79600
rect 156328 79620 156380 79626
rect 155972 78628 156092 78656
rect 155868 77376 155920 77382
rect 155868 77318 155920 77324
rect 155776 76016 155828 76022
rect 155776 75958 155828 75964
rect 155592 71324 155644 71330
rect 155592 71266 155644 71272
rect 155224 71256 155276 71262
rect 155224 71198 155276 71204
rect 155132 66972 155184 66978
rect 155132 66914 155184 66920
rect 155040 61532 155092 61538
rect 155040 61474 155092 61480
rect 154948 60104 155000 60110
rect 154948 60046 155000 60052
rect 154856 55888 154908 55894
rect 154856 55830 154908 55836
rect 155222 44840 155278 44849
rect 155222 44775 155278 44784
rect 154764 26920 154816 26926
rect 154764 26862 154816 26868
rect 154672 25560 154724 25566
rect 154672 25502 154724 25508
rect 154580 21548 154632 21554
rect 154580 21490 154632 21496
rect 155236 3670 155264 44775
rect 155972 6458 156000 78628
rect 156052 77988 156104 77994
rect 156052 77930 156104 77936
rect 156064 14550 156092 77930
rect 156156 77294 156184 79591
rect 156380 79580 156460 79608
rect 156328 79562 156380 79568
rect 156326 78704 156382 78713
rect 156326 78639 156382 78648
rect 156156 77266 156276 77294
rect 156144 76696 156196 76702
rect 156144 76638 156196 76644
rect 156156 19990 156184 76638
rect 156248 46306 156276 77266
rect 156340 76634 156368 78639
rect 156432 78266 156460 79580
rect 156512 79552 156564 79558
rect 156512 79494 156564 79500
rect 156420 78260 156472 78266
rect 156420 78202 156472 78208
rect 156524 78062 156552 79494
rect 156512 78056 156564 78062
rect 156512 77998 156564 78004
rect 156616 77994 156644 79698
rect 156604 77988 156656 77994
rect 156604 77930 156656 77936
rect 156708 77602 156736 79750
rect 157432 79766 157484 79772
rect 156786 79727 156842 79736
rect 156880 79688 156932 79694
rect 156880 79630 156932 79636
rect 157156 79688 157208 79694
rect 157444 79665 157472 79766
rect 157582 79744 157610 80036
rect 157674 79966 157702 80036
rect 157766 79966 157794 80036
rect 157662 79960 157714 79966
rect 157662 79902 157714 79908
rect 157754 79960 157806 79966
rect 157754 79902 157806 79908
rect 157858 79898 157886 80036
rect 157950 79966 157978 80036
rect 157938 79960 157990 79966
rect 157938 79902 157990 79908
rect 158042 79898 158070 80036
rect 157846 79892 157898 79898
rect 157846 79834 157898 79840
rect 158030 79892 158082 79898
rect 158030 79834 158082 79840
rect 157708 79824 157760 79830
rect 158134 79801 158162 80036
rect 158226 79830 158254 80036
rect 158214 79824 158266 79830
rect 157708 79766 157760 79772
rect 158120 79792 158176 79801
rect 157582 79716 157656 79744
rect 157156 79630 157208 79636
rect 157430 79656 157486 79665
rect 156788 79620 156840 79626
rect 156788 79562 156840 79568
rect 156432 77574 156736 77602
rect 156328 76628 156380 76634
rect 156328 76570 156380 76576
rect 156328 75132 156380 75138
rect 156328 75074 156380 75080
rect 156340 50658 156368 75074
rect 156432 54534 156460 77574
rect 156604 77376 156656 77382
rect 156604 77318 156656 77324
rect 156512 76628 156564 76634
rect 156512 76570 156564 76576
rect 156524 57254 156552 76570
rect 156616 65686 156644 77318
rect 156800 75138 156828 79562
rect 156892 76702 156920 79630
rect 157064 79620 157116 79626
rect 157064 79562 157116 79568
rect 156972 79552 157024 79558
rect 156972 79494 157024 79500
rect 156880 76696 156932 76702
rect 156880 76638 156932 76644
rect 156984 76106 157012 79494
rect 157076 77897 157104 79562
rect 157168 78713 157196 79630
rect 157430 79591 157486 79600
rect 157524 79620 157576 79626
rect 157524 79562 157576 79568
rect 157154 78704 157210 78713
rect 157154 78639 157210 78648
rect 157248 78328 157300 78334
rect 157248 78270 157300 78276
rect 157062 77888 157118 77897
rect 157062 77823 157118 77832
rect 157064 77648 157116 77654
rect 157064 77590 157116 77596
rect 156892 76078 157012 76106
rect 156892 75449 156920 76078
rect 156972 76016 157024 76022
rect 156972 75958 157024 75964
rect 156878 75440 156934 75449
rect 156878 75375 156934 75384
rect 156788 75132 156840 75138
rect 156788 75074 156840 75080
rect 156604 65680 156656 65686
rect 156604 65622 156656 65628
rect 156512 57248 156564 57254
rect 156512 57190 156564 57196
rect 156420 54528 156472 54534
rect 156420 54470 156472 54476
rect 156328 50652 156380 50658
rect 156328 50594 156380 50600
rect 156984 49230 157012 75958
rect 157076 68746 157104 77590
rect 157260 75478 157288 78270
rect 157340 78192 157392 78198
rect 157340 78134 157392 78140
rect 157248 75472 157300 75478
rect 157248 75414 157300 75420
rect 157064 68740 157116 68746
rect 157064 68682 157116 68688
rect 156972 49224 157024 49230
rect 156972 49166 157024 49172
rect 156236 46300 156288 46306
rect 156236 46242 156288 46248
rect 156604 46232 156656 46238
rect 156604 46174 156656 46180
rect 156144 19984 156196 19990
rect 156144 19926 156196 19932
rect 156052 14544 156104 14550
rect 156052 14486 156104 14492
rect 156144 11824 156196 11830
rect 156144 11766 156196 11772
rect 155960 6452 156012 6458
rect 155960 6394 156012 6400
rect 155408 3732 155460 3738
rect 155408 3674 155460 3680
rect 155224 3664 155276 3670
rect 155224 3606 155276 3612
rect 153844 3120 153896 3126
rect 153844 3062 153896 3068
rect 155420 480 155448 3674
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 11766
rect 156616 3738 156644 46174
rect 157352 9314 157380 78134
rect 157536 77294 157564 79562
rect 157628 77790 157656 79716
rect 157720 78198 157748 79766
rect 158214 79766 158266 79772
rect 158120 79727 158176 79736
rect 158318 79744 158346 80036
rect 158410 79971 158438 80036
rect 158396 79962 158452 79971
rect 158396 79897 158452 79906
rect 158502 79830 158530 80036
rect 158490 79824 158542 79830
rect 158594 79801 158622 80036
rect 158686 79971 158714 80036
rect 158672 79962 158728 79971
rect 158672 79897 158728 79906
rect 158778 79898 158806 80036
rect 158766 79892 158818 79898
rect 158766 79834 158818 79840
rect 158490 79766 158542 79772
rect 158580 79792 158636 79801
rect 158318 79716 158392 79744
rect 158580 79727 158636 79736
rect 158718 79792 158774 79801
rect 158718 79727 158720 79736
rect 157892 79688 157944 79694
rect 157892 79630 157944 79636
rect 158122 79688 158174 79694
rect 158364 79665 158392 79716
rect 158772 79727 158774 79736
rect 158870 79744 158898 80036
rect 158962 79812 158990 80036
rect 159054 79966 159082 80036
rect 159042 79960 159094 79966
rect 159042 79902 159094 79908
rect 158962 79784 159036 79812
rect 158870 79716 158944 79744
rect 158720 79698 158772 79704
rect 158444 79688 158496 79694
rect 158350 79656 158406 79665
rect 158174 79636 158208 79642
rect 158122 79630 158208 79636
rect 157800 79280 157852 79286
rect 157800 79222 157852 79228
rect 157812 79014 157840 79222
rect 157800 79008 157852 79014
rect 157800 78950 157852 78956
rect 157904 78690 157932 79630
rect 157984 79620 158036 79626
rect 158134 79614 158208 79630
rect 157984 79562 158036 79568
rect 157812 78662 157932 78690
rect 157708 78192 157760 78198
rect 157708 78134 157760 78140
rect 157708 77988 157760 77994
rect 157708 77930 157760 77936
rect 157616 77784 157668 77790
rect 157616 77726 157668 77732
rect 157536 77266 157656 77294
rect 157524 76696 157576 76702
rect 157524 76638 157576 76644
rect 157432 76628 157484 76634
rect 157432 76570 157484 76576
rect 157444 22914 157472 76570
rect 157536 76430 157564 76638
rect 157524 76424 157576 76430
rect 157524 76366 157576 76372
rect 157524 76288 157576 76294
rect 157524 76230 157576 76236
rect 157536 38010 157564 76230
rect 157628 39438 157656 77266
rect 157720 42158 157748 77930
rect 157812 51746 157840 78662
rect 157890 78432 157946 78441
rect 157890 78367 157946 78376
rect 157904 62898 157932 78367
rect 157996 77994 158024 79562
rect 158076 79552 158128 79558
rect 158076 79494 158128 79500
rect 157984 77988 158036 77994
rect 157984 77930 158036 77936
rect 157984 77308 158036 77314
rect 157984 77250 158036 77256
rect 157996 72554 158024 77250
rect 157984 72548 158036 72554
rect 157984 72490 158036 72496
rect 158088 64874 158116 79494
rect 158180 76634 158208 79614
rect 158444 79630 158496 79636
rect 158536 79688 158588 79694
rect 158588 79636 158668 79642
rect 158536 79630 158668 79636
rect 158350 79591 158406 79600
rect 158260 79552 158312 79558
rect 158260 79494 158312 79500
rect 158168 76628 158220 76634
rect 158168 76570 158220 76576
rect 158272 76294 158300 79494
rect 158352 79144 158404 79150
rect 158352 79086 158404 79092
rect 158364 77450 158392 79086
rect 158456 78962 158484 79630
rect 158548 79614 158668 79630
rect 158456 78934 158576 78962
rect 158352 77444 158404 77450
rect 158352 77386 158404 77392
rect 158548 77294 158576 78934
rect 158640 78334 158668 79614
rect 158812 79076 158864 79082
rect 158812 79018 158864 79024
rect 158824 78946 158852 79018
rect 158812 78940 158864 78946
rect 158812 78882 158864 78888
rect 158812 78668 158864 78674
rect 158812 78610 158864 78616
rect 158628 78328 158680 78334
rect 158628 78270 158680 78276
rect 158456 77266 158576 77294
rect 158260 76288 158312 76294
rect 158260 76230 158312 76236
rect 158456 70394 158484 77266
rect 158364 70366 158484 70394
rect 158364 65618 158392 70366
rect 158352 65612 158404 65618
rect 158352 65554 158404 65560
rect 157996 64846 158116 64874
rect 157996 64326 158024 64846
rect 157984 64320 158036 64326
rect 157984 64262 158036 64268
rect 157892 62892 157944 62898
rect 157892 62834 157944 62840
rect 157800 51740 157852 51746
rect 157800 51682 157852 51688
rect 157708 42152 157760 42158
rect 157708 42094 157760 42100
rect 157616 39432 157668 39438
rect 157616 39374 157668 39380
rect 157524 38004 157576 38010
rect 157524 37946 157576 37952
rect 157432 22908 157484 22914
rect 157432 22850 157484 22856
rect 158824 18766 158852 78610
rect 158916 29646 158944 79716
rect 159008 78674 159036 79784
rect 159146 79744 159174 80036
rect 159238 79937 159266 80036
rect 159224 79928 159280 79937
rect 159224 79863 159280 79872
rect 159330 79778 159358 80036
rect 159422 79898 159450 80036
rect 159514 79898 159542 80036
rect 159606 79898 159634 80036
rect 159698 79966 159726 80036
rect 159686 79960 159738 79966
rect 159686 79902 159738 79908
rect 159410 79892 159462 79898
rect 159410 79834 159462 79840
rect 159502 79892 159554 79898
rect 159502 79834 159554 79840
rect 159594 79892 159646 79898
rect 159594 79834 159646 79840
rect 159790 79778 159818 80036
rect 159882 79830 159910 80036
rect 159974 79937 160002 80036
rect 159960 79928 160016 79937
rect 160066 79898 160094 80036
rect 160158 79898 160186 80036
rect 159960 79863 160016 79872
rect 160054 79892 160106 79898
rect 160054 79834 160106 79840
rect 160146 79892 160198 79898
rect 160146 79834 160198 79840
rect 159284 79750 159358 79778
rect 159744 79750 159818 79778
rect 159870 79824 159922 79830
rect 159870 79766 159922 79772
rect 160098 79792 160154 79801
rect 159146 79716 159220 79744
rect 159088 79416 159140 79422
rect 159088 79358 159140 79364
rect 159100 78674 159128 79358
rect 158996 78668 159048 78674
rect 158996 78610 159048 78616
rect 159088 78668 159140 78674
rect 159088 78610 159140 78616
rect 158996 78328 159048 78334
rect 158996 78270 159048 78276
rect 159008 77217 159036 78270
rect 158994 77208 159050 77217
rect 158994 77143 159050 77152
rect 158994 76528 159050 76537
rect 158994 76463 159050 76472
rect 159008 47802 159036 76463
rect 159088 76220 159140 76226
rect 159088 76162 159140 76168
rect 159100 58818 159128 76162
rect 159192 76106 159220 79716
rect 159284 76226 159312 79750
rect 159364 79688 159416 79694
rect 159362 79656 159364 79665
rect 159416 79656 159418 79665
rect 159362 79591 159418 79600
rect 159456 79620 159508 79626
rect 159456 79562 159508 79568
rect 159548 79620 159600 79626
rect 159548 79562 159600 79568
rect 159364 79552 159416 79558
rect 159364 79494 159416 79500
rect 159376 79234 159404 79494
rect 159468 79370 159496 79562
rect 159560 79472 159588 79562
rect 159560 79444 159680 79472
rect 159468 79342 159588 79370
rect 159376 79206 159496 79234
rect 159364 79076 159416 79082
rect 159364 79018 159416 79024
rect 159376 78946 159404 79018
rect 159364 78940 159416 78946
rect 159364 78882 159416 78888
rect 159468 78810 159496 79206
rect 159456 78804 159508 78810
rect 159456 78746 159508 78752
rect 159362 78704 159418 78713
rect 159362 78639 159418 78648
rect 159272 76220 159324 76226
rect 159272 76162 159324 76168
rect 159192 76078 159312 76106
rect 159180 75268 159232 75274
rect 159180 75210 159232 75216
rect 159192 62830 159220 75210
rect 159284 68542 159312 76078
rect 159376 75177 159404 78639
rect 159560 78402 159588 79342
rect 159548 78396 159600 78402
rect 159548 78338 159600 78344
rect 159454 78160 159510 78169
rect 159454 78095 159510 78104
rect 159362 75168 159418 75177
rect 159362 75103 159418 75112
rect 159468 72486 159496 78095
rect 159456 72480 159508 72486
rect 159456 72422 159508 72428
rect 159652 70394 159680 79444
rect 159744 78305 159772 79750
rect 160098 79727 160154 79736
rect 159824 79688 159876 79694
rect 159824 79630 159876 79636
rect 159916 79688 159968 79694
rect 159916 79630 159968 79636
rect 159730 78296 159786 78305
rect 159730 78231 159786 78240
rect 159836 75274 159864 79630
rect 159928 75313 159956 79630
rect 160112 79506 160140 79727
rect 160250 79642 160278 80036
rect 160342 79744 160370 80036
rect 160434 79898 160462 80036
rect 160526 79937 160554 80036
rect 160512 79928 160568 79937
rect 160422 79892 160474 79898
rect 160512 79863 160568 79872
rect 160422 79834 160474 79840
rect 160618 79812 160646 80036
rect 160710 79966 160738 80036
rect 160698 79960 160750 79966
rect 160698 79902 160750 79908
rect 160802 79812 160830 80036
rect 160894 79966 160922 80036
rect 160986 79966 161014 80036
rect 161078 79971 161106 80036
rect 160882 79960 160934 79966
rect 160882 79902 160934 79908
rect 160974 79960 161026 79966
rect 160974 79902 161026 79908
rect 161064 79962 161120 79971
rect 161064 79897 161120 79906
rect 161170 79898 161198 80036
rect 161262 79937 161290 80036
rect 161354 79966 161382 80036
rect 161446 79966 161474 80036
rect 161538 79971 161566 80036
rect 161342 79960 161394 79966
rect 161248 79928 161304 79937
rect 161158 79892 161210 79898
rect 161342 79902 161394 79908
rect 161434 79960 161486 79966
rect 161434 79902 161486 79908
rect 161524 79962 161580 79971
rect 161524 79897 161580 79906
rect 161248 79863 161304 79872
rect 161158 79834 161210 79840
rect 161630 79812 161658 80036
rect 161722 79971 161750 80036
rect 161708 79962 161764 79971
rect 161814 79966 161842 80036
rect 161708 79897 161764 79906
rect 161802 79960 161854 79966
rect 161802 79902 161854 79908
rect 161906 79830 161934 80036
rect 161894 79824 161946 79830
rect 160618 79784 160692 79812
rect 160802 79784 160968 79812
rect 161630 79784 161796 79812
rect 160664 79778 160692 79784
rect 160468 79756 160520 79762
rect 160342 79716 160416 79744
rect 160250 79614 160324 79642
rect 160020 79478 160140 79506
rect 160020 78554 160048 79478
rect 160020 78526 160140 78554
rect 160008 78396 160060 78402
rect 160008 78338 160060 78344
rect 159914 75304 159970 75313
rect 159824 75268 159876 75274
rect 159914 75239 159970 75248
rect 159824 75210 159876 75216
rect 159376 70366 159680 70394
rect 159376 69970 159404 70366
rect 159364 69964 159416 69970
rect 159364 69906 159416 69912
rect 159272 68536 159324 68542
rect 159272 68478 159324 68484
rect 159180 62824 159232 62830
rect 159180 62766 159232 62772
rect 159088 58812 159140 58818
rect 159088 58754 159140 58760
rect 158996 47796 159048 47802
rect 158996 47738 159048 47744
rect 158904 29640 158956 29646
rect 158904 29582 158956 29588
rect 158812 18760 158864 18766
rect 158812 18702 158864 18708
rect 160020 11966 160048 78338
rect 160112 77654 160140 78526
rect 160190 78432 160246 78441
rect 160190 78367 160246 78376
rect 160100 77648 160152 77654
rect 160100 77590 160152 77596
rect 160100 75948 160152 75954
rect 160100 75890 160152 75896
rect 160008 11960 160060 11966
rect 160008 11902 160060 11908
rect 160112 11898 160140 75890
rect 160204 16114 160232 78367
rect 160296 75834 160324 79614
rect 160388 75954 160416 79716
rect 160664 79750 160738 79778
rect 160710 79744 160738 79750
rect 160710 79716 160876 79744
rect 160468 79698 160520 79704
rect 160480 75954 160508 79698
rect 160560 79620 160612 79626
rect 160560 79562 160612 79568
rect 160744 79620 160796 79626
rect 160744 79562 160796 79568
rect 160376 75948 160428 75954
rect 160376 75890 160428 75896
rect 160468 75948 160520 75954
rect 160468 75890 160520 75896
rect 160296 75806 160508 75834
rect 160284 75336 160336 75342
rect 160284 75278 160336 75284
rect 160192 16108 160244 16114
rect 160192 16050 160244 16056
rect 160296 16046 160324 75278
rect 160376 75268 160428 75274
rect 160376 75210 160428 75216
rect 160388 17406 160416 75210
rect 160480 17474 160508 75806
rect 160572 47734 160600 79562
rect 160652 79552 160704 79558
rect 160652 79494 160704 79500
rect 160664 77314 160692 79494
rect 160652 77308 160704 77314
rect 160652 77250 160704 77256
rect 160652 75948 160704 75954
rect 160652 75890 160704 75896
rect 160664 50590 160692 75890
rect 160756 53242 160784 79562
rect 160848 78878 160876 79716
rect 160836 78872 160888 78878
rect 160836 78814 160888 78820
rect 160836 78396 160888 78402
rect 160836 78338 160888 78344
rect 160848 75342 160876 78338
rect 160836 75336 160888 75342
rect 160836 75278 160888 75284
rect 160940 75274 160968 79784
rect 161112 79756 161164 79762
rect 161112 79698 161164 79704
rect 161204 79756 161256 79762
rect 161204 79698 161256 79704
rect 161020 79688 161072 79694
rect 161020 79630 161072 79636
rect 161032 78402 161060 79630
rect 161124 78402 161152 79698
rect 161216 79150 161244 79698
rect 161572 79688 161624 79694
rect 161492 79648 161572 79676
rect 161388 79552 161440 79558
rect 161388 79494 161440 79500
rect 161296 79416 161348 79422
rect 161296 79358 161348 79364
rect 161204 79144 161256 79150
rect 161204 79086 161256 79092
rect 161204 78872 161256 78878
rect 161204 78814 161256 78820
rect 161020 78396 161072 78402
rect 161020 78338 161072 78344
rect 161112 78396 161164 78402
rect 161112 78338 161164 78344
rect 161020 78260 161072 78266
rect 161020 78202 161072 78208
rect 160928 75268 160980 75274
rect 160928 75210 160980 75216
rect 160834 75168 160890 75177
rect 160834 75103 160890 75112
rect 160848 64258 160876 75103
rect 161032 70394 161060 78202
rect 161110 77480 161166 77489
rect 161110 77415 161166 77424
rect 161124 77382 161152 77415
rect 161112 77376 161164 77382
rect 161112 77318 161164 77324
rect 161216 77217 161244 78814
rect 161308 78674 161336 79358
rect 161296 78668 161348 78674
rect 161296 78610 161348 78616
rect 161202 77208 161258 77217
rect 161202 77143 161258 77152
rect 161400 76401 161428 79494
rect 161386 76392 161442 76401
rect 161386 76327 161442 76336
rect 161492 75313 161520 79648
rect 161572 79630 161624 79636
rect 161572 79484 161624 79490
rect 161572 79426 161624 79432
rect 161664 79484 161716 79490
rect 161664 79426 161716 79432
rect 161584 79286 161612 79426
rect 161572 79280 161624 79286
rect 161572 79222 161624 79228
rect 161572 79144 161624 79150
rect 161572 79086 161624 79092
rect 161584 76090 161612 79086
rect 161572 76084 161624 76090
rect 161572 76026 161624 76032
rect 161570 75984 161626 75993
rect 161570 75919 161626 75928
rect 161478 75304 161534 75313
rect 161478 75239 161534 75248
rect 161480 73432 161532 73438
rect 161480 73374 161532 73380
rect 161032 70366 161152 70394
rect 160836 64252 160888 64258
rect 160836 64194 160888 64200
rect 161124 60042 161152 70366
rect 161112 60036 161164 60042
rect 161112 59978 161164 59984
rect 160744 53236 160796 53242
rect 160744 53178 160796 53184
rect 160652 50584 160704 50590
rect 160652 50526 160704 50532
rect 160742 50280 160798 50289
rect 160742 50215 160798 50224
rect 160560 47728 160612 47734
rect 160560 47670 160612 47676
rect 160468 17468 160520 17474
rect 160468 17410 160520 17416
rect 160376 17400 160428 17406
rect 160376 17342 160428 17348
rect 160284 16040 160336 16046
rect 160284 15982 160336 15988
rect 160100 11892 160152 11898
rect 160100 11834 160152 11840
rect 157340 9308 157392 9314
rect 157340 9250 157392 9256
rect 158902 4856 158958 4865
rect 157800 4820 157852 4826
rect 158902 4791 158958 4800
rect 157800 4762 157852 4768
rect 156604 3732 156656 3738
rect 156604 3674 156656 3680
rect 157812 480 157840 4762
rect 158916 480 158944 4791
rect 160756 3670 160784 50215
rect 161492 6322 161520 73374
rect 161584 6390 161612 75919
rect 161676 9246 161704 79426
rect 161768 76158 161796 79784
rect 161894 79766 161946 79772
rect 161998 79778 162026 80036
rect 162090 79898 162118 80036
rect 162182 79966 162210 80036
rect 162170 79960 162222 79966
rect 162170 79902 162222 79908
rect 162274 79898 162302 80036
rect 162078 79892 162130 79898
rect 162078 79834 162130 79840
rect 162262 79892 162314 79898
rect 162262 79834 162314 79840
rect 161998 79750 162072 79778
rect 161848 79688 161900 79694
rect 161848 79630 161900 79636
rect 161756 76152 161808 76158
rect 161756 76094 161808 76100
rect 161756 76016 161808 76022
rect 161756 75958 161808 75964
rect 161664 9240 161716 9246
rect 161664 9182 161716 9188
rect 161768 9178 161796 75958
rect 161860 73438 161888 79630
rect 161940 79552 161992 79558
rect 161940 79494 161992 79500
rect 161952 79150 161980 79494
rect 161940 79144 161992 79150
rect 161940 79086 161992 79092
rect 161940 76288 161992 76294
rect 161940 76230 161992 76236
rect 161848 73432 161900 73438
rect 161848 73374 161900 73380
rect 161848 73296 161900 73302
rect 161848 73238 161900 73244
rect 161756 9172 161808 9178
rect 161756 9114 161808 9120
rect 161860 9110 161888 73238
rect 161952 11762 161980 76230
rect 162044 72894 162072 79750
rect 162366 79744 162394 80036
rect 162458 79830 162486 80036
rect 162446 79824 162498 79830
rect 162446 79766 162498 79772
rect 162228 79716 162394 79744
rect 162228 79608 162256 79716
rect 162550 79676 162578 80036
rect 162642 79966 162670 80036
rect 162630 79960 162682 79966
rect 162630 79902 162682 79908
rect 162734 79801 162762 80036
rect 162720 79792 162776 79801
rect 162826 79778 162854 80036
rect 162918 79937 162946 80036
rect 162904 79928 162960 79937
rect 162904 79863 162960 79872
rect 163010 79812 163038 80036
rect 162964 79801 163038 79812
rect 162950 79792 163038 79801
rect 162826 79750 162900 79778
rect 162720 79727 162776 79736
rect 162504 79648 162578 79676
rect 162676 79688 162728 79694
rect 162400 79620 162452 79626
rect 162228 79580 162348 79608
rect 162124 79484 162176 79490
rect 162124 79426 162176 79432
rect 162136 76294 162164 79426
rect 162216 79144 162268 79150
rect 162216 79086 162268 79092
rect 162228 78130 162256 79086
rect 162216 78124 162268 78130
rect 162216 78066 162268 78072
rect 162216 77240 162268 77246
rect 162216 77182 162268 77188
rect 162228 76498 162256 77182
rect 162216 76492 162268 76498
rect 162216 76434 162268 76440
rect 162124 76288 162176 76294
rect 162124 76230 162176 76236
rect 162124 76152 162176 76158
rect 162124 76094 162176 76100
rect 162032 72888 162084 72894
rect 162032 72830 162084 72836
rect 162136 70394 162164 76094
rect 162320 73302 162348 79580
rect 162504 79608 162532 79648
rect 162676 79630 162728 79636
rect 162768 79688 162820 79694
rect 162768 79630 162820 79636
rect 162504 79580 162624 79608
rect 162400 79562 162452 79568
rect 162412 79121 162440 79562
rect 162492 79484 162544 79490
rect 162492 79426 162544 79432
rect 162398 79112 162454 79121
rect 162398 79047 162454 79056
rect 162400 78736 162452 78742
rect 162400 78678 162452 78684
rect 162308 73296 162360 73302
rect 162308 73238 162360 73244
rect 162044 70366 162164 70394
rect 162044 11830 162072 70366
rect 162412 70038 162440 78678
rect 162504 76362 162532 79426
rect 162596 78334 162624 79580
rect 162584 78328 162636 78334
rect 162584 78270 162636 78276
rect 162492 76356 162544 76362
rect 162492 76298 162544 76304
rect 162688 75041 162716 79630
rect 162674 75032 162730 75041
rect 162674 74967 162730 74976
rect 162780 70394 162808 79630
rect 162872 77294 162900 79750
rect 163006 79784 163038 79792
rect 162950 79727 163006 79736
rect 163102 79744 163130 80036
rect 163194 79898 163222 80036
rect 163182 79892 163234 79898
rect 163182 79834 163234 79840
rect 163286 79830 163314 80036
rect 163378 79966 163406 80036
rect 163366 79960 163418 79966
rect 163366 79902 163418 79908
rect 163274 79824 163326 79830
rect 163274 79766 163326 79772
rect 163470 79744 163498 80036
rect 163562 79830 163590 80036
rect 163654 79966 163682 80036
rect 163746 79966 163774 80036
rect 163642 79960 163694 79966
rect 163642 79902 163694 79908
rect 163734 79960 163786 79966
rect 163734 79902 163786 79908
rect 163838 79898 163866 80036
rect 163826 79892 163878 79898
rect 163826 79834 163878 79840
rect 163550 79824 163602 79830
rect 163550 79766 163602 79772
rect 163930 79778 163958 80036
rect 164022 79937 164050 80036
rect 164008 79928 164064 79937
rect 164008 79863 164064 79872
rect 164114 79801 164142 80036
rect 164206 79898 164234 80036
rect 164298 79966 164326 80036
rect 164286 79960 164338 79966
rect 164286 79902 164338 79908
rect 164194 79892 164246 79898
rect 164194 79834 164246 79840
rect 164100 79792 164156 79801
rect 163102 79716 163176 79744
rect 163042 79656 163098 79665
rect 163042 79591 163098 79600
rect 162872 77266 162992 77294
rect 162964 75721 162992 77266
rect 162950 75712 163006 75721
rect 162950 75647 163006 75656
rect 163056 75614 163084 79591
rect 163148 78130 163176 79716
rect 163424 79716 163498 79744
rect 163780 79756 163832 79762
rect 163228 79688 163280 79694
rect 163228 79630 163280 79636
rect 163320 79688 163372 79694
rect 163320 79630 163372 79636
rect 163136 78124 163188 78130
rect 163136 78066 163188 78072
rect 163136 76016 163188 76022
rect 163136 75958 163188 75964
rect 163044 75608 163096 75614
rect 163044 75550 163096 75556
rect 162952 75404 163004 75410
rect 162952 75346 163004 75352
rect 162780 70366 162900 70394
rect 162400 70032 162452 70038
rect 162400 69974 162452 69980
rect 162032 11824 162084 11830
rect 162032 11766 162084 11772
rect 161940 11756 161992 11762
rect 161940 11698 161992 11704
rect 161848 9104 161900 9110
rect 161848 9046 161900 9052
rect 161572 6384 161624 6390
rect 161572 6326 161624 6332
rect 161480 6316 161532 6322
rect 161480 6258 161532 6264
rect 162872 4894 162900 70366
rect 162964 17338 162992 75346
rect 163044 75268 163096 75274
rect 163044 75210 163096 75216
rect 163056 35222 163084 75210
rect 163148 46238 163176 75958
rect 163240 47666 163268 79630
rect 163332 53174 163360 79630
rect 163424 78316 163452 79716
rect 163930 79750 164004 79778
rect 163780 79698 163832 79704
rect 163686 79656 163742 79665
rect 163596 79620 163648 79626
rect 163686 79591 163742 79600
rect 163596 79562 163648 79568
rect 163608 78441 163636 79562
rect 163594 78432 163650 78441
rect 163594 78367 163650 78376
rect 163424 78288 163636 78316
rect 163504 78124 163556 78130
rect 163504 78066 163556 78072
rect 163412 75608 163464 75614
rect 163412 75550 163464 75556
rect 163424 61470 163452 75550
rect 163516 68474 163544 78066
rect 163608 75274 163636 78288
rect 163700 78198 163728 79591
rect 163688 78192 163740 78198
rect 163688 78134 163740 78140
rect 163596 75268 163648 75274
rect 163596 75210 163648 75216
rect 163792 72962 163820 79698
rect 163872 79688 163924 79694
rect 163872 79630 163924 79636
rect 163884 76022 163912 79630
rect 163872 76016 163924 76022
rect 163872 75958 163924 75964
rect 163976 75410 164004 79750
rect 164390 79778 164418 80036
rect 164482 79812 164510 80036
rect 164574 79966 164602 80036
rect 164562 79960 164614 79966
rect 164562 79902 164614 79908
rect 164666 79903 164694 80036
rect 164758 79966 164786 80036
rect 164746 79960 164798 79966
rect 164652 79894 164708 79903
rect 164746 79902 164798 79908
rect 164652 79829 164708 79838
rect 164482 79784 164556 79812
rect 164100 79727 164156 79736
rect 164344 79750 164418 79778
rect 164238 79656 164294 79665
rect 164148 79620 164200 79626
rect 164238 79591 164294 79600
rect 164148 79562 164200 79568
rect 164056 79552 164108 79558
rect 164056 79494 164108 79500
rect 163964 75404 164016 75410
rect 163964 75346 164016 75352
rect 164068 74186 164096 79494
rect 164160 75410 164188 79562
rect 164148 75404 164200 75410
rect 164148 75346 164200 75352
rect 164056 74180 164108 74186
rect 164056 74122 164108 74128
rect 163780 72956 163832 72962
rect 163780 72898 163832 72904
rect 163504 68468 163556 68474
rect 163504 68410 163556 68416
rect 163412 61464 163464 61470
rect 163412 61406 163464 61412
rect 163320 53168 163372 53174
rect 163320 53110 163372 53116
rect 163228 47660 163280 47666
rect 163228 47602 163280 47608
rect 163136 46232 163188 46238
rect 163136 46174 163188 46180
rect 163044 35216 163096 35222
rect 163044 35158 163096 35164
rect 162952 17332 163004 17338
rect 162952 17274 163004 17280
rect 164252 6254 164280 79591
rect 164344 75342 164372 79750
rect 164424 79688 164476 79694
rect 164422 79656 164424 79665
rect 164476 79656 164478 79665
rect 164422 79591 164478 79600
rect 164424 79552 164476 79558
rect 164424 79494 164476 79500
rect 164436 79286 164464 79494
rect 164424 79280 164476 79286
rect 164424 79222 164476 79228
rect 164422 77616 164478 77625
rect 164422 77551 164478 77560
rect 164436 77450 164464 77551
rect 164424 77444 164476 77450
rect 164424 77386 164476 77392
rect 164332 75336 164384 75342
rect 164332 75278 164384 75284
rect 164424 75200 164476 75206
rect 164424 75142 164476 75148
rect 164332 75132 164384 75138
rect 164332 75074 164384 75080
rect 164344 7614 164372 75074
rect 164436 9042 164464 75142
rect 164528 31210 164556 79784
rect 164850 79778 164878 80036
rect 164942 79830 164970 80036
rect 164700 79756 164752 79762
rect 164620 79716 164700 79744
rect 164620 37942 164648 79716
rect 164700 79698 164752 79704
rect 164804 79750 164878 79778
rect 164930 79824 164982 79830
rect 164930 79766 164982 79772
rect 165034 79778 165062 80036
rect 165126 79898 165154 80036
rect 165114 79892 165166 79898
rect 165114 79834 165166 79840
rect 165218 79830 165246 80036
rect 165310 79898 165338 80036
rect 165402 79966 165430 80036
rect 165494 79966 165522 80036
rect 165390 79960 165442 79966
rect 165390 79902 165442 79908
rect 165482 79960 165534 79966
rect 165586 79937 165614 80036
rect 165678 79966 165706 80036
rect 165770 79971 165798 80036
rect 165666 79960 165718 79966
rect 165482 79902 165534 79908
rect 165572 79928 165628 79937
rect 165298 79892 165350 79898
rect 165666 79902 165718 79908
rect 165756 79962 165812 79971
rect 165862 79966 165890 80036
rect 165756 79897 165812 79906
rect 165850 79960 165902 79966
rect 165850 79902 165902 79908
rect 165572 79863 165628 79872
rect 165298 79834 165350 79840
rect 165206 79824 165258 79830
rect 165034 79750 165108 79778
rect 165482 79824 165534 79830
rect 165206 79766 165258 79772
rect 165480 79792 165482 79801
rect 165712 79824 165764 79830
rect 165534 79792 165536 79801
rect 164700 79280 164752 79286
rect 164700 79222 164752 79228
rect 164712 79082 164740 79222
rect 164700 79076 164752 79082
rect 164700 79018 164752 79024
rect 164804 78928 164832 79750
rect 164884 79688 164936 79694
rect 164884 79630 164936 79636
rect 164974 79656 165030 79665
rect 164712 78900 164832 78928
rect 164712 75682 164740 78900
rect 164790 78704 164846 78713
rect 164790 78639 164846 78648
rect 164804 78266 164832 78639
rect 164792 78260 164844 78266
rect 164792 78202 164844 78208
rect 164700 75676 164752 75682
rect 164700 75618 164752 75624
rect 164700 75336 164752 75342
rect 164700 75278 164752 75284
rect 164712 49094 164740 75278
rect 164896 75138 164924 79630
rect 164974 79591 164976 79600
rect 165028 79591 165030 79600
rect 164976 79562 165028 79568
rect 165080 79472 165108 79750
rect 165954 79812 165982 80036
rect 166046 79966 166074 80036
rect 166034 79960 166086 79966
rect 166034 79902 166086 79908
rect 166138 79830 166166 80036
rect 165712 79766 165764 79772
rect 165816 79784 165982 79812
rect 166126 79824 166178 79830
rect 165480 79727 165536 79736
rect 165252 79688 165304 79694
rect 165252 79630 165304 79636
rect 165528 79688 165580 79694
rect 165528 79630 165580 79636
rect 165160 79620 165212 79626
rect 165160 79562 165212 79568
rect 164988 79444 165108 79472
rect 164988 78713 165016 79444
rect 165172 78826 165200 79562
rect 165080 78798 165200 78826
rect 164974 78704 165030 78713
rect 164974 78639 165030 78648
rect 164976 78600 165028 78606
rect 164976 78542 165028 78548
rect 164988 75206 165016 78542
rect 164976 75200 165028 75206
rect 164976 75142 165028 75148
rect 164884 75132 164936 75138
rect 164884 75074 164936 75080
rect 165080 70394 165108 78798
rect 165158 78704 165214 78713
rect 165158 78639 165214 78648
rect 165172 75138 165200 78639
rect 165264 78606 165292 79630
rect 165436 79620 165488 79626
rect 165436 79562 165488 79568
rect 165252 78600 165304 78606
rect 165252 78542 165304 78548
rect 165448 75993 165476 79562
rect 165434 75984 165490 75993
rect 165434 75919 165490 75928
rect 165252 75676 165304 75682
rect 165252 75618 165304 75624
rect 165160 75132 165212 75138
rect 165160 75074 165212 75080
rect 165264 71194 165292 75618
rect 165540 71774 165568 79630
rect 165618 79384 165674 79393
rect 165618 79319 165674 79328
rect 165632 79121 165660 79319
rect 165618 79112 165674 79121
rect 165618 79047 165674 79056
rect 165540 71746 165660 71774
rect 165252 71188 165304 71194
rect 165252 71130 165304 71136
rect 164804 70366 165108 70394
rect 164804 58750 164832 70366
rect 164792 58744 164844 58750
rect 164792 58686 164844 58692
rect 164700 49088 164752 49094
rect 164700 49030 164752 49036
rect 164608 37936 164660 37942
rect 164608 37878 164660 37884
rect 164516 31204 164568 31210
rect 164516 31146 164568 31152
rect 165632 14482 165660 71746
rect 165724 15978 165752 79766
rect 165816 75954 165844 79784
rect 166126 79766 166178 79772
rect 165896 79688 165948 79694
rect 166230 79676 166258 80036
rect 166322 79830 166350 80036
rect 166414 79937 166442 80036
rect 166400 79928 166456 79937
rect 166400 79863 166456 79872
rect 166310 79824 166362 79830
rect 166506 79778 166534 80036
rect 166598 79937 166626 80036
rect 166584 79928 166640 79937
rect 166584 79863 166640 79872
rect 166690 79778 166718 80036
rect 166310 79766 166362 79772
rect 166460 79750 166534 79778
rect 166644 79750 166718 79778
rect 165896 79630 165948 79636
rect 166078 79656 166134 79665
rect 165804 75948 165856 75954
rect 165804 75890 165856 75896
rect 165804 75200 165856 75206
rect 165804 75142 165856 75148
rect 165712 15972 165764 15978
rect 165712 15914 165764 15920
rect 165816 15910 165844 75142
rect 165908 22846 165936 79630
rect 166230 79648 166396 79676
rect 166078 79591 166134 79600
rect 166092 79472 166120 79591
rect 166092 79444 166212 79472
rect 166078 79384 166134 79393
rect 166078 79319 166134 79328
rect 165986 79248 166042 79257
rect 165986 79183 166042 79192
rect 166000 78878 166028 79183
rect 165988 78872 166040 78878
rect 165988 78814 166040 78820
rect 165986 78568 166042 78577
rect 165986 78503 166042 78512
rect 166000 78062 166028 78503
rect 165988 78056 166040 78062
rect 165988 77998 166040 78004
rect 165986 77888 166042 77897
rect 165986 77823 166042 77832
rect 166000 77625 166028 77823
rect 165986 77616 166042 77625
rect 165986 77551 166042 77560
rect 166092 77500 166120 79319
rect 166000 77472 166120 77500
rect 166000 24138 166028 77472
rect 166080 75336 166132 75342
rect 166080 75278 166132 75284
rect 166092 39370 166120 75278
rect 166184 53106 166212 79444
rect 166262 79248 166318 79257
rect 166262 79183 166318 79192
rect 166276 79014 166304 79183
rect 166264 79008 166316 79014
rect 166264 78950 166316 78956
rect 166264 78668 166316 78674
rect 166264 78610 166316 78616
rect 166276 78169 166304 78610
rect 166262 78160 166318 78169
rect 166262 78095 166318 78104
rect 166264 75268 166316 75274
rect 166264 75210 166316 75216
rect 166276 66910 166304 75210
rect 166368 69902 166396 79648
rect 166460 75274 166488 79750
rect 166540 79688 166592 79694
rect 166540 79630 166592 79636
rect 166448 75268 166500 75274
rect 166448 75210 166500 75216
rect 166552 75206 166580 79630
rect 166644 77489 166672 79750
rect 166782 79744 166810 80036
rect 166874 79898 166902 80036
rect 166966 79937 166994 80036
rect 166952 79928 167008 79937
rect 166862 79892 166914 79898
rect 166952 79863 167008 79872
rect 166862 79834 166914 79840
rect 167058 79812 167086 80036
rect 167012 79784 167086 79812
rect 166782 79716 166948 79744
rect 166722 79656 166778 79665
rect 166722 79591 166778 79600
rect 166816 79620 166868 79626
rect 166630 77480 166686 77489
rect 166630 77415 166686 77424
rect 166632 75948 166684 75954
rect 166632 75890 166684 75896
rect 166540 75200 166592 75206
rect 166540 75142 166592 75148
rect 166644 71126 166672 75890
rect 166736 75342 166764 79591
rect 166816 79562 166868 79568
rect 166828 77353 166856 79562
rect 166920 77897 166948 79716
rect 167012 78713 167040 79784
rect 167150 79744 167178 80036
rect 167242 79830 167270 80036
rect 167230 79824 167282 79830
rect 167334 79812 167362 80036
rect 167426 79966 167454 80036
rect 167414 79960 167466 79966
rect 167414 79902 167466 79908
rect 167334 79784 167408 79812
rect 167230 79766 167282 79772
rect 167104 79716 167178 79744
rect 166998 78704 167054 78713
rect 166998 78639 167054 78648
rect 167000 78600 167052 78606
rect 167000 78542 167052 78548
rect 166906 77888 166962 77897
rect 166906 77823 166962 77832
rect 167012 77518 167040 78542
rect 167000 77512 167052 77518
rect 167000 77454 167052 77460
rect 166814 77344 166870 77353
rect 166814 77279 166870 77288
rect 166908 77308 166960 77314
rect 166908 77250 166960 77256
rect 166920 75410 166948 77250
rect 166908 75404 166960 75410
rect 166908 75346 166960 75352
rect 166724 75336 166776 75342
rect 166724 75278 166776 75284
rect 167104 75070 167132 79716
rect 167276 79688 167328 79694
rect 167182 79656 167238 79665
rect 167276 79630 167328 79636
rect 167182 79591 167238 79600
rect 167196 78792 167224 79591
rect 167288 78860 167316 79630
rect 167380 79014 167408 79784
rect 167518 79744 167546 80036
rect 167610 79898 167638 80036
rect 167702 79937 167730 80036
rect 167688 79928 167744 79937
rect 167598 79892 167650 79898
rect 167688 79863 167744 79872
rect 167598 79834 167650 79840
rect 167794 79812 167822 80036
rect 167886 79830 167914 80036
rect 167748 79784 167822 79812
rect 167874 79824 167926 79830
rect 167518 79716 167592 79744
rect 167460 79620 167512 79626
rect 167460 79562 167512 79568
rect 167368 79008 167420 79014
rect 167368 78950 167420 78956
rect 167288 78832 167408 78860
rect 167196 78764 167316 78792
rect 167182 78704 167238 78713
rect 167182 78639 167238 78648
rect 167196 78130 167224 78639
rect 167184 78124 167236 78130
rect 167184 78066 167236 78072
rect 167182 75984 167238 75993
rect 167182 75919 167238 75928
rect 167092 75064 167144 75070
rect 167092 75006 167144 75012
rect 167092 74928 167144 74934
rect 167092 74870 167144 74876
rect 166632 71120 166684 71126
rect 166632 71062 166684 71068
rect 166356 69896 166408 69902
rect 166356 69838 166408 69844
rect 166264 66904 166316 66910
rect 166264 66846 166316 66852
rect 166172 53100 166224 53106
rect 166172 53042 166224 53048
rect 166080 39364 166132 39370
rect 166080 39306 166132 39312
rect 165988 24132 166040 24138
rect 165988 24074 166040 24080
rect 165896 22840 165948 22846
rect 165896 22782 165948 22788
rect 165804 15904 165856 15910
rect 165804 15846 165856 15852
rect 165620 14476 165672 14482
rect 165620 14418 165672 14424
rect 166080 10328 166132 10334
rect 166080 10270 166132 10276
rect 164424 9036 164476 9042
rect 164424 8978 164476 8984
rect 164332 7608 164384 7614
rect 164332 7550 164384 7556
rect 164240 6248 164292 6254
rect 164240 6190 164292 6196
rect 162860 4888 162912 4894
rect 162860 4830 162912 4836
rect 160100 3664 160152 3670
rect 160100 3606 160152 3612
rect 160744 3664 160796 3670
rect 160744 3606 160796 3612
rect 160112 480 160140 3606
rect 162492 3596 162544 3602
rect 162492 3538 162544 3544
rect 161296 3120 161348 3126
rect 161296 3062 161348 3068
rect 161308 480 161336 3062
rect 162504 480 162532 3538
rect 163688 3528 163740 3534
rect 163688 3470 163740 3476
rect 163700 480 163728 3470
rect 164882 3360 164938 3369
rect 164882 3295 164938 3304
rect 164896 480 164924 3295
rect 166092 480 166120 10270
rect 167104 6186 167132 74870
rect 167196 8974 167224 75919
rect 167288 17270 167316 78764
rect 167380 31142 167408 78832
rect 167472 76090 167500 79562
rect 167564 79393 167592 79716
rect 167550 79384 167606 79393
rect 167550 79319 167606 79328
rect 167748 79200 167776 79784
rect 167874 79766 167926 79772
rect 167828 79688 167880 79694
rect 167978 79676 168006 80036
rect 167828 79630 167880 79636
rect 167932 79648 168006 79676
rect 167564 79172 167776 79200
rect 167460 76084 167512 76090
rect 167460 76026 167512 76032
rect 167564 75970 167592 79172
rect 167840 79098 167868 79630
rect 167472 75942 167592 75970
rect 167656 79070 167868 79098
rect 167472 50454 167500 75942
rect 167552 75064 167604 75070
rect 167552 75006 167604 75012
rect 167564 50522 167592 75006
rect 167656 68406 167684 79070
rect 167736 79008 167788 79014
rect 167736 78950 167788 78956
rect 167748 69834 167776 78950
rect 167932 76242 167960 79648
rect 168070 79472 168098 80036
rect 168162 79937 168190 80036
rect 168254 79966 168282 80036
rect 168242 79960 168294 79966
rect 168148 79928 168204 79937
rect 168242 79902 168294 79908
rect 168148 79863 168204 79872
rect 168196 79824 168248 79830
rect 168346 79801 168374 80036
rect 168438 79971 168466 80036
rect 168424 79962 168480 79971
rect 168424 79897 168480 79906
rect 168196 79766 168248 79772
rect 168332 79792 168388 79801
rect 168024 79444 168098 79472
rect 168024 79393 168052 79444
rect 168010 79384 168066 79393
rect 168010 79319 168066 79328
rect 168010 78704 168066 78713
rect 168010 78639 168066 78648
rect 168024 78169 168052 78639
rect 168010 78160 168066 78169
rect 168010 78095 168066 78104
rect 167840 76214 167960 76242
rect 167840 74934 167868 76214
rect 167920 76084 167972 76090
rect 167920 76026 167972 76032
rect 167828 74928 167880 74934
rect 167828 74870 167880 74876
rect 167932 70394 167960 76026
rect 168208 75993 168236 79766
rect 168530 79744 168558 80036
rect 168332 79727 168388 79736
rect 168484 79716 168558 79744
rect 168622 79744 168650 80036
rect 168714 79966 168742 80036
rect 168702 79960 168754 79966
rect 168702 79902 168754 79908
rect 168806 79744 168834 80036
rect 168898 79966 168926 80036
rect 168990 79971 169018 80036
rect 168886 79960 168938 79966
rect 168886 79902 168938 79908
rect 168976 79962 169032 79971
rect 168976 79897 169032 79906
rect 169082 79812 169110 80036
rect 169174 79898 169202 80036
rect 169162 79892 169214 79898
rect 169162 79834 169214 79840
rect 168622 79716 168696 79744
rect 168288 79688 168340 79694
rect 168288 79630 168340 79636
rect 168380 79688 168432 79694
rect 168380 79630 168432 79636
rect 168194 75984 168250 75993
rect 168194 75919 168250 75928
rect 168300 71058 168328 79630
rect 168288 71052 168340 71058
rect 168288 70994 168340 71000
rect 167932 70366 168328 70394
rect 167736 69828 167788 69834
rect 167736 69770 167788 69776
rect 167644 68400 167696 68406
rect 167644 68342 167696 68348
rect 167552 50516 167604 50522
rect 167552 50458 167604 50464
rect 167460 50448 167512 50454
rect 167460 50390 167512 50396
rect 167368 31136 167420 31142
rect 167368 31078 167420 31084
rect 167276 17264 167328 17270
rect 167276 17206 167328 17212
rect 167184 8968 167236 8974
rect 167184 8910 167236 8916
rect 167092 6180 167144 6186
rect 167092 6122 167144 6128
rect 167184 5024 167236 5030
rect 167184 4966 167236 4972
rect 167196 480 167224 4966
rect 168300 4826 168328 70366
rect 168392 18698 168420 79630
rect 168484 75274 168512 79716
rect 168668 79393 168696 79716
rect 168760 79716 168834 79744
rect 168944 79784 169110 79812
rect 168654 79384 168710 79393
rect 168654 79319 168710 79328
rect 168760 78384 168788 79716
rect 168944 79472 168972 79784
rect 169266 79744 169294 80036
rect 169358 79830 169386 80036
rect 169450 79830 169478 80036
rect 169542 79898 169570 80036
rect 169634 79898 169662 80036
rect 169726 79937 169754 80036
rect 169712 79928 169768 79937
rect 169530 79892 169582 79898
rect 169530 79834 169582 79840
rect 169622 79892 169674 79898
rect 169712 79863 169768 79872
rect 169622 79834 169674 79840
rect 169346 79824 169398 79830
rect 169346 79766 169398 79772
rect 169438 79824 169490 79830
rect 169438 79766 169490 79772
rect 169818 79744 169846 80036
rect 169910 79971 169938 80036
rect 169896 79962 169952 79971
rect 170002 79966 170030 80036
rect 170094 79966 170122 80036
rect 170186 79966 170214 80036
rect 169896 79897 169952 79906
rect 169990 79960 170042 79966
rect 169990 79902 170042 79908
rect 170082 79960 170134 79966
rect 170082 79902 170134 79908
rect 170174 79960 170226 79966
rect 170174 79902 170226 79908
rect 170278 79778 170306 80036
rect 170370 79966 170398 80036
rect 170462 79971 170490 80036
rect 170358 79960 170410 79966
rect 170358 79902 170410 79908
rect 170448 79962 170504 79971
rect 170448 79897 170504 79906
rect 170554 79898 170582 80036
rect 170542 79892 170594 79898
rect 170542 79834 170594 79840
rect 170646 79778 170674 80036
rect 170738 79898 170766 80036
rect 170830 79937 170858 80036
rect 170922 79966 170950 80036
rect 170910 79960 170962 79966
rect 170816 79928 170872 79937
rect 170726 79892 170778 79898
rect 170910 79902 170962 79908
rect 170816 79863 170872 79872
rect 170726 79834 170778 79840
rect 171014 79830 171042 80036
rect 171002 79824 171054 79830
rect 169220 79716 169294 79744
rect 169772 79716 169846 79744
rect 170128 79756 170180 79762
rect 169116 79620 169168 79626
rect 169116 79562 169168 79568
rect 168852 79444 168972 79472
rect 168852 78674 168880 79444
rect 168930 79384 168986 79393
rect 168930 79319 168986 79328
rect 168840 78668 168892 78674
rect 168840 78610 168892 78616
rect 168668 78356 168788 78384
rect 168472 75268 168524 75274
rect 168472 75210 168524 75216
rect 168472 75064 168524 75070
rect 168472 75006 168524 75012
rect 168380 18692 168432 18698
rect 168380 18634 168432 18640
rect 168484 18630 168512 75006
rect 168668 70394 168696 78356
rect 168746 78296 168802 78305
rect 168746 78231 168802 78240
rect 168576 70366 168696 70394
rect 168576 21418 168604 70366
rect 168760 44878 168788 78231
rect 168840 75268 168892 75274
rect 168840 75210 168892 75216
rect 168852 49026 168880 75210
rect 168944 50386 168972 79319
rect 169024 77512 169076 77518
rect 169024 77454 169076 77460
rect 169036 77314 169064 77454
rect 169024 77308 169076 77314
rect 169024 77250 169076 77256
rect 169128 75070 169156 79562
rect 169116 75064 169168 75070
rect 169116 75006 169168 75012
rect 169220 70394 169248 79716
rect 169392 79688 169444 79694
rect 169392 79630 169444 79636
rect 169484 79688 169536 79694
rect 169484 79630 169536 79636
rect 169668 79688 169720 79694
rect 169668 79630 169720 79636
rect 169300 79620 169352 79626
rect 169300 79562 169352 79568
rect 169312 79014 169340 79562
rect 169300 79008 169352 79014
rect 169300 78950 169352 78956
rect 169404 75206 169432 79630
rect 169392 75200 169444 75206
rect 169392 75142 169444 75148
rect 169036 70366 169248 70394
rect 169036 64190 169064 70366
rect 169496 69698 169524 79630
rect 169576 79620 169628 79626
rect 169576 79562 169628 79568
rect 169588 79490 169616 79562
rect 169576 79484 169628 79490
rect 169576 79426 169628 79432
rect 169680 79370 169708 79630
rect 169588 79342 169708 79370
rect 169588 76537 169616 79342
rect 169668 79008 169720 79014
rect 169668 78950 169720 78956
rect 169574 76528 169630 76537
rect 169574 76463 169630 76472
rect 169484 69692 169536 69698
rect 169484 69634 169536 69640
rect 169024 64184 169076 64190
rect 169024 64126 169076 64132
rect 168932 50380 168984 50386
rect 168932 50322 168984 50328
rect 168840 49020 168892 49026
rect 168840 48962 168892 48968
rect 168748 44872 168800 44878
rect 168748 44814 168800 44820
rect 169680 43450 169708 78950
rect 169772 75070 169800 79716
rect 170278 79750 170536 79778
rect 170646 79750 170720 79778
rect 171106 79812 171134 80036
rect 171198 79937 171226 80036
rect 171184 79928 171240 79937
rect 171184 79863 171240 79872
rect 171106 79784 171180 79812
rect 171002 79766 171054 79772
rect 170128 79698 170180 79704
rect 170036 79688 170088 79694
rect 170036 79630 170088 79636
rect 169850 79384 169906 79393
rect 169850 79319 169906 79328
rect 169944 79348 169996 79354
rect 169760 75064 169812 75070
rect 169760 75006 169812 75012
rect 169760 74928 169812 74934
rect 169760 74870 169812 74876
rect 169668 43444 169720 43450
rect 169668 43386 169720 43392
rect 169772 31074 169800 74870
rect 169864 40730 169892 79319
rect 169944 79290 169996 79296
rect 169956 78810 169984 79290
rect 169944 78804 169996 78810
rect 169944 78746 169996 78752
rect 169944 75268 169996 75274
rect 169944 75210 169996 75216
rect 169956 42090 169984 75210
rect 170048 47598 170076 79630
rect 170140 58682 170168 79698
rect 170220 79688 170272 79694
rect 170220 79630 170272 79636
rect 170312 79688 170364 79694
rect 170312 79630 170364 79636
rect 170232 75274 170260 79630
rect 170324 77489 170352 79630
rect 170402 79520 170458 79529
rect 170402 79455 170458 79464
rect 170416 79218 170444 79455
rect 170508 79393 170536 79750
rect 170588 79688 170640 79694
rect 170588 79630 170640 79636
rect 170494 79384 170550 79393
rect 170494 79319 170550 79328
rect 170404 79212 170456 79218
rect 170404 79154 170456 79160
rect 170600 78713 170628 79630
rect 170586 78704 170642 78713
rect 170586 78639 170642 78648
rect 170494 78296 170550 78305
rect 170494 78231 170550 78240
rect 170310 77480 170366 77489
rect 170310 77415 170366 77424
rect 170220 75268 170272 75274
rect 170220 75210 170272 75216
rect 170220 75064 170272 75070
rect 170220 75006 170272 75012
rect 170232 65550 170260 75006
rect 170508 74934 170536 78231
rect 170586 78160 170642 78169
rect 170586 78095 170642 78104
rect 170496 74928 170548 74934
rect 170496 74870 170548 74876
rect 170600 68338 170628 78095
rect 170692 78062 170720 79750
rect 171048 79688 171100 79694
rect 171048 79630 171100 79636
rect 170772 79552 170824 79558
rect 170772 79494 170824 79500
rect 170784 79354 170812 79494
rect 170864 79484 170916 79490
rect 170864 79426 170916 79432
rect 170772 79348 170824 79354
rect 170772 79290 170824 79296
rect 170772 78668 170824 78674
rect 170772 78610 170824 78616
rect 170680 78056 170732 78062
rect 170680 77998 170732 78004
rect 170784 69766 170812 78610
rect 170876 77294 170904 79426
rect 170876 77266 170996 77294
rect 170968 75993 170996 77266
rect 170954 75984 171010 75993
rect 170954 75919 171010 75928
rect 171060 75834 171088 79630
rect 171152 79490 171180 79784
rect 171290 79744 171318 80036
rect 171382 79898 171410 80036
rect 171474 79971 171502 80036
rect 171460 79962 171516 79971
rect 171566 79966 171594 80036
rect 171370 79892 171422 79898
rect 171460 79897 171516 79906
rect 171554 79960 171606 79966
rect 171554 79902 171606 79908
rect 171370 79834 171422 79840
rect 171658 79812 171686 80036
rect 171750 79937 171778 80036
rect 171736 79928 171792 79937
rect 171736 79863 171792 79872
rect 171520 79784 171686 79812
rect 171290 79716 171364 79744
rect 171232 79620 171284 79626
rect 171232 79562 171284 79568
rect 171140 79484 171192 79490
rect 171140 79426 171192 79432
rect 171244 79286 171272 79562
rect 171232 79280 171284 79286
rect 171232 79222 171284 79228
rect 171336 78713 171364 79716
rect 171416 79688 171468 79694
rect 171416 79630 171468 79636
rect 171520 79642 171548 79784
rect 171842 79778 171870 80036
rect 171934 79937 171962 80036
rect 171920 79928 171976 79937
rect 171920 79863 171976 79872
rect 172026 79812 172054 80036
rect 172118 79830 172146 80036
rect 172210 79937 172238 80036
rect 172196 79928 172252 79937
rect 172196 79863 172252 79872
rect 171980 79784 172054 79812
rect 172106 79824 172158 79830
rect 171842 79750 171916 79778
rect 171692 79688 171744 79694
rect 171322 78704 171378 78713
rect 171322 78639 171378 78648
rect 171230 78024 171286 78033
rect 171230 77959 171286 77968
rect 171244 76566 171272 77959
rect 171428 77926 171456 79630
rect 171520 79614 171594 79642
rect 171692 79630 171744 79636
rect 171566 79540 171594 79614
rect 171566 79512 171640 79540
rect 171612 78606 171640 79512
rect 171600 78600 171652 78606
rect 171600 78542 171652 78548
rect 171416 77920 171468 77926
rect 171416 77862 171468 77868
rect 171704 77738 171732 79630
rect 171784 79416 171836 79422
rect 171782 79384 171784 79393
rect 171836 79384 171838 79393
rect 171782 79319 171838 79328
rect 171888 78674 171916 79750
rect 171876 78668 171928 78674
rect 171876 78610 171928 78616
rect 171784 78532 171836 78538
rect 171784 78474 171836 78480
rect 171416 77716 171468 77722
rect 171416 77658 171468 77664
rect 171520 77710 171732 77738
rect 171232 76560 171284 76566
rect 171232 76502 171284 76508
rect 171060 75806 171180 75834
rect 171152 73166 171180 75806
rect 171140 73160 171192 73166
rect 171140 73102 171192 73108
rect 170772 69760 170824 69766
rect 170772 69702 170824 69708
rect 171140 68876 171192 68882
rect 171140 68818 171192 68824
rect 170588 68332 170640 68338
rect 170588 68274 170640 68280
rect 170220 65544 170272 65550
rect 170220 65486 170272 65492
rect 170128 58676 170180 58682
rect 170128 58618 170180 58624
rect 170036 47592 170088 47598
rect 170036 47534 170088 47540
rect 169944 42084 169996 42090
rect 169944 42026 169996 42032
rect 169852 40724 169904 40730
rect 169852 40666 169904 40672
rect 169760 31068 169812 31074
rect 169760 31010 169812 31016
rect 168656 21616 168708 21622
rect 168656 21558 168708 21564
rect 168564 21412 168616 21418
rect 168564 21354 168616 21360
rect 168472 18624 168524 18630
rect 168472 18566 168524 18572
rect 168668 16574 168696 21558
rect 168668 16546 169616 16574
rect 168288 4820 168340 4826
rect 168288 4762 168340 4768
rect 168380 3732 168432 3738
rect 168380 3674 168432 3680
rect 168392 480 168420 3674
rect 169588 480 169616 16546
rect 171152 6914 171180 68818
rect 171428 9382 171456 77658
rect 171520 75750 171548 77710
rect 171692 77648 171744 77654
rect 171692 77590 171744 77596
rect 171704 77466 171732 77590
rect 171796 77518 171824 78474
rect 171980 78305 172008 79784
rect 172106 79766 172158 79772
rect 172302 79676 172330 80036
rect 172394 79744 172422 80036
rect 172486 79937 172514 80036
rect 172472 79928 172528 79937
rect 172472 79863 172528 79872
rect 172578 79744 172606 80036
rect 172670 79812 172698 80036
rect 172762 79966 172790 80036
rect 172854 79966 172882 80036
rect 172750 79960 172802 79966
rect 172750 79902 172802 79908
rect 172842 79960 172894 79966
rect 172842 79902 172894 79908
rect 172946 79898 172974 80036
rect 173038 79898 173066 80036
rect 172934 79892 172986 79898
rect 172934 79834 172986 79840
rect 173026 79892 173078 79898
rect 173026 79834 173078 79840
rect 172670 79784 172744 79812
rect 172394 79716 172468 79744
rect 172302 79648 172376 79676
rect 172060 79620 172112 79626
rect 172060 79562 172112 79568
rect 172072 78538 172100 79562
rect 172060 78532 172112 78538
rect 172060 78474 172112 78480
rect 171966 78296 172022 78305
rect 171966 78231 172022 78240
rect 172058 77888 172114 77897
rect 171968 77852 172020 77858
rect 172058 77823 172114 77832
rect 171968 77794 172020 77800
rect 171876 77784 171928 77790
rect 171876 77726 171928 77732
rect 171612 77438 171732 77466
rect 171784 77512 171836 77518
rect 171784 77454 171836 77460
rect 171508 75744 171560 75750
rect 171508 75686 171560 75692
rect 171612 70394 171640 77438
rect 171692 77308 171744 77314
rect 171692 77250 171744 77256
rect 171520 70366 171640 70394
rect 171520 43518 171548 70366
rect 171704 49162 171732 77250
rect 171888 76480 171916 77726
rect 171796 76452 171916 76480
rect 171692 49156 171744 49162
rect 171692 49098 171744 49104
rect 171508 43512 171560 43518
rect 171508 43454 171560 43460
rect 171796 16574 171824 76452
rect 171980 70394 172008 77794
rect 171888 70366 172008 70394
rect 171888 44946 171916 70366
rect 171876 44940 171928 44946
rect 171876 44882 171928 44888
rect 172072 21486 172100 77823
rect 172244 77580 172296 77586
rect 172244 77522 172296 77528
rect 172152 77376 172204 77382
rect 172152 77318 172204 77324
rect 172164 28286 172192 77318
rect 172152 28280 172204 28286
rect 172152 28222 172204 28228
rect 172060 21480 172112 21486
rect 172060 21422 172112 21428
rect 171796 16546 172100 16574
rect 171416 9376 171468 9382
rect 171416 9318 171468 9324
rect 171152 6886 171732 6914
rect 171704 3482 171732 6886
rect 170772 3460 170824 3466
rect 171704 3454 172008 3482
rect 170772 3402 170824 3408
rect 170784 480 170812 3402
rect 171980 480 172008 3454
rect 172072 3194 172100 16546
rect 172256 3262 172284 77522
rect 172348 77217 172376 79648
rect 172440 79393 172468 79716
rect 172532 79716 172606 79744
rect 172426 79384 172482 79393
rect 172426 79319 172482 79328
rect 172428 79076 172480 79082
rect 172428 79018 172480 79024
rect 172334 77208 172390 77217
rect 172334 77143 172390 77152
rect 172440 64874 172468 79018
rect 172532 79014 172560 79716
rect 172612 79620 172664 79626
rect 172612 79562 172664 79568
rect 172520 79008 172572 79014
rect 172520 78950 172572 78956
rect 172624 75818 172652 79562
rect 172716 79082 172744 79784
rect 172980 79756 173032 79762
rect 173130 79744 173158 80036
rect 173222 79937 173250 80036
rect 173314 79966 173342 80036
rect 173406 79966 173434 80036
rect 173302 79960 173354 79966
rect 173208 79928 173264 79937
rect 173302 79902 173354 79908
rect 173394 79960 173446 79966
rect 173394 79902 173446 79908
rect 173498 79898 173526 80036
rect 173590 79966 173618 80036
rect 173578 79960 173630 79966
rect 173578 79902 173630 79908
rect 173208 79863 173264 79872
rect 173486 79892 173538 79898
rect 173486 79834 173538 79840
rect 173302 79756 173354 79762
rect 173130 79716 173204 79744
rect 172980 79698 173032 79704
rect 172888 79620 172940 79626
rect 172808 79580 172888 79608
rect 172704 79076 172756 79082
rect 172704 79018 172756 79024
rect 172808 78946 172836 79580
rect 172888 79562 172940 79568
rect 172886 79248 172942 79257
rect 172886 79183 172942 79192
rect 172900 78946 172928 79183
rect 172796 78940 172848 78946
rect 172796 78882 172848 78888
rect 172888 78940 172940 78946
rect 172888 78882 172940 78888
rect 172794 77752 172850 77761
rect 172794 77687 172850 77696
rect 172808 77586 172836 77687
rect 172796 77580 172848 77586
rect 172796 77522 172848 77528
rect 172992 75914 173020 79698
rect 173070 79656 173126 79665
rect 173070 79591 173126 79600
rect 173084 79393 173112 79591
rect 173176 79472 173204 79716
rect 173682 79744 173710 80036
rect 173774 79971 173802 80036
rect 173760 79962 173816 79971
rect 173760 79897 173816 79906
rect 173866 79830 173894 80036
rect 173958 79971 173986 80036
rect 173944 79962 174000 79971
rect 173944 79897 174000 79906
rect 173854 79824 173906 79830
rect 173854 79766 173906 79772
rect 173354 79716 173572 79744
rect 173302 79698 173354 79704
rect 173348 79620 173400 79626
rect 173348 79562 173400 79568
rect 173440 79620 173492 79626
rect 173440 79562 173492 79568
rect 173176 79444 173296 79472
rect 173070 79384 173126 79393
rect 173070 79319 173126 79328
rect 173268 78849 173296 79444
rect 173360 79393 173388 79562
rect 173346 79384 173402 79393
rect 173346 79319 173402 79328
rect 173346 79248 173402 79257
rect 173346 79183 173402 79192
rect 173254 78840 173310 78849
rect 173360 78810 173388 79183
rect 173452 79121 173480 79562
rect 173438 79112 173494 79121
rect 173438 79047 173494 79056
rect 173544 78985 173572 79716
rect 173636 79716 173710 79744
rect 173762 79756 173814 79762
rect 173636 79558 173664 79716
rect 173762 79698 173814 79704
rect 173774 79642 173802 79698
rect 173774 79614 173894 79642
rect 173866 79608 173894 79614
rect 174050 79608 174078 80036
rect 174142 79966 174170 80036
rect 174130 79960 174182 79966
rect 174130 79902 174182 79908
rect 174234 79914 174262 80036
rect 174340 80022 174584 80050
rect 174360 79960 174412 79966
rect 174234 79886 174308 79914
rect 174360 79902 174412 79908
rect 173866 79580 173940 79608
rect 173624 79552 173676 79558
rect 173624 79494 173676 79500
rect 173530 78976 173586 78985
rect 173912 78946 173940 79580
rect 174004 79580 174078 79608
rect 174004 79218 174032 79580
rect 174280 79370 174308 79886
rect 174188 79342 174308 79370
rect 174372 79354 174400 79902
rect 174452 79824 174504 79830
rect 174452 79766 174504 79772
rect 174360 79348 174412 79354
rect 174084 79280 174136 79286
rect 174084 79222 174136 79228
rect 173992 79212 174044 79218
rect 173992 79154 174044 79160
rect 174096 78946 174124 79222
rect 173530 78911 173586 78920
rect 173900 78940 173952 78946
rect 173900 78882 173952 78888
rect 174084 78940 174136 78946
rect 174084 78882 174136 78888
rect 173254 78775 173310 78784
rect 173348 78804 173400 78810
rect 173348 78746 173400 78752
rect 173162 76392 173218 76401
rect 173162 76327 173218 76336
rect 173256 76356 173308 76362
rect 172992 75886 173112 75914
rect 173072 75880 173124 75886
rect 173072 75822 173124 75828
rect 172612 75812 172664 75818
rect 172612 75754 172664 75760
rect 172348 64846 172468 64874
rect 172348 6662 172376 64846
rect 172336 6656 172388 6662
rect 172336 6598 172388 6604
rect 173176 5250 173204 76327
rect 173256 76298 173308 76304
rect 173268 5386 173296 76298
rect 173346 75712 173402 75721
rect 173346 75647 173402 75656
rect 173360 6914 173388 75647
rect 173440 74180 173492 74186
rect 173440 74122 173492 74128
rect 173452 11778 173480 74122
rect 173900 74112 173952 74118
rect 173900 74054 173952 74060
rect 173532 72956 173584 72962
rect 173532 72898 173584 72904
rect 173544 11914 173572 72898
rect 173544 11886 173756 11914
rect 173452 11750 173664 11778
rect 173532 11688 173584 11694
rect 173532 11630 173584 11636
rect 173360 6886 173480 6914
rect 173268 5358 173388 5386
rect 173176 5222 173296 5250
rect 173268 3670 173296 5222
rect 173164 3664 173216 3670
rect 173164 3606 173216 3612
rect 173256 3664 173308 3670
rect 173256 3606 173308 3612
rect 172244 3256 172296 3262
rect 172244 3198 172296 3204
rect 172060 3188 172112 3194
rect 172060 3130 172112 3136
rect 173176 480 173204 3606
rect 173360 3602 173388 5358
rect 173348 3596 173400 3602
rect 173348 3538 173400 3544
rect 173452 3466 173480 6886
rect 173544 3738 173572 11630
rect 173532 3732 173584 3738
rect 173532 3674 173584 3680
rect 173440 3460 173492 3466
rect 173440 3402 173492 3408
rect 173636 3369 173664 11750
rect 173728 11694 173756 11886
rect 173716 11688 173768 11694
rect 173716 11630 173768 11636
rect 173622 3360 173678 3369
rect 173622 3295 173678 3304
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 173912 354 173940 74054
rect 174188 70394 174216 79342
rect 174360 79290 174412 79296
rect 174268 79280 174320 79286
rect 174268 79222 174320 79228
rect 174280 78742 174308 79222
rect 174268 78736 174320 78742
rect 174268 78678 174320 78684
rect 174464 77994 174492 79766
rect 174452 77988 174504 77994
rect 174452 77930 174504 77936
rect 174450 71088 174506 71097
rect 174450 71023 174506 71032
rect 174004 70366 174216 70394
rect 174004 45558 174032 70366
rect 174464 64874 174492 71023
rect 174556 70106 174584 80022
rect 174648 79966 174676 80378
rect 174740 80238 174768 80514
rect 174924 80306 174952 80543
rect 174912 80300 174964 80306
rect 174912 80242 174964 80248
rect 174728 80232 174780 80238
rect 174728 80174 174780 80180
rect 177396 80096 177448 80102
rect 177396 80038 177448 80044
rect 174636 79960 174688 79966
rect 174636 79902 174688 79908
rect 177408 79354 177436 80038
rect 177396 79348 177448 79354
rect 177396 79290 177448 79296
rect 178052 78674 178080 80582
rect 178040 78668 178092 78674
rect 178040 78610 178092 78616
rect 178972 78538 179000 82078
rect 179420 80844 179472 80850
rect 179420 80786 179472 80792
rect 179432 78577 179460 80786
rect 179418 78568 179474 78577
rect 178960 78532 179012 78538
rect 179418 78503 179474 78512
rect 178960 78474 179012 78480
rect 178040 77512 178092 77518
rect 178040 77454 178092 77460
rect 176658 75576 176714 75585
rect 176658 75511 176714 75520
rect 174544 70100 174596 70106
rect 174544 70042 174596 70048
rect 174464 64846 174584 64874
rect 173992 45552 174044 45558
rect 173992 45494 174044 45500
rect 174556 3534 174584 64846
rect 176672 3602 176700 75511
rect 176752 71392 176804 71398
rect 176752 71334 176804 71340
rect 176660 3596 176712 3602
rect 176660 3538 176712 3544
rect 174544 3528 174596 3534
rect 174544 3470 174596 3476
rect 175464 3528 175516 3534
rect 176764 3482 176792 71334
rect 178052 16574 178080 77454
rect 178684 75268 178736 75274
rect 178684 75210 178736 75216
rect 178696 75138 178724 75210
rect 178684 75132 178736 75138
rect 178684 75074 178736 75080
rect 179512 60308 179564 60314
rect 179512 60250 179564 60256
rect 179524 16574 179552 60250
rect 179708 22778 179736 130455
rect 180064 125656 180116 125662
rect 180064 125598 180116 125604
rect 180076 80481 180104 125598
rect 180168 114578 180196 139334
rect 180812 114753 180840 231134
rect 192484 218068 192536 218074
rect 192484 218010 192536 218016
rect 180892 209092 180944 209098
rect 180892 209034 180944 209040
rect 180904 122913 180932 209034
rect 189724 178084 189776 178090
rect 189724 178026 189776 178032
rect 182272 169040 182324 169046
rect 182272 168982 182324 168988
rect 180984 159384 181036 159390
rect 180984 159326 181036 159332
rect 180890 122904 180946 122913
rect 180890 122839 180946 122848
rect 180798 114744 180854 114753
rect 180798 114679 180854 114688
rect 180156 114572 180208 114578
rect 180156 114514 180208 114520
rect 180996 112033 181024 159326
rect 181444 151836 181496 151842
rect 181444 151778 181496 151784
rect 181076 139460 181128 139466
rect 181076 139402 181128 139408
rect 181088 128353 181116 139402
rect 181074 128344 181130 128353
rect 181074 128279 181130 128288
rect 180982 112024 181038 112033
rect 180982 111959 181038 111968
rect 180156 111852 180208 111858
rect 180156 111794 180208 111800
rect 180062 80472 180118 80481
rect 180062 80407 180118 80416
rect 180168 79694 180196 111794
rect 180156 79688 180208 79694
rect 180156 79630 180208 79636
rect 181456 79422 181484 151778
rect 181536 140140 181588 140146
rect 181536 140082 181588 140088
rect 181548 119882 181576 140082
rect 182180 139324 182232 139330
rect 182180 139266 182232 139272
rect 182192 126993 182220 139266
rect 182178 126984 182234 126993
rect 182178 126919 182234 126928
rect 182284 124273 182312 168982
rect 182364 164892 182416 164898
rect 182364 164834 182416 164840
rect 182270 124264 182326 124273
rect 182270 124199 182326 124208
rect 182376 121553 182404 164834
rect 182732 162172 182784 162178
rect 182732 162114 182784 162120
rect 182456 141568 182508 141574
rect 182456 141510 182508 141516
rect 182362 121544 182418 121553
rect 182362 121479 182418 121488
rect 181536 119876 181588 119882
rect 181536 119818 181588 119824
rect 182272 119876 182324 119882
rect 182272 119818 182324 119824
rect 182180 114504 182232 114510
rect 182180 114446 182232 114452
rect 182192 109313 182220 114446
rect 182178 109304 182234 109313
rect 182178 109239 182234 109248
rect 182284 107953 182312 119818
rect 182468 110673 182496 141510
rect 182548 141500 182600 141506
rect 182548 141442 182600 141448
rect 182560 118833 182588 141442
rect 182640 140072 182692 140078
rect 182640 140014 182692 140020
rect 182546 118824 182602 118833
rect 182546 118759 182602 118768
rect 182652 117473 182680 140014
rect 182744 120193 182772 162114
rect 188344 138032 188396 138038
rect 188344 137974 188396 137980
rect 183006 129704 183062 129713
rect 183006 129639 183062 129648
rect 182730 120184 182786 120193
rect 182730 120119 182786 120128
rect 182638 117464 182694 117473
rect 182638 117399 182694 117408
rect 182454 110664 182510 110673
rect 182454 110599 182510 110608
rect 182270 107944 182326 107953
rect 182270 107879 182326 107888
rect 182824 99408 182876 99414
rect 182824 99350 182876 99356
rect 182548 86556 182600 86562
rect 182548 86498 182600 86504
rect 182560 86193 182588 86498
rect 182546 86184 182602 86193
rect 182546 86119 182602 86128
rect 182732 84924 182784 84930
rect 182732 84866 182784 84872
rect 182744 84833 182772 84866
rect 182730 84824 182786 84833
rect 182730 84759 182786 84768
rect 182836 83473 182864 99350
rect 182822 83464 182878 83473
rect 182822 83399 182878 83408
rect 182822 82104 182878 82113
rect 182822 82039 182878 82048
rect 182178 80744 182234 80753
rect 182178 80679 182234 80688
rect 182192 80102 182220 80679
rect 182180 80096 182232 80102
rect 182180 80038 182232 80044
rect 181444 79416 181496 79422
rect 181444 79358 181496 79364
rect 181444 72888 181496 72894
rect 181444 72830 181496 72836
rect 180800 59016 180852 59022
rect 180800 58958 180852 58964
rect 179696 22772 179748 22778
rect 179696 22714 179748 22720
rect 180812 16574 180840 58958
rect 178052 16546 178632 16574
rect 179524 16546 180288 16574
rect 180812 16546 181024 16574
rect 178132 3732 178184 3738
rect 178132 3674 178184 3680
rect 177856 3596 177908 3602
rect 177856 3538 177908 3544
rect 175464 3470 175516 3476
rect 175476 480 175504 3470
rect 176672 3454 176792 3482
rect 176672 480 176700 3454
rect 177868 480 177896 3538
rect 178144 3466 178172 3674
rect 178132 3460 178184 3466
rect 178132 3402 178184 3408
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181456 3262 181484 72830
rect 182836 60722 182864 82039
rect 183020 68678 183048 129639
rect 183284 107636 183336 107642
rect 183284 107578 183336 107584
rect 183296 106593 183324 107578
rect 183282 106584 183338 106593
rect 183282 106519 183338 106528
rect 183284 106276 183336 106282
rect 183284 106218 183336 106224
rect 183296 105233 183324 106218
rect 183282 105224 183338 105233
rect 183282 105159 183338 105168
rect 183284 104848 183336 104854
rect 183284 104790 183336 104796
rect 183296 103873 183324 104790
rect 183282 103864 183338 103873
rect 183282 103799 183338 103808
rect 183284 103488 183336 103494
rect 183284 103430 183336 103436
rect 183296 102513 183324 103430
rect 183282 102504 183338 102513
rect 183282 102439 183338 102448
rect 183284 102128 183336 102134
rect 183284 102070 183336 102076
rect 183296 101153 183324 102070
rect 183282 101144 183338 101153
rect 183282 101079 183338 101088
rect 183192 100700 183244 100706
rect 183192 100642 183244 100648
rect 183204 99793 183232 100642
rect 183190 99784 183246 99793
rect 183190 99719 183246 99728
rect 183192 99340 183244 99346
rect 183192 99282 183244 99288
rect 183204 98433 183232 99282
rect 183190 98424 183246 98433
rect 183190 98359 183246 98368
rect 183192 97980 183244 97986
rect 183192 97922 183244 97928
rect 183204 97073 183232 97922
rect 183190 97064 183246 97073
rect 183190 96999 183246 97008
rect 183192 96620 183244 96626
rect 183192 96562 183244 96568
rect 183204 95713 183232 96562
rect 183190 95704 183246 95713
rect 183190 95639 183246 95648
rect 183468 95192 183520 95198
rect 183468 95134 183520 95140
rect 183480 94353 183508 95134
rect 183466 94344 183522 94353
rect 183466 94279 183522 94288
rect 183468 93832 183520 93838
rect 183468 93774 183520 93780
rect 183480 92993 183508 93774
rect 183466 92984 183522 92993
rect 183466 92919 183522 92928
rect 183468 92472 183520 92478
rect 183468 92414 183520 92420
rect 183480 91633 183508 92414
rect 183466 91624 183522 91633
rect 183466 91559 183522 91568
rect 183468 91044 183520 91050
rect 183468 90986 183520 90992
rect 183480 90273 183508 90986
rect 183466 90264 183522 90273
rect 183466 90199 183522 90208
rect 183468 89684 183520 89690
rect 183468 89626 183520 89632
rect 183480 88913 183508 89626
rect 183466 88904 183522 88913
rect 183466 88839 183522 88848
rect 183468 88324 183520 88330
rect 183468 88266 183520 88272
rect 183480 87553 183508 88266
rect 183466 87544 183522 87553
rect 183466 87479 183522 87488
rect 188356 84930 188384 137974
rect 189736 86562 189764 178026
rect 192496 88330 192524 218010
rect 207032 198082 207060 230588
rect 236012 230574 236578 230602
rect 266372 230574 266570 230602
rect 236012 202162 236040 230574
rect 266372 203590 266400 230574
rect 296732 228478 296760 230588
rect 296720 228472 296772 228478
rect 296720 228414 296772 228420
rect 266360 203584 266412 203590
rect 266360 203526 266412 203532
rect 236000 202156 236052 202162
rect 236000 202098 236052 202104
rect 207020 198076 207072 198082
rect 207020 198018 207072 198024
rect 327092 196654 327120 230588
rect 356072 230574 356546 230602
rect 356072 198014 356100 230574
rect 383660 221876 383712 221882
rect 383660 221818 383712 221824
rect 383672 218142 383700 221818
rect 382280 218136 382332 218142
rect 382280 218078 382332 218084
rect 383660 218136 383712 218142
rect 383660 218078 383712 218084
rect 382292 209846 382320 218078
rect 382280 209840 382332 209846
rect 382280 209782 382332 209788
rect 378784 209772 378836 209778
rect 378784 209714 378836 209720
rect 356060 198008 356112 198014
rect 356060 197950 356112 197956
rect 378796 197402 378824 209714
rect 384304 205760 384356 205766
rect 384304 205702 384356 205708
rect 376024 197396 376076 197402
rect 376024 197338 376076 197344
rect 378784 197396 378836 197402
rect 378784 197338 378836 197344
rect 327080 196648 327132 196654
rect 327080 196590 327132 196596
rect 371884 191140 371936 191146
rect 371884 191082 371936 191088
rect 371896 175982 371924 191082
rect 355324 175976 355376 175982
rect 355324 175918 355376 175924
rect 371884 175976 371936 175982
rect 371884 175918 371936 175924
rect 355336 163538 355364 175918
rect 345664 163532 345716 163538
rect 345664 163474 345716 163480
rect 355324 163532 355376 163538
rect 355324 163474 355376 163480
rect 345676 149802 345704 163474
rect 376036 160138 376064 197338
rect 379520 193792 379572 193798
rect 379520 193734 379572 193740
rect 379532 191146 379560 193734
rect 379520 191140 379572 191146
rect 379520 191082 379572 191088
rect 376024 160132 376076 160138
rect 376024 160074 376076 160080
rect 373264 160064 373316 160070
rect 373264 160006 373316 160012
rect 319444 149796 319496 149802
rect 319444 149738 319496 149744
rect 345664 149796 345716 149802
rect 345664 149738 345716 149744
rect 319456 139466 319484 149738
rect 316684 139460 316736 139466
rect 316684 139402 316736 139408
rect 319444 139460 319496 139466
rect 319444 139402 319496 139408
rect 304264 123480 304316 123486
rect 304264 123422 304316 123428
rect 304276 107642 304304 123422
rect 304264 107636 304316 107642
rect 304264 107578 304316 107584
rect 316696 89010 316724 139402
rect 373276 131170 373304 160006
rect 384316 151910 384344 205702
rect 384408 193798 384436 231134
rect 386524 228410 386552 230588
rect 390560 230512 390612 230518
rect 390560 230454 390612 230460
rect 390572 229094 390600 230454
rect 390480 229066 390600 229094
rect 386512 228404 386564 228410
rect 386512 228346 386564 228352
rect 390480 225078 390508 229066
rect 391940 228404 391992 228410
rect 391940 228346 391992 228352
rect 387800 225072 387852 225078
rect 387800 225014 387852 225020
rect 390468 225072 390520 225078
rect 390468 225014 390520 225020
rect 387064 225004 387116 225010
rect 387064 224946 387116 224952
rect 387076 205766 387104 224946
rect 387812 221882 387840 225014
rect 391952 225010 391980 228346
rect 391940 225004 391992 225010
rect 391940 224946 391992 224952
rect 387800 221876 387852 221882
rect 387800 221818 387852 221824
rect 387064 205760 387116 205766
rect 387064 205702 387116 205708
rect 384396 193792 384448 193798
rect 384396 193734 384448 193740
rect 381544 151904 381596 151910
rect 381544 151846 381596 151852
rect 384304 151904 384356 151910
rect 384304 151846 384356 151852
rect 381556 144294 381584 151846
rect 373356 144288 373408 144294
rect 373356 144230 373408 144236
rect 381544 144288 381596 144294
rect 381544 144230 381596 144236
rect 369860 131164 369912 131170
rect 369860 131106 369912 131112
rect 373264 131164 373316 131170
rect 373264 131106 373316 131112
rect 369872 129062 369900 131106
rect 355968 129056 356020 129062
rect 355968 128998 356020 129004
rect 369860 129056 369912 129062
rect 369860 128998 369912 129004
rect 355980 127634 356008 128998
rect 328920 127628 328972 127634
rect 328920 127570 328972 127576
rect 355968 127628 356020 127634
rect 355968 127570 356020 127576
rect 328932 126070 328960 127570
rect 326712 126064 326764 126070
rect 326712 126006 326764 126012
rect 328920 126064 328972 126070
rect 328920 126006 328972 126012
rect 326724 124506 326752 126006
rect 322940 124500 322992 124506
rect 322940 124442 322992 124448
rect 326712 124500 326764 124506
rect 326712 124442 326764 124448
rect 322952 123486 322980 124442
rect 373368 123690 373396 144230
rect 367744 123684 367796 123690
rect 367744 123626 367796 123632
rect 373356 123684 373408 123690
rect 373356 123626 373408 123632
rect 322940 123480 322992 123486
rect 322940 123422 322992 123428
rect 305644 89004 305696 89010
rect 305644 88946 305696 88952
rect 316684 89004 316736 89010
rect 316684 88946 316736 88952
rect 192484 88324 192536 88330
rect 192484 88266 192536 88272
rect 189724 86556 189776 86562
rect 189724 86498 189776 86504
rect 188344 84924 188396 84930
rect 188344 84866 188396 84872
rect 305656 83502 305684 88946
rect 293960 83496 294012 83502
rect 293960 83438 294012 83444
rect 305644 83496 305696 83502
rect 305644 83438 305696 83444
rect 252560 80300 252612 80306
rect 252560 80242 252612 80248
rect 184204 80096 184256 80102
rect 184204 80038 184256 80044
rect 183008 68672 183060 68678
rect 183008 68614 183060 68620
rect 182824 60716 182876 60722
rect 182824 60658 182876 60664
rect 183560 60240 183612 60246
rect 183560 60182 183612 60188
rect 183572 16574 183600 60182
rect 184216 22778 184244 80038
rect 184940 79416 184992 79422
rect 184940 79358 184992 79364
rect 184952 78305 184980 79358
rect 195980 78464 196032 78470
rect 195980 78406 196032 78412
rect 184938 78296 184994 78305
rect 184938 78231 184994 78240
rect 194598 74352 194654 74361
rect 194598 74287 194654 74296
rect 184940 70236 184992 70242
rect 184940 70178 184992 70184
rect 184204 22772 184256 22778
rect 184204 22714 184256 22720
rect 183572 16546 183784 16574
rect 181444 3256 181496 3262
rect 181444 3198 181496 3204
rect 182548 3188 182600 3194
rect 182548 3130 182600 3136
rect 182560 480 182588 3130
rect 183756 480 183784 16546
rect 184952 3738 184980 70178
rect 189080 67176 189132 67182
rect 189080 67118 189132 67124
rect 185032 53304 185084 53310
rect 185032 53246 185084 53252
rect 184940 3732 184992 3738
rect 184940 3674 184992 3680
rect 185044 3482 185072 53246
rect 187700 42220 187752 42226
rect 187700 42162 187752 42168
rect 186320 23044 186372 23050
rect 186320 22986 186372 22992
rect 186332 16574 186360 22986
rect 187712 16574 187740 42162
rect 189092 16574 189120 67118
rect 193218 65512 193274 65521
rect 193218 65447 193274 65456
rect 190460 62960 190512 62966
rect 190460 62902 190512 62908
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 189092 16546 189304 16574
rect 186136 3732 186188 3738
rect 186136 3674 186188 3680
rect 186228 3732 186280 3738
rect 186228 3674 186280 3680
rect 184952 3454 185072 3482
rect 184952 480 184980 3454
rect 186148 480 186176 3674
rect 186240 3262 186268 3674
rect 186228 3256 186280 3262
rect 186228 3198 186280 3204
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 181414 -960 181526 326
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 62902
rect 191838 40896 191894 40905
rect 191838 40831 191894 40840
rect 191852 16574 191880 40831
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 480 193260 65447
rect 193310 24440 193366 24449
rect 193310 24375 193366 24384
rect 193324 16574 193352 24375
rect 194612 16574 194640 74287
rect 195992 16574 196020 78406
rect 197360 77240 197412 77246
rect 197360 77182 197412 77188
rect 197372 16574 197400 77182
rect 213920 77172 213972 77178
rect 213920 77114 213972 77120
rect 211158 77072 211214 77081
rect 211158 77007 211214 77016
rect 209780 74044 209832 74050
rect 209780 73986 209832 73992
rect 202880 68808 202932 68814
rect 202880 68750 202932 68756
rect 201500 57316 201552 57322
rect 201500 57258 201552 57264
rect 198740 18828 198792 18834
rect 198740 18770 198792 18776
rect 193324 16546 194456 16574
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 194428 480 194456 16546
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 18770
rect 200304 3324 200356 3330
rect 200304 3266 200356 3272
rect 200316 480 200344 3266
rect 201512 480 201540 57258
rect 202892 16574 202920 68750
rect 207020 67108 207072 67114
rect 207020 67050 207072 67056
rect 204260 51876 204312 51882
rect 204260 51818 204312 51824
rect 204272 16574 204300 51818
rect 205640 31408 205692 31414
rect 205640 31350 205692 31356
rect 205652 16574 205680 31350
rect 202892 16546 203472 16574
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 202696 12368 202748 12374
rect 202696 12310 202748 12316
rect 202708 480 202736 12310
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 67050
rect 208400 46436 208452 46442
rect 208400 46378 208452 46384
rect 208412 16574 208440 46378
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 480 209820 73986
rect 209872 70168 209924 70174
rect 209872 70110 209924 70116
rect 209884 16574 209912 70110
rect 211172 16574 211200 77007
rect 212538 17368 212594 17377
rect 212538 17303 212594 17312
rect 212552 16574 212580 17303
rect 213932 16574 213960 77114
rect 226340 77104 226392 77110
rect 226340 77046 226392 77052
rect 223580 73976 223632 73982
rect 223580 73918 223632 73924
rect 219440 54732 219492 54738
rect 219440 54674 219492 54680
rect 215300 47864 215352 47870
rect 215300 47806 215352 47812
rect 209884 16546 211016 16574
rect 211172 16546 211752 16574
rect 212552 16546 213408 16574
rect 213932 16546 214512 16574
rect 210988 480 211016 16546
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213380 480 213408 16546
rect 214484 480 214512 16546
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 47806
rect 218152 45076 218204 45082
rect 218152 45018 218204 45024
rect 216680 31340 216732 31346
rect 216680 31282 216732 31288
rect 216692 16574 216720 31282
rect 218164 16574 218192 45018
rect 219452 16574 219480 54674
rect 222200 24268 222252 24274
rect 222200 24210 222252 24216
rect 222212 16574 222240 24210
rect 216692 16546 216904 16574
rect 218164 16546 219296 16574
rect 219452 16546 220032 16574
rect 222212 16546 222792 16574
rect 216876 480 216904 16546
rect 218060 3392 218112 3398
rect 218060 3334 218112 3340
rect 218072 480 218100 3334
rect 219268 480 219296 16546
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 221556 4140 221608 4146
rect 221556 4082 221608 4088
rect 221568 480 221596 4082
rect 222764 480 222792 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 220422 -960 220534 326
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223592 354 223620 73918
rect 225142 3632 225198 3641
rect 225142 3567 225198 3576
rect 225156 480 225184 3567
rect 226352 480 226380 77046
rect 231860 77036 231912 77042
rect 231860 76978 231912 76984
rect 230478 74216 230534 74225
rect 230478 74151 230534 74160
rect 227718 58576 227774 58585
rect 227718 58511 227774 58520
rect 227732 16574 227760 58511
rect 230492 16574 230520 74151
rect 227732 16546 228312 16574
rect 230492 16546 231072 16574
rect 227534 7848 227590 7857
rect 227534 7783 227590 7792
rect 227548 480 227576 7783
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 229374 13696 229430 13705
rect 229374 13631 229430 13640
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 13631
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 76978
rect 240140 76968 240192 76974
rect 240140 76910 240192 76916
rect 247038 76936 247094 76945
rect 233240 46368 233292 46374
rect 233240 46310 233292 46316
rect 233252 16574 233280 46310
rect 237380 31272 237432 31278
rect 237380 31214 237432 31220
rect 236000 25696 236052 25702
rect 236000 25638 236052 25644
rect 236012 16574 236040 25638
rect 237392 16574 237420 31214
rect 233252 16546 233464 16574
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 233436 480 233464 16546
rect 234620 4956 234672 4962
rect 234620 4898 234672 4904
rect 234632 480 234660 4898
rect 235816 4072 235868 4078
rect 235816 4014 235868 4020
rect 235828 480 235856 4014
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239312 4004 239364 4010
rect 239312 3946 239364 3952
rect 239324 480 239352 3946
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 76910
rect 247038 76871 247094 76880
rect 244278 74080 244334 74089
rect 244278 74015 244334 74024
rect 242990 40760 243046 40769
rect 242990 40695 243046 40704
rect 241520 20256 241572 20262
rect 241520 20198 241572 20204
rect 241532 16574 241560 20198
rect 243004 16574 243032 40695
rect 244292 16574 244320 74015
rect 247052 16574 247080 76871
rect 251180 73908 251232 73914
rect 251180 73850 251232 73856
rect 249800 68740 249852 68746
rect 249800 68682 249852 68688
rect 248418 19952 248474 19961
rect 248418 19887 248474 19896
rect 241532 16546 241744 16574
rect 243004 16546 244136 16574
rect 244292 16546 245240 16574
rect 247052 16546 247632 16574
rect 241716 480 241744 16546
rect 242900 3936 242952 3942
rect 242900 3878 242952 3884
rect 242912 480 242940 3878
rect 244108 480 244136 16546
rect 245212 480 245240 16546
rect 246394 3496 246450 3505
rect 246394 3431 246450 3440
rect 246408 480 246436 3431
rect 247604 480 247632 16546
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 354 248460 19887
rect 249812 16574 249840 68682
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 3942 251220 73850
rect 251272 25628 251324 25634
rect 251272 25570 251324 25576
rect 251180 3936 251232 3942
rect 251180 3878 251232 3884
rect 251284 3482 251312 25570
rect 252572 16574 252600 80242
rect 288440 79280 288492 79286
rect 288440 79222 288492 79228
rect 255964 78396 256016 78402
rect 255964 78338 256016 78344
rect 255976 20058 256004 78338
rect 260840 76900 260892 76906
rect 260840 76842 260892 76848
rect 256700 64388 256752 64394
rect 256700 64330 256752 64336
rect 255320 20052 255372 20058
rect 255320 19994 255372 20000
rect 255964 20052 256016 20058
rect 255964 19994 256016 20000
rect 255332 16574 255360 19994
rect 252572 16546 253520 16574
rect 255332 16546 255912 16574
rect 252376 3936 252428 3942
rect 252376 3878 252428 3884
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3878
rect 253492 480 253520 16546
rect 254216 14816 254268 14822
rect 254216 14758 254268 14764
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 14758
rect 255884 480 255912 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 64330
rect 259460 61600 259512 61606
rect 259460 61542 259512 61548
rect 258080 26988 258132 26994
rect 258080 26930 258132 26936
rect 258092 16574 258120 26930
rect 258092 16546 258304 16574
rect 258276 480 258304 16546
rect 259472 3942 259500 61542
rect 259552 49292 259604 49298
rect 259552 49234 259604 49240
rect 259460 3936 259512 3942
rect 259460 3878 259512 3884
rect 259564 3482 259592 49234
rect 260852 16574 260880 76842
rect 267740 76832 267792 76838
rect 267740 76774 267792 76780
rect 282918 76800 282974 76809
rect 263598 57488 263654 57497
rect 263598 57423 263654 57432
rect 262220 20188 262272 20194
rect 262220 20130 262272 20136
rect 262232 16574 262260 20130
rect 263612 16574 263640 57423
rect 266358 42120 266414 42129
rect 266358 42055 266414 42064
rect 266372 16574 266400 42055
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 263612 16546 264192 16574
rect 266372 16546 266584 16574
rect 260656 3936 260708 3942
rect 260656 3878 260708 3884
rect 259472 3454 259592 3482
rect 259472 480 259500 3454
rect 260668 480 260696 3878
rect 261772 480 261800 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264164 480 264192 16546
rect 264978 13560 265034 13569
rect 264978 13495 265034 13504
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 13495
rect 266556 480 266584 16546
rect 267752 480 267780 76774
rect 282918 76735 282974 76744
rect 284300 76764 284352 76770
rect 282932 16574 282960 76735
rect 284300 76706 284352 76712
rect 282932 16546 283144 16574
rect 280710 12336 280766 12345
rect 273260 12300 273312 12306
rect 280710 12271 280766 12280
rect 273260 12242 273312 12248
rect 272432 9648 272484 9654
rect 272432 9590 272484 9596
rect 268844 8900 268896 8906
rect 268844 8842 268896 8848
rect 268856 480 268884 8842
rect 270040 6044 270092 6050
rect 270040 5986 270092 5992
rect 270052 480 270080 5986
rect 271236 3868 271288 3874
rect 271236 3810 271288 3816
rect 271248 480 271276 3810
rect 272444 480 272472 9590
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 12242
rect 276664 12232 276716 12238
rect 276664 12174 276716 12180
rect 276020 9580 276072 9586
rect 276020 9522 276072 9528
rect 274824 6112 274876 6118
rect 274824 6054 274876 6060
rect 274836 480 274864 6054
rect 276032 480 276060 9522
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 12174
rect 279514 9208 279570 9217
rect 279514 9143 279570 9152
rect 278320 6860 278372 6866
rect 278320 6802 278372 6808
rect 278332 480 278360 6802
rect 279528 480 279556 9143
rect 280724 480 280752 12271
rect 281906 6352 281962 6361
rect 281906 6287 281962 6296
rect 281920 480 281948 6287
rect 283116 480 283144 16546
rect 284312 3874 284340 76706
rect 285680 43580 285732 43586
rect 285680 43522 285732 43528
rect 285692 16574 285720 43522
rect 288452 16574 288480 79222
rect 293972 79082 294000 83438
rect 320180 80232 320232 80238
rect 320180 80174 320232 80180
rect 293960 79076 294012 79082
rect 293960 79018 294012 79024
rect 315304 78328 315356 78334
rect 315304 78270 315356 78276
rect 296720 76696 296772 76702
rect 296720 76638 296772 76644
rect 292580 65748 292632 65754
rect 292580 65690 292632 65696
rect 289820 45008 289872 45014
rect 289820 44950 289872 44956
rect 285692 16546 286640 16574
rect 288452 16546 289032 16574
rect 284390 14784 284446 14793
rect 284390 14719 284446 14728
rect 284300 3868 284352 3874
rect 284300 3810 284352 3816
rect 284404 3482 284432 14719
rect 285036 3868 285088 3874
rect 285036 3810 285088 3816
rect 284312 3454 284432 3482
rect 284312 480 284340 3454
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285048 354 285076 3810
rect 286612 480 286640 16546
rect 287336 12164 287388 12170
rect 287336 12106 287388 12112
rect 285374 354 285486 480
rect 285048 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 12106
rect 289004 480 289032 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 44950
rect 291200 32496 291252 32502
rect 291200 32438 291252 32444
rect 291212 16574 291240 32438
rect 291212 16546 291424 16574
rect 291396 480 291424 16546
rect 292592 480 292620 65690
rect 295340 60172 295392 60178
rect 295340 60114 295392 60120
rect 293960 32428 294012 32434
rect 293960 32370 294012 32376
rect 292672 24200 292724 24206
rect 292672 24142 292724 24148
rect 292684 16574 292712 24142
rect 293972 16574 294000 32370
rect 295352 16574 295380 60114
rect 296732 16574 296760 76638
rect 302240 76628 302292 76634
rect 302240 76570 302292 76576
rect 298098 73944 298154 73953
rect 298098 73879 298154 73888
rect 292684 16546 293264 16574
rect 293972 16546 294920 16574
rect 295352 16546 295656 16574
rect 296732 16546 297312 16574
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 297284 480 297312 16546
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 73879
rect 299478 55856 299534 55865
rect 299478 55791 299534 55800
rect 299492 3482 299520 55791
rect 299570 25664 299626 25673
rect 299570 25599 299626 25608
rect 299584 3874 299612 25599
rect 302252 16574 302280 76570
rect 302252 16546 303200 16574
rect 301502 10704 301558 10713
rect 301502 10639 301558 10648
rect 299572 3868 299624 3874
rect 299572 3810 299624 3816
rect 300768 3868 300820 3874
rect 300768 3810 300820 3816
rect 299492 3454 299704 3482
rect 299676 480 299704 3454
rect 300780 480 300808 3810
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 10639
rect 303172 480 303200 16546
rect 305552 14748 305604 14754
rect 305552 14690 305604 14696
rect 304356 9512 304408 9518
rect 304356 9454 304408 9460
rect 304368 480 304396 9454
rect 305564 480 305592 14690
rect 307760 14680 307812 14686
rect 307760 14622 307812 14628
rect 306748 3800 306800 3806
rect 306748 3742 306800 3748
rect 306760 480 306788 3742
rect 307772 3398 307800 14622
rect 315316 14618 315344 78270
rect 318798 76664 318854 76673
rect 318798 76599 318854 76608
rect 316038 17232 316094 17241
rect 316038 17167 316094 17176
rect 316052 16574 316080 17167
rect 318812 16574 318840 76599
rect 320192 16574 320220 80174
rect 324320 79144 324372 79150
rect 324320 79086 324372 79092
rect 322940 75540 322992 75546
rect 322940 75482 322992 75488
rect 321560 28416 321612 28422
rect 321560 28358 321612 28364
rect 321572 16574 321600 28358
rect 316052 16546 316264 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 312176 14612 312228 14618
rect 312176 14554 312228 14560
rect 315304 14612 315356 14618
rect 315304 14554 315356 14560
rect 311440 12096 311492 12102
rect 311440 12038 311492 12044
rect 307944 9444 307996 9450
rect 307944 9386 307996 9392
rect 307760 3392 307812 3398
rect 307760 3334 307812 3340
rect 307956 480 307984 9386
rect 310244 6792 310296 6798
rect 310244 6734 310296 6740
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 310256 480 310284 6734
rect 311452 480 311480 12038
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 14554
rect 314660 12028 314712 12034
rect 314660 11970 314712 11976
rect 313832 6724 313884 6730
rect 313832 6666 313884 6672
rect 313844 480 313872 6666
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 11970
rect 316236 480 316264 16546
rect 318062 12200 318118 12209
rect 318062 12135 318118 12144
rect 317326 6216 317382 6225
rect 317326 6151 317382 6160
rect 317340 480 317368 6151
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 12135
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 75482
rect 324332 3210 324360 79086
rect 367756 79014 367784 123626
rect 367744 79008 367796 79014
rect 367744 78950 367796 78956
rect 393976 78946 394004 231814
rect 394160 230518 394188 232358
rect 396460 231198 396488 240042
rect 396448 231192 396500 231198
rect 396448 231134 396500 231140
rect 394148 230512 394200 230518
rect 394148 230454 394200 230460
rect 396552 228410 396580 469202
rect 396540 228404 396592 228410
rect 396540 228346 396592 228352
rect 396644 106282 396672 700266
rect 396724 430636 396776 430642
rect 396724 430578 396776 430584
rect 396632 106276 396684 106282
rect 396632 106218 396684 106224
rect 393964 78940 394016 78946
rect 393964 78882 394016 78888
rect 341524 78260 341576 78266
rect 341524 78202 341576 78208
rect 325700 72820 325752 72826
rect 325700 72762 325752 72768
rect 324412 29844 324464 29850
rect 324412 29786 324464 29792
rect 324424 3398 324452 29786
rect 325712 16574 325740 72762
rect 332600 72752 332652 72758
rect 332600 72694 332652 72700
rect 327080 58948 327132 58954
rect 327080 58890 327132 58896
rect 327092 16574 327120 58890
rect 331220 55956 331272 55962
rect 331220 55898 331272 55904
rect 328460 22976 328512 22982
rect 328460 22918 328512 22924
rect 328472 16574 328500 22918
rect 325712 16546 326384 16574
rect 327092 16546 328040 16574
rect 328472 16546 328776 16574
rect 324412 3392 324464 3398
rect 324412 3334 324464 3340
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324332 3182 324452 3210
rect 324424 480 324452 3182
rect 325620 480 325648 3334
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328012 480 328040 16546
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330392 7676 330444 7682
rect 330392 7618 330444 7624
rect 330404 480 330432 7618
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 55898
rect 332612 3398 332640 72694
rect 341536 72690 341564 78202
rect 396736 77586 396764 430578
rect 397000 404320 397052 404326
rect 397000 404262 397052 404268
rect 396816 378208 396868 378214
rect 396816 378150 396868 378156
rect 396828 78606 396856 378150
rect 396908 271924 396960 271930
rect 396908 271866 396960 271872
rect 396920 80617 396948 271866
rect 397012 232422 397040 404262
rect 397000 232416 397052 232422
rect 397000 232358 397052 232364
rect 396906 80608 396962 80617
rect 396906 80543 396962 80552
rect 397472 78713 397500 703520
rect 413664 700466 413692 703520
rect 405004 700460 405056 700466
rect 405004 700402 405056 700408
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 397552 700392 397604 700398
rect 397552 700334 397604 700340
rect 403624 700392 403676 700398
rect 403624 700334 403676 700340
rect 397564 231130 397592 700334
rect 400864 700324 400916 700330
rect 400864 700266 400916 700272
rect 399484 683188 399536 683194
rect 399484 683130 399536 683136
rect 397552 231124 397604 231130
rect 397552 231066 397604 231072
rect 399496 100706 399524 683130
rect 399576 244316 399628 244322
rect 399576 244258 399628 244264
rect 399588 152522 399616 244258
rect 399576 152516 399628 152522
rect 399576 152458 399628 152464
rect 400876 102134 400904 700266
rect 400956 298172 401008 298178
rect 400956 298114 401008 298120
rect 400968 153882 400996 298114
rect 400956 153876 401008 153882
rect 400956 153818 401008 153824
rect 403636 103494 403664 700334
rect 405016 104854 405044 700402
rect 413284 670744 413336 670750
rect 413284 670686 413336 670692
rect 410524 418192 410576 418198
rect 410524 418134 410576 418140
rect 409144 364404 409196 364410
rect 409144 364346 409196 364352
rect 407764 311908 407816 311914
rect 407764 311850 407816 311856
rect 406384 258120 406436 258126
rect 406384 258062 406436 258068
rect 405004 104848 405056 104854
rect 405004 104790 405056 104796
rect 403624 103488 403676 103494
rect 403624 103430 403676 103436
rect 400864 102128 400916 102134
rect 400864 102070 400916 102076
rect 399484 100700 399536 100706
rect 399484 100642 399536 100648
rect 406396 89690 406424 258062
rect 407776 91050 407804 311850
rect 409156 92478 409184 364346
rect 410536 93838 410564 418134
rect 413296 141438 413324 670686
rect 417424 404388 417476 404394
rect 417424 404330 417476 404336
rect 414664 351960 414716 351966
rect 414664 351902 414716 351908
rect 414676 155242 414704 351902
rect 417436 156670 417464 404330
rect 417424 156664 417476 156670
rect 417424 156606 417476 156612
rect 414664 155236 414716 155242
rect 414664 155178 414716 155184
rect 429212 149734 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 429200 149728 429252 149734
rect 429200 149670 429252 149676
rect 413284 141432 413336 141438
rect 413284 141374 413336 141380
rect 410524 93832 410576 93838
rect 410524 93774 410576 93780
rect 409144 92472 409196 92478
rect 409144 92414 409196 92420
rect 407764 91044 407816 91050
rect 407764 90986 407816 90992
rect 406384 89684 406436 89690
rect 406384 89626 406436 89632
rect 426440 80164 426492 80170
rect 426440 80106 426492 80112
rect 397458 78704 397514 78713
rect 397458 78639 397514 78648
rect 396816 78600 396868 78606
rect 396816 78542 396868 78548
rect 396724 77580 396776 77586
rect 396724 77522 396776 77528
rect 374000 76560 374052 76566
rect 374000 76502 374052 76508
rect 361580 75472 361632 75478
rect 361580 75414 361632 75420
rect 357440 73840 357492 73846
rect 357440 73782 357492 73788
rect 340880 72684 340932 72690
rect 340880 72626 340932 72632
rect 341524 72684 341576 72690
rect 341524 72626 341576 72632
rect 332692 68604 332744 68610
rect 332692 68546 332744 68552
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 68546
rect 333978 62928 334034 62937
rect 333978 62863 334034 62872
rect 333992 16574 334020 62863
rect 339500 29776 339552 29782
rect 339500 29718 339552 29724
rect 333992 16546 334664 16574
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336278 12064 336334 12073
rect 336278 11999 336334 12008
rect 336292 480 336320 11999
rect 337014 10568 337070 10577
rect 337014 10503 337070 10512
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 10503
rect 338672 6588 338724 6594
rect 338672 6530 338724 6536
rect 338684 480 338712 6530
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 29718
rect 340892 16574 340920 72626
rect 347780 72616 347832 72622
rect 347780 72558 347832 72564
rect 345020 40792 345072 40798
rect 345020 40734 345072 40740
rect 343640 20120 343692 20126
rect 343640 20062 343692 20068
rect 343652 16574 343680 20062
rect 345032 16574 345060 40734
rect 346400 29708 346452 29714
rect 346400 29650 346452 29656
rect 346412 16574 346440 29650
rect 347792 16574 347820 72558
rect 356060 67040 356112 67046
rect 356060 66982 356112 66988
rect 349160 54664 349212 54670
rect 349160 54606 349212 54612
rect 340892 16546 341012 16574
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 340984 480 341012 16546
rect 342904 16176 342956 16182
rect 342904 16118 342956 16124
rect 342168 6656 342220 6662
rect 342168 6598 342220 6604
rect 342180 480 342208 6598
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16118
rect 344572 480 344600 16546
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349172 3210 349200 54606
rect 351918 53408 351974 53417
rect 351918 53343 351974 53352
rect 350538 21448 350594 21457
rect 350538 21383 350594 21392
rect 350552 16574 350580 21383
rect 351932 16574 351960 53343
rect 353300 50720 353352 50726
rect 353300 50662 353352 50668
rect 353312 16574 353340 50662
rect 354678 21312 354734 21321
rect 354678 21247 354734 21256
rect 354692 16574 354720 21247
rect 356072 16574 356100 66982
rect 350552 16546 351224 16574
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 356072 16546 356376 16574
rect 349250 15872 349306 15881
rect 349250 15807 349306 15816
rect 349264 3398 349292 15807
rect 349252 3392 349304 3398
rect 349252 3334 349304 3340
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 349172 3182 349292 3210
rect 349264 480 349292 3182
rect 350460 480 350488 3334
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352852 480 352880 16546
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356348 480 356376 16546
rect 357452 3398 357480 73782
rect 358820 58880 358872 58886
rect 358820 58822 358872 58828
rect 357532 39500 357584 39506
rect 357532 39442 357584 39448
rect 357440 3392 357492 3398
rect 357440 3334 357492 3340
rect 357544 480 357572 39442
rect 358832 16574 358860 58822
rect 360200 28348 360252 28354
rect 360200 28290 360252 28296
rect 360212 16574 360240 28290
rect 361592 16574 361620 75414
rect 368480 72548 368532 72554
rect 368480 72490 368532 72496
rect 367100 71324 367152 71330
rect 367100 71266 367152 71272
rect 362960 54596 363012 54602
rect 362960 54538 363012 54544
rect 362972 16574 363000 54538
rect 365720 51808 365772 51814
rect 365720 51750 365772 51756
rect 358832 16546 359504 16574
rect 360212 16546 361160 16574
rect 361592 16546 361896 16574
rect 362972 16546 363552 16574
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358740 480 358768 3334
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 361132 480 361160 16546
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363524 480 363552 16546
rect 364616 6520 364668 6526
rect 364616 6462 364668 6468
rect 364628 480 364656 6462
rect 365732 3398 365760 51750
rect 367112 16574 367140 71266
rect 368492 16574 368520 72490
rect 369858 37904 369914 37913
rect 369858 37839 369914 37848
rect 369872 16574 369900 37839
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 369872 16546 370176 16574
rect 365810 14648 365866 14657
rect 365810 14583 365866 14592
rect 365720 3392 365772 3398
rect 365720 3334 365772 3340
rect 365824 480 365852 14583
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367020 480 367048 3334
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 372894 14512 372950 14521
rect 372894 14447 372950 14456
rect 371238 13424 371294 13433
rect 371238 13359 371294 13368
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 13359
rect 372908 480 372936 14447
rect 374012 1170 374040 76502
rect 402978 75440 403034 75449
rect 402978 75375 403034 75384
rect 382280 72480 382332 72486
rect 382280 72422 382332 72428
rect 375380 70032 375432 70038
rect 375380 69974 375432 69980
rect 374092 66972 374144 66978
rect 374092 66914 374144 66920
rect 374104 3398 374132 66914
rect 375392 16574 375420 69974
rect 380900 61532 380952 61538
rect 380900 61474 380952 61480
rect 376760 60104 376812 60110
rect 376760 60046 376812 60052
rect 376772 16574 376800 60046
rect 378140 26920 378192 26926
rect 378140 26862 378192 26868
rect 378152 16574 378180 26862
rect 379520 21548 379572 21554
rect 379520 21490 379572 21496
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 378152 16546 378456 16574
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374012 1142 374132 1170
rect 374104 480 374132 1142
rect 375300 480 375328 3334
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 21490
rect 380912 16574 380940 61474
rect 380912 16546 381216 16574
rect 381188 480 381216 16546
rect 382292 3398 382320 72422
rect 382372 71256 382424 71262
rect 382372 71198 382424 71204
rect 382280 3392 382332 3398
rect 382280 3334 382332 3340
rect 382384 480 382412 71198
rect 390560 65680 390612 65686
rect 390560 65622 390612 65628
rect 383660 55888 383712 55894
rect 383660 55830 383712 55836
rect 383672 16574 383700 55830
rect 389180 49224 389232 49230
rect 389180 49166 389232 49172
rect 387798 44840 387854 44849
rect 387798 44775 387854 44784
rect 386418 26888 386474 26897
rect 386418 26823 386474 26832
rect 385040 25560 385092 25566
rect 385040 25502 385092 25508
rect 385052 16574 385080 25502
rect 386432 16574 386460 26823
rect 383672 16546 384344 16574
rect 385052 16546 386000 16574
rect 386432 16546 386736 16574
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 383580 480 383608 3334
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 16546
rect 385972 480 386000 16546
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 44775
rect 389192 16574 389220 49166
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 3398 390600 65622
rect 396080 65612 396132 65618
rect 396080 65554 396132 65560
rect 390652 60036 390704 60042
rect 390652 59978 390704 59984
rect 390560 3392 390612 3398
rect 390560 3334 390612 3340
rect 390664 480 390692 59978
rect 394700 57248 394752 57254
rect 394700 57190 394752 57196
rect 391940 46300 391992 46306
rect 391940 46242 391992 46248
rect 391952 16574 391980 46242
rect 394712 16574 394740 57190
rect 391952 16546 392624 16574
rect 394712 16546 395384 16574
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391860 480 391888 3334
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394240 6452 394292 6458
rect 394240 6394 394292 6400
rect 394252 480 394280 6394
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 65554
rect 398840 54528 398892 54534
rect 398840 54470 398892 54476
rect 397460 44940 397512 44946
rect 397460 44882 397512 44888
rect 397472 16574 397500 44882
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398852 3210 398880 54470
rect 401600 50652 401652 50658
rect 401600 50594 401652 50600
rect 400220 19984 400272 19990
rect 400220 19926 400272 19932
rect 400232 16574 400260 19926
rect 401612 16574 401640 50594
rect 402992 16574 403020 75375
rect 412640 64320 412692 64326
rect 412640 64262 412692 64268
rect 408500 62892 408552 62898
rect 408500 62834 408552 62840
rect 405738 29608 405794 29617
rect 405738 29543 405794 29552
rect 404360 21480 404412 21486
rect 404360 21422 404412 21428
rect 400232 16546 400904 16574
rect 401612 16546 402560 16574
rect 402992 16546 403664 16574
rect 398932 14544 398984 14550
rect 398932 14486 398984 14492
rect 398944 3398 398972 14486
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 398852 3182 398972 3210
rect 398944 480 398972 3182
rect 400140 480 400168 3334
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 402532 480 402560 16546
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 21422
rect 405752 16574 405780 29543
rect 407118 24304 407174 24313
rect 407118 24239 407174 24248
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 3210 407160 24239
rect 407210 24168 407266 24177
rect 407210 24103 407266 24112
rect 407224 3398 407252 24103
rect 408512 16574 408540 62834
rect 409880 39432 409932 39438
rect 409880 39374 409932 39380
rect 409892 16574 409920 39374
rect 408512 16546 409184 16574
rect 409892 16546 410840 16574
rect 407212 3392 407264 3398
rect 407212 3334 407264 3340
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 407132 3182 407252 3210
rect 407224 480 407252 3182
rect 408420 480 408448 3334
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410812 480 410840 16546
rect 411904 9376 411956 9382
rect 411904 9318 411956 9324
rect 411916 480 411944 9318
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 64262
rect 415400 51740 415452 51746
rect 415400 51682 415452 51688
rect 414296 9308 414348 9314
rect 414296 9250 414348 9256
rect 414308 480 414336 9250
rect 415412 1970 415440 51682
rect 425060 49156 425112 49162
rect 425060 49098 425112 49104
rect 423678 48920 423734 48929
rect 423678 48855 423734 48864
rect 415492 42152 415544 42158
rect 415492 42094 415544 42100
rect 415400 1964 415452 1970
rect 415400 1906 415452 1912
rect 415504 480 415532 42094
rect 419540 38004 419592 38010
rect 419540 37946 419592 37952
rect 418160 28280 418212 28286
rect 418160 28222 418212 28228
rect 416780 22908 416832 22914
rect 416780 22850 416832 22856
rect 416792 16574 416820 22850
rect 418172 16574 418200 28222
rect 419552 16574 419580 37946
rect 422298 22672 422354 22681
rect 422298 22607 422354 22616
rect 422312 16574 422340 22607
rect 423692 16574 423720 48855
rect 425072 16574 425100 49098
rect 426452 16574 426480 80106
rect 462332 80073 462360 703520
rect 478524 700398 478552 703520
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 494072 145586 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 526444 524476 526496 524482
rect 526444 524418 526496 524424
rect 525064 470620 525116 470626
rect 525064 470562 525116 470568
rect 494060 145580 494112 145586
rect 494060 145522 494112 145528
rect 525076 95198 525104 470562
rect 526456 96626 526484 524418
rect 526444 96620 526496 96626
rect 526444 96562 526496 96568
rect 525064 95192 525116 95198
rect 525064 95134 525116 95140
rect 462318 80064 462374 80073
rect 462318 79999 462374 80008
rect 498200 79892 498252 79898
rect 498200 79834 498252 79840
rect 430580 78872 430632 78878
rect 430580 78814 430632 78820
rect 427820 29640 427872 29646
rect 427820 29582 427872 29588
rect 427832 16574 427860 29582
rect 429200 18760 429252 18766
rect 429200 18702 429252 18708
rect 416792 16546 417464 16574
rect 418172 16546 418568 16574
rect 419552 16546 420224 16574
rect 422312 16546 422616 16574
rect 423692 16546 423812 16574
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 416688 1964 416740 1970
rect 416688 1906 416740 1912
rect 416700 480 416728 1906
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420196 480 420224 16546
rect 421378 4992 421434 5001
rect 421378 4927 421434 4936
rect 421392 480 421420 4927
rect 422588 480 422616 16546
rect 423784 480 423812 16546
rect 424966 7712 425022 7721
rect 424966 7647 425022 7656
rect 424980 480 425008 7647
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 18702
rect 430592 16574 430620 78814
rect 480260 78192 480312 78198
rect 480260 78134 480312 78140
rect 438860 75404 438912 75410
rect 438860 75346 438912 75352
rect 437480 69964 437532 69970
rect 437480 69906 437532 69912
rect 431960 68536 432012 68542
rect 431960 68478 432012 68484
rect 430592 16546 430896 16574
rect 430868 480 430896 16546
rect 431972 1986 432000 68478
rect 433340 58812 433392 58818
rect 433340 58754 433392 58760
rect 432052 43512 432104 43518
rect 432052 43454 432104 43460
rect 432064 2106 432092 43454
rect 433352 16574 433380 58754
rect 436100 47796 436152 47802
rect 436100 47738 436152 47744
rect 436112 16574 436140 47738
rect 433352 16546 434024 16574
rect 436112 16546 436784 16574
rect 432052 2100 432104 2106
rect 432052 2042 432104 2048
rect 433248 2100 433300 2106
rect 433248 2042 433300 2048
rect 431972 1958 432092 1986
rect 432064 480 432092 1958
rect 433260 480 433288 2042
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 435088 11960 435140 11966
rect 435088 11902 435140 11908
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 11902
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 69906
rect 438872 16574 438900 75346
rect 459558 75304 459614 75313
rect 459558 75239 459614 75248
rect 444380 64252 444432 64258
rect 444380 64194 444432 64200
rect 440240 62824 440292 62830
rect 440240 62766 440292 62772
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 1970 440280 62766
rect 440330 59936 440386 59945
rect 440330 59871 440386 59880
rect 440240 1964 440292 1970
rect 440240 1906 440292 1912
rect 440344 480 440372 59871
rect 444392 16574 444420 64194
rect 449898 57352 449954 57361
rect 449898 57287 449954 57296
rect 448520 50584 448572 50590
rect 448520 50526 448572 50532
rect 445760 17468 445812 17474
rect 445760 17410 445812 17416
rect 444392 16546 445064 16574
rect 442630 10432 442686 10441
rect 442630 10367 442686 10376
rect 441528 1964 441580 1970
rect 441528 1906 441580 1912
rect 441540 480 441568 1906
rect 442644 480 442672 10367
rect 443366 10296 443422 10305
rect 443366 10231 443422 10240
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 10231
rect 445036 480 445064 16546
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 17410
rect 447416 11892 447468 11898
rect 447416 11834 447468 11840
rect 447428 480 447456 11834
rect 448532 3210 448560 50526
rect 449912 16574 449940 57287
rect 458178 54496 458234 54505
rect 458178 54431 458234 54440
rect 455420 53236 455472 53242
rect 455420 53178 455472 53184
rect 451280 47728 451332 47734
rect 451280 47670 451332 47676
rect 451292 16574 451320 47670
rect 452660 17400 452712 17406
rect 452660 17342 452712 17348
rect 452672 16574 452700 17342
rect 455432 16574 455460 53178
rect 456800 20052 456852 20058
rect 456800 19994 456852 20000
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 455432 16546 455736 16574
rect 448612 16108 448664 16114
rect 448612 16050 448664 16056
rect 448624 3398 448652 16050
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 454040 16040 454092 16046
rect 454040 15982 454092 15988
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 15982
rect 455708 480 455736 16546
rect 456812 1970 456840 19994
rect 458192 16574 458220 54431
rect 459572 16574 459600 75239
rect 465080 72684 465132 72690
rect 465080 72626 465132 72632
rect 465092 16574 465120 72626
rect 480272 16574 480300 78134
rect 483018 77888 483074 77897
rect 483018 77823 483074 77832
rect 481640 68468 481692 68474
rect 481640 68410 481692 68416
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 465092 16546 465212 16574
rect 480272 16546 480576 16574
rect 456890 13288 456946 13297
rect 456890 13223 456946 13232
rect 456800 1964 456852 1970
rect 456800 1906 456852 1912
rect 456904 480 456932 13223
rect 458088 1964 458140 1970
rect 458088 1906 458140 1912
rect 458100 480 458128 1906
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 463976 11824 464028 11830
rect 463976 11766 464028 11772
rect 462780 6384 462832 6390
rect 462780 6326 462832 6332
rect 461584 3664 461636 3670
rect 461584 3606 461636 3612
rect 461596 480 461624 3606
rect 462792 480 462820 6326
rect 463988 480 464016 11766
rect 465184 480 465212 16546
rect 475752 14612 475804 14618
rect 475752 14554 475804 14560
rect 474094 11928 474150 11937
rect 474094 11863 474150 11872
rect 470600 11756 470652 11762
rect 470600 11698 470652 11704
rect 466276 9240 466328 9246
rect 466276 9182 466328 9188
rect 466288 480 466316 9182
rect 469864 9172 469916 9178
rect 469864 9114 469916 9120
rect 467472 6316 467524 6322
rect 467472 6258 467524 6264
rect 467484 480 467512 6258
rect 468668 3732 468720 3738
rect 468668 3674 468720 3680
rect 468680 480 468708 3674
rect 469876 480 469904 9114
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 11698
rect 473452 9104 473504 9110
rect 473452 9046 473504 9052
rect 472256 3596 472308 3602
rect 472256 3538 472308 3544
rect 472268 480 472296 3538
rect 473464 480 473492 9046
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 11863
rect 475764 480 475792 14554
rect 478142 11792 478198 11801
rect 478142 11727 478198 11736
rect 476946 9072 477002 9081
rect 476946 9007 477002 9016
rect 476960 480 476988 9007
rect 478156 480 478184 11727
rect 479340 3528 479392 3534
rect 479340 3470 479392 3476
rect 479352 480 479380 3470
rect 480548 480 480576 16546
rect 481652 3534 481680 68410
rect 481732 61464 481784 61470
rect 481732 61406 481784 61412
rect 481640 3528 481692 3534
rect 481640 3470 481692 3476
rect 481744 480 481772 61406
rect 483032 16574 483060 77823
rect 490012 75336 490064 75342
rect 490012 75278 490064 75284
rect 488540 53168 488592 53174
rect 488540 53110 488592 53116
rect 484400 47660 484452 47666
rect 484400 47602 484452 47608
rect 484412 16574 484440 47602
rect 487160 35216 487212 35222
rect 487160 35158 487212 35164
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 482468 3528 482520 3534
rect 482468 3470 482520 3476
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482480 354 482508 3470
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486424 4888 486476 4894
rect 486424 4830 486476 4836
rect 486436 480 486464 4830
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 35158
rect 488552 16574 488580 53110
rect 488552 16546 488856 16574
rect 488828 480 488856 16546
rect 490024 6914 490052 75278
rect 496818 75168 496874 75177
rect 496818 75103 496874 75112
rect 494058 57216 494114 57225
rect 494058 57151 494114 57160
rect 491300 46232 491352 46238
rect 491300 46174 491352 46180
rect 491312 16574 491340 46174
rect 492680 17332 492732 17338
rect 492680 17274 492732 17280
rect 492692 16574 492720 17274
rect 494072 16574 494100 57151
rect 496832 16574 496860 75103
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 496832 16546 497136 16574
rect 489932 6886 490052 6914
rect 489932 480 489960 6886
rect 491116 3460 491168 3466
rect 491116 3402 491168 3408
rect 491128 480 491156 3402
rect 492324 480 492352 16546
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 495898 4856 495954 4865
rect 495898 4791 495954 4800
rect 495912 480 495940 4791
rect 497108 480 497136 16546
rect 498212 480 498240 79834
rect 514760 79824 514812 79830
rect 514760 79766 514812 79772
rect 506480 75268 506532 75274
rect 506480 75210 506532 75216
rect 505100 71188 505152 71194
rect 505100 71130 505152 71136
rect 498292 49088 498344 49094
rect 498292 49030 498344 49036
rect 498304 16574 498332 49030
rect 503720 37936 503772 37942
rect 503720 37878 503772 37884
rect 499580 31204 499632 31210
rect 499580 31146 499632 31152
rect 499592 16574 499620 31146
rect 498304 16546 498976 16574
rect 499592 16546 500632 16574
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500604 480 500632 16546
rect 502984 6248 503036 6254
rect 502984 6190 503036 6196
rect 501786 3360 501842 3369
rect 501786 3295 501842 3304
rect 501800 480 501828 3295
rect 502996 480 503024 6190
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 37878
rect 505112 16574 505140 71130
rect 506492 16574 506520 75210
rect 511998 64152 512054 64161
rect 511998 64087 512054 64096
rect 507860 58744 507912 58750
rect 507860 58686 507912 58692
rect 507872 16574 507900 58686
rect 510618 40624 510674 40633
rect 510618 40559 510674 40568
rect 510632 16574 510660 40559
rect 505112 16546 505416 16574
rect 506492 16546 507256 16574
rect 507872 16546 508912 16574
rect 510632 16546 511304 16574
rect 505388 480 505416 16546
rect 506480 7608 506532 7614
rect 506480 7550 506532 7556
rect 506492 480 506520 7550
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 16546
rect 508884 480 508912 16546
rect 510068 9036 510120 9042
rect 510068 8978 510120 8984
rect 510080 480 510108 8978
rect 511276 480 511304 16546
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512012 354 512040 64087
rect 513378 13152 513434 13161
rect 513378 13087 513434 13096
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 13087
rect 514772 3534 514800 79766
rect 527192 77217 527220 703520
rect 543476 700330 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 531964 630692 532016 630698
rect 531964 630634 532016 630640
rect 530584 576904 530636 576910
rect 530584 576846 530636 576852
rect 530596 97986 530624 576846
rect 531976 99346 532004 630634
rect 558932 144226 558960 702406
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580262 644056 580318 644065
rect 580262 643991 580318 644000
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580078 431624 580134 431633
rect 580078 431559 580134 431568
rect 580092 430642 580120 431559
rect 580080 430636 580132 430642
rect 580080 430578 580132 430584
rect 580078 418296 580134 418305
rect 580078 418231 580134 418240
rect 580092 418198 580120 418231
rect 580080 418192 580132 418198
rect 580080 418134 580132 418140
rect 580078 404968 580134 404977
rect 580078 404903 580134 404912
rect 580092 404394 580120 404903
rect 580080 404388 580132 404394
rect 580080 404330 580132 404336
rect 580078 378448 580134 378457
rect 580078 378383 580134 378392
rect 580092 378214 580120 378383
rect 580080 378208 580132 378214
rect 580080 378150 580132 378156
rect 579802 365120 579858 365129
rect 579802 365055 579858 365064
rect 579816 364410 579844 365055
rect 579804 364404 579856 364410
rect 579804 364346 579856 364352
rect 580080 351960 580132 351966
rect 580078 351928 580080 351937
rect 580132 351928 580134 351937
rect 580078 351863 580134 351872
rect 580078 312080 580134 312089
rect 580078 312015 580134 312024
rect 580092 311914 580120 312015
rect 580080 311908 580132 311914
rect 580080 311850 580132 311856
rect 580078 298752 580134 298761
rect 580078 298687 580134 298696
rect 580092 298178 580120 298687
rect 580080 298172 580132 298178
rect 580080 298114 580132 298120
rect 579802 272232 579858 272241
rect 579802 272167 579858 272176
rect 579816 271930 579844 272167
rect 579804 271924 579856 271930
rect 579804 271866 579856 271872
rect 579986 258904 580042 258913
rect 579986 258839 580042 258848
rect 580000 258126 580028 258839
rect 579988 258120 580040 258126
rect 579988 258062 580040 258068
rect 579986 245576 580042 245585
rect 579986 245511 580042 245520
rect 580000 244322 580028 245511
rect 579988 244316 580040 244322
rect 579988 244258 580040 244264
rect 580078 232384 580134 232393
rect 580078 232319 580134 232328
rect 580092 231878 580120 232319
rect 580080 231872 580132 231878
rect 580080 231814 580132 231820
rect 580184 227050 580212 458079
rect 580172 227044 580224 227050
rect 580172 226986 580224 226992
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580184 218074 580212 218991
rect 580172 218068 580224 218074
rect 580172 218010 580224 218016
rect 580170 205728 580226 205737
rect 580170 205663 580172 205672
rect 580224 205663 580226 205672
rect 580172 205634 580224 205640
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 579986 152688 580042 152697
rect 579986 152623 580042 152632
rect 580000 151842 580028 152623
rect 579988 151836 580040 151842
rect 579988 151778 580040 151784
rect 558920 144220 558972 144226
rect 558920 144162 558972 144168
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 580184 138038 580212 139295
rect 580172 138032 580224 138038
rect 580172 137974 580224 137980
rect 579802 126032 579858 126041
rect 579802 125967 579858 125976
rect 579816 125662 579844 125967
rect 579804 125656 579856 125662
rect 579804 125598 579856 125604
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580184 111858 580212 112775
rect 580172 111852 580224 111858
rect 580172 111794 580224 111800
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580184 99414 580212 99447
rect 580172 99408 580224 99414
rect 580172 99350 580224 99356
rect 531964 99340 532016 99346
rect 531964 99282 532016 99288
rect 530584 97980 530636 97986
rect 530584 97922 530636 97928
rect 579986 86184 580042 86193
rect 579986 86119 580042 86128
rect 580000 80782 580028 86119
rect 580276 82142 580304 643991
rect 580722 617536 580778 617545
rect 580722 617471 580778 617480
rect 580354 591016 580410 591025
rect 580354 590951 580410 590960
rect 580264 82136 580316 82142
rect 580264 82078 580316 82084
rect 579988 80776 580040 80782
rect 579988 80718 580040 80724
rect 554780 80368 554832 80374
rect 554780 80310 554832 80316
rect 532700 78124 532752 78130
rect 532700 78066 532752 78072
rect 527178 77208 527234 77217
rect 527178 77143 527234 77152
rect 518900 71120 518952 71126
rect 518900 71062 518952 71068
rect 514850 53272 514906 53281
rect 514850 53207 514906 53216
rect 514760 3528 514812 3534
rect 514760 3470 514812 3476
rect 514864 3346 514892 53207
rect 516140 53100 516192 53106
rect 516140 53042 516192 53048
rect 516152 16574 516180 53042
rect 518912 16574 518940 71062
rect 523040 69896 523092 69902
rect 523040 69838 523092 69844
rect 521660 22840 521712 22846
rect 521660 22782 521712 22788
rect 516152 16546 517192 16574
rect 518912 16546 519584 16574
rect 515588 3528 515640 3534
rect 515588 3470 515640 3476
rect 514772 3318 514892 3346
rect 514772 480 514800 3318
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515600 354 515628 3470
rect 517164 480 517192 16546
rect 517888 15972 517940 15978
rect 517888 15914 517940 15920
rect 515926 354 516038 480
rect 515600 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 15914
rect 519556 480 519584 16546
rect 520280 14476 520332 14482
rect 520280 14418 520332 14424
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 14418
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 22782
rect 523052 480 523080 69838
rect 529938 69592 529994 69601
rect 529938 69527 529994 69536
rect 525800 66904 525852 66910
rect 525800 66846 525852 66852
rect 524420 24132 524472 24138
rect 524420 24074 524472 24080
rect 524432 16574 524460 24074
rect 525812 16574 525840 66846
rect 528558 51776 528614 51785
rect 528558 51711 528614 51720
rect 527180 39364 527232 39370
rect 527180 39306 527232 39312
rect 527192 16574 527220 39306
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 523776 15904 523828 15910
rect 523776 15846 523828 15852
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 15846
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527836 480 527864 16546
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 51711
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 69527
rect 531318 39264 531374 39273
rect 531318 39199 531374 39208
rect 531332 480 531360 39199
rect 531410 25528 531466 25537
rect 531410 25463 531466 25472
rect 531424 16574 531452 25463
rect 532712 16574 532740 78066
rect 538864 78056 538916 78062
rect 538864 77998 538916 78004
rect 536840 69828 536892 69834
rect 536840 69770 536892 69776
rect 534080 50516 534132 50522
rect 534080 50458 534132 50464
rect 534092 16574 534120 50458
rect 535460 31136 535512 31142
rect 535460 31078 535512 31084
rect 535472 16574 535500 31078
rect 536852 16574 536880 69770
rect 531424 16546 532096 16574
rect 532712 16546 533752 16574
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533724 480 533752 16546
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 538876 6254 538904 77998
rect 539600 71052 539652 71058
rect 539600 70994 539652 71000
rect 539612 16574 539640 70994
rect 543740 68400 543792 68406
rect 543740 68342 543792 68348
rect 542360 50448 542412 50454
rect 542360 50390 542412 50396
rect 540980 17264 541032 17270
rect 540980 17206 541032 17212
rect 540992 16574 541020 17206
rect 542372 16574 542400 50390
rect 543752 16574 543780 68342
rect 550640 68332 550692 68338
rect 550640 68274 550692 68280
rect 547878 62792 547934 62801
rect 547878 62727 547934 62736
rect 546498 18592 546554 18601
rect 546498 18527 546554 18536
rect 539612 16546 540376 16574
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 539600 8968 539652 8974
rect 539600 8910 539652 8916
rect 538864 6248 538916 6254
rect 538864 6190 538916 6196
rect 538404 4820 538456 4826
rect 538404 4762 538456 4768
rect 538416 480 538444 4762
rect 539612 480 539640 8910
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540348 354 540376 16546
rect 542004 480 542032 16546
rect 540766 354 540878 480
rect 540348 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545488 6180 545540 6186
rect 545488 6122 545540 6128
rect 545500 480 545528 6122
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 18527
rect 547892 480 547920 62727
rect 549258 46200 549314 46209
rect 549258 46135 549314 46144
rect 549272 16574 549300 46135
rect 550652 16574 550680 68274
rect 552020 49020 552072 49026
rect 552020 48962 552072 48968
rect 552032 16574 552060 48962
rect 553400 44872 553452 44878
rect 553400 44814 553452 44820
rect 553412 16574 553440 44814
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 549074 7576 549130 7585
rect 549074 7511 549130 7520
rect 549088 480 549116 7511
rect 550284 480 550312 16546
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 80310
rect 580368 79422 580396 590951
rect 580538 564360 580594 564369
rect 580538 564295 580594 564304
rect 580446 537840 580502 537849
rect 580446 537775 580502 537784
rect 580460 80850 580488 537775
rect 580552 151094 580580 564295
rect 580630 484664 580686 484673
rect 580630 484599 580686 484608
rect 580540 151088 580592 151094
rect 580540 151030 580592 151036
rect 580448 80844 580500 80850
rect 580448 80786 580500 80792
rect 580644 80646 580672 484599
rect 580736 229770 580764 617471
rect 580814 511320 580870 511329
rect 580814 511255 580870 511264
rect 580724 229764 580776 229770
rect 580724 229706 580776 229712
rect 580828 224262 580856 511255
rect 580906 325272 580962 325281
rect 580906 325207 580962 325216
rect 580816 224256 580868 224262
rect 580816 224198 580868 224204
rect 580722 192536 580778 192545
rect 580722 192471 580778 192480
rect 580736 80714 580764 192471
rect 580724 80708 580776 80714
rect 580724 80650 580776 80656
rect 580632 80640 580684 80646
rect 580632 80582 580684 80588
rect 580356 79416 580408 79422
rect 580356 79358 580408 79364
rect 580920 79354 580948 325207
rect 580908 79348 580960 79354
rect 580908 79290 580960 79296
rect 581000 77988 581052 77994
rect 581000 77930 581052 77936
rect 565818 76528 565874 76537
rect 565818 76463 565874 76472
rect 564440 75200 564492 75206
rect 564440 75142 564492 75148
rect 558920 69760 558972 69766
rect 558920 69702 558972 69708
rect 557540 50380 557592 50386
rect 557540 50322 557592 50328
rect 556160 21412 556212 21418
rect 556160 21354 556212 21360
rect 556172 480 556200 21354
rect 556252 18692 556304 18698
rect 556252 18634 556304 18640
rect 556264 16574 556292 18634
rect 557552 16574 557580 50322
rect 558932 16574 558960 69702
rect 561680 64184 561732 64190
rect 561680 64126 561732 64132
rect 560300 18624 560352 18630
rect 560300 18566 560352 18572
rect 560312 16574 560340 18566
rect 561692 16574 561720 64126
rect 563060 43444 563112 43450
rect 563060 43386 563112 43392
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 43386
rect 564452 480 564480 75142
rect 564532 69692 564584 69698
rect 564532 69634 564584 69640
rect 564544 16574 564572 69634
rect 565832 16574 565860 76463
rect 578238 73808 578294 73817
rect 578238 73743 578294 73752
rect 568580 65544 568632 65550
rect 568580 65486 568632 65492
rect 568592 16574 568620 65486
rect 572720 58676 572772 58682
rect 572720 58618 572772 58624
rect 571340 47592 571392 47598
rect 571340 47534 571392 47540
rect 569960 40724 570012 40730
rect 569960 40666 570012 40672
rect 569972 16574 570000 40666
rect 564544 16546 565216 16574
rect 565832 16546 566872 16574
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 566844 480 566872 16546
rect 567566 13016 567622 13025
rect 567566 12951 567622 12960
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 12951
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 570340 480 570368 16546
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571352 354 571380 47534
rect 572732 480 572760 58618
rect 575478 53136 575534 53145
rect 575478 53071 575534 53080
rect 572812 42084 572864 42090
rect 572812 42026 572864 42032
rect 572824 16574 572852 42026
rect 574100 31068 574152 31074
rect 574100 31010 574152 31016
rect 574112 16574 574140 31010
rect 575492 16574 575520 53071
rect 578252 16574 578280 73743
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580264 61396 580316 61402
rect 580264 61338 580316 61344
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580172 22772 580224 22778
rect 580172 22714 580224 22720
rect 580184 19825 580212 22714
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 572824 16546 573496 16574
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 578252 16546 578648 16574
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 575124 480 575152 16546
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 577410 8936 577466 8945
rect 577410 8871 577466 8880
rect 577424 480 577452 8871
rect 578620 480 578648 16546
rect 580276 6633 580304 61338
rect 581012 16574 581040 77930
rect 581012 16546 581776 16574
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 581000 6248 581052 6254
rect 581000 6190 581052 6196
rect 581012 480 581040 6190
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576278 -960 576390 326
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583390 11656 583446 11665
rect 583390 11591 583446 11600
rect 583404 480 583432 11591
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3330 632068 3332 632088
rect 3332 632068 3384 632088
rect 3384 632068 3386 632088
rect 3330 632032 3386 632068
rect 3330 579944 3386 580000
rect 2962 527856 3018 527912
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 3238 501744 3294 501800
rect 3054 475632 3110 475688
rect 3330 462576 3386 462632
rect 3330 449520 3386 449576
rect 2962 423544 3018 423600
rect 3330 410488 3386 410544
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3330 371320 3386 371376
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 3146 319232 3202 319288
rect 3238 267144 3294 267200
rect 3330 254088 3386 254144
rect 2778 241032 2834 241088
rect 3054 227976 3110 228032
rect 3330 214920 3386 214976
rect 2962 188808 3018 188864
rect 3330 175888 3386 175944
rect 3330 162868 3332 162888
rect 3332 162868 3384 162888
rect 3384 162868 3386 162888
rect 3330 162832 3386 162868
rect 2962 110608 3018 110664
rect 3330 84632 3386 84688
rect 3698 619112 3754 619168
rect 3606 606056 3662 606112
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 3514 97552 3570 97608
rect 3882 566888 3938 566944
rect 3790 553832 3846 553888
rect 3698 201864 3754 201920
rect 4066 306176 4122 306232
rect 3974 293120 4030 293176
rect 3790 79056 3846 79112
rect 3606 78920 3662 78976
rect 3422 78784 3478 78840
rect 6918 79192 6974 79248
rect 4894 78512 4950 78568
rect 17222 77832 17278 77888
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 2870 32408 2926 32464
rect 2778 21256 2834 21312
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3514 19352 3570 19408
rect 3422 6432 3478 6488
rect 20718 76472 20774 76528
rect 19338 35128 19394 35184
rect 43442 79464 43498 79520
rect 37922 79328 37978 79384
rect 19430 7520 19486 7576
rect 37278 74160 37334 74216
rect 35990 71032 36046 71088
rect 40038 71168 40094 71224
rect 41878 8880 41934 8936
rect 57978 73888 58034 73944
rect 55218 68176 55274 68232
rect 57242 9016 57298 9072
rect 75918 72392 75974 72448
rect 73158 69536 73214 69592
rect 74998 9152 75054 9208
rect 93858 76608 93914 76664
rect 91098 68312 91154 68368
rect 92478 10240 92534 10296
rect 117318 137536 117374 137592
rect 117318 136040 117374 136096
rect 117318 134544 117374 134600
rect 117410 133048 117466 133104
rect 117318 131552 117374 131608
rect 117318 130056 117374 130112
rect 117318 128560 117374 128616
rect 117318 127064 117374 127120
rect 117318 125568 117374 125624
rect 117318 124108 117320 124128
rect 117320 124108 117372 124128
rect 117372 124108 117374 124128
rect 117318 124072 117374 124108
rect 117318 122576 117374 122632
rect 117318 121080 117374 121136
rect 117318 119584 117374 119640
rect 117318 118088 117374 118144
rect 117318 116592 117374 116648
rect 117318 115096 117374 115152
rect 117318 113600 117374 113656
rect 117318 112104 117374 112160
rect 117318 110608 117374 110664
rect 117962 103128 118018 103184
rect 118054 89664 118110 89720
rect 118238 95648 118294 95704
rect 118330 94152 118386 94208
rect 118606 109112 118662 109168
rect 118974 106120 119030 106176
rect 118882 104624 118938 104680
rect 118790 100136 118846 100192
rect 118698 98640 118754 98696
rect 118514 92656 118570 92712
rect 118422 91160 118478 91216
rect 118146 88168 118202 88224
rect 118514 86672 118570 86728
rect 118422 83680 118478 83736
rect 118330 82184 118386 82240
rect 109314 7656 109370 7712
rect 113822 78104 113878 78160
rect 111798 76744 111854 76800
rect 118606 85176 118662 85232
rect 118514 80416 118570 80472
rect 120630 108296 120686 108352
rect 120814 102040 120870 102096
rect 120722 97688 120778 97744
rect 143538 200640 143594 200696
rect 147494 196424 147550 196480
rect 153290 196152 153346 196208
rect 139398 195900 139454 195936
rect 139398 195880 139400 195900
rect 139400 195880 139452 195900
rect 139452 195880 139454 195900
rect 142342 195880 142398 195936
rect 153198 195880 153254 195936
rect 138110 195744 138166 195800
rect 140778 195744 140834 195800
rect 150346 195644 150348 195664
rect 150348 195644 150400 195664
rect 150400 195644 150402 195664
rect 150346 195608 150402 195644
rect 153934 195880 153990 195936
rect 155958 195880 156014 195936
rect 158258 195880 158314 195936
rect 158902 195880 158958 195936
rect 163502 199280 163558 199336
rect 161386 195880 161442 195936
rect 159822 195744 159878 195800
rect 153934 194656 153990 194712
rect 155222 194656 155278 194712
rect 151634 193568 151690 193624
rect 153290 193568 153346 193624
rect 149794 190576 149850 190632
rect 166078 196152 166134 196208
rect 144642 186904 144698 186960
rect 146114 180684 146116 180704
rect 146116 180684 146168 180704
rect 146168 180684 146170 180704
rect 146114 180648 146170 180684
rect 148046 179016 148102 179072
rect 142666 178744 142722 178800
rect 135258 173984 135314 174040
rect 137834 173984 137890 174040
rect 142066 176704 142122 176760
rect 144182 174528 144238 174584
rect 156050 174528 156106 174584
rect 145654 173848 145710 173904
rect 142618 173712 142674 173768
rect 142066 171128 142122 171184
rect 142066 170992 142122 171048
rect 142066 161472 142122 161528
rect 143538 142432 143594 142488
rect 142066 142160 142122 142216
rect 148690 173712 148746 173768
rect 146758 173576 146814 173632
rect 146482 143384 146538 143440
rect 148046 143248 148102 143304
rect 149610 143112 149666 143168
rect 151174 142976 151230 143032
rect 151358 142976 151414 143032
rect 151358 142568 151414 142624
rect 160558 142976 160614 143032
rect 164330 166368 164386 166424
rect 166170 196016 166226 196072
rect 166998 166232 167054 166288
rect 171506 142840 171562 142896
rect 173070 142704 173126 142760
rect 179418 126112 179474 126168
rect 179510 116592 179566 116648
rect 179694 130464 179750 130520
rect 179602 113872 179658 113928
rect 121090 108296 121146 108352
rect 120998 107616 121054 107672
rect 120906 77560 120962 77616
rect 114006 10376 114062 10432
rect 123482 80144 123538 80200
rect 122378 79736 122434 79792
rect 122930 73888 122986 73944
rect 123298 78104 123354 78160
rect 124126 77968 124182 78024
rect 174910 80552 174966 80608
rect 174542 80280 174598 80336
rect 125828 79906 125884 79962
rect 126150 78240 126206 78296
rect 126058 77832 126114 77888
rect 127024 79736 127080 79792
rect 128036 79872 128092 79928
rect 126794 76472 126850 76528
rect 127070 75928 127126 75984
rect 128404 79872 128460 79928
rect 128680 79872 128736 79928
rect 129048 79872 129104 79928
rect 129508 79906 129564 79962
rect 128450 74160 128506 74216
rect 128726 78104 128782 78160
rect 129094 74432 129150 74488
rect 129462 79736 129518 79792
rect 129968 79872 130024 79928
rect 130290 79736 130346 79792
rect 129922 79600 129978 79656
rect 129646 77288 129702 77344
rect 130704 79872 130760 79928
rect 131164 79906 131220 79962
rect 131532 79872 131588 79928
rect 131256 79772 131258 79792
rect 131258 79772 131310 79792
rect 131310 79772 131312 79792
rect 131256 79736 131312 79772
rect 131716 79906 131772 79962
rect 130290 79600 130346 79656
rect 131210 79600 131266 79656
rect 131578 79600 131634 79656
rect 131394 77288 131450 77344
rect 131302 77152 131358 77208
rect 132176 79838 132232 79894
rect 132544 79872 132600 79928
rect 132820 79906 132876 79962
rect 132498 79600 132554 79656
rect 132590 78376 132646 78432
rect 132774 78104 132830 78160
rect 132682 76608 132738 76664
rect 131762 69536 131818 69592
rect 133648 79906 133704 79962
rect 134016 79906 134072 79962
rect 134200 79906 134256 79962
rect 134660 79906 134716 79962
rect 132866 77152 132922 77208
rect 133234 78240 133290 78296
rect 133602 78648 133658 78704
rect 133970 79600 134026 79656
rect 134338 79736 134394 79792
rect 134660 79736 134716 79792
rect 134246 78648 134302 78704
rect 134154 76744 134210 76800
rect 135120 79770 135176 79826
rect 135488 79906 135544 79962
rect 135948 79872 136004 79928
rect 135074 79600 135130 79656
rect 135258 77288 135314 77344
rect 135994 79600 136050 79656
rect 136592 79906 136648 79962
rect 136546 77832 136602 77888
rect 137052 79872 137108 79928
rect 136914 78648 136970 78704
rect 137972 79906 138028 79962
rect 137282 77832 137338 77888
rect 137282 77560 137338 77616
rect 137926 79772 137928 79792
rect 137928 79772 137980 79792
rect 137980 79772 137982 79792
rect 137926 79736 137982 79772
rect 138156 79872 138212 79928
rect 138018 78648 138074 78704
rect 138616 79872 138672 79928
rect 138800 79906 138856 79962
rect 138570 79736 138626 79792
rect 139352 79872 139408 79928
rect 138294 78240 138350 78296
rect 139168 79736 139224 79792
rect 139214 78240 139270 78296
rect 139536 79838 139592 79894
rect 140824 79906 140880 79962
rect 139398 79600 139454 79656
rect 140318 79620 140374 79656
rect 140318 79600 140320 79620
rect 140320 79600 140372 79620
rect 140372 79600 140374 79620
rect 140042 67496 140098 67552
rect 140502 77696 140558 77752
rect 140686 79600 140742 79656
rect 140778 78648 140834 78704
rect 140594 77424 140650 77480
rect 141468 79872 141524 79928
rect 141514 79736 141570 79792
rect 142020 79906 142076 79962
rect 142480 79906 142536 79962
rect 142756 79906 142812 79962
rect 142066 79736 142122 79792
rect 142066 79600 142122 79656
rect 142342 76744 142398 76800
rect 142710 79736 142766 79792
rect 142434 10920 142490 10976
rect 143400 79872 143456 79928
rect 143584 79872 143640 79928
rect 143768 79906 143824 79962
rect 144044 79872 144100 79928
rect 144320 79906 144376 79962
rect 143078 78104 143134 78160
rect 144872 79906 144928 79962
rect 144274 79736 144330 79792
rect 143354 78648 143410 78704
rect 143262 78240 143318 78296
rect 143538 79600 143594 79656
rect 143814 79600 143870 79656
rect 143906 78648 143962 78704
rect 144504 79736 144560 79792
rect 144872 79736 144928 79792
rect 144734 76880 144790 76936
rect 144642 74024 144698 74080
rect 145056 79906 145112 79962
rect 145102 78648 145158 78704
rect 144826 73616 144882 73672
rect 145792 79872 145848 79928
rect 145194 76336 145250 76392
rect 146022 79600 146078 79656
rect 146022 78648 146078 78704
rect 146114 78104 146170 78160
rect 146436 79872 146492 79928
rect 146712 79906 146768 79962
rect 147264 79872 147320 79928
rect 146758 79736 146814 79792
rect 146666 79600 146722 79656
rect 146298 76608 146354 76664
rect 146206 76472 146262 76528
rect 146850 77832 146906 77888
rect 147448 79906 147504 79962
rect 147494 79600 147550 79656
rect 147402 76608 147458 76664
rect 147586 76744 147642 76800
rect 147494 76472 147550 76528
rect 148276 79872 148332 79928
rect 148230 79736 148286 79792
rect 147862 76472 147918 76528
rect 148322 79600 148378 79656
rect 148920 79736 148976 79792
rect 149564 79872 149620 79928
rect 148782 78240 148838 78296
rect 148690 73888 148746 73944
rect 149242 77968 149298 78024
rect 148966 77832 149022 77888
rect 150116 79872 150172 79928
rect 149702 78104 149758 78160
rect 150668 79906 150724 79962
rect 150162 78104 150218 78160
rect 150254 77832 150310 77888
rect 150346 76608 150402 76664
rect 150898 79736 150954 79792
rect 151220 79872 151276 79928
rect 150990 78104 151046 78160
rect 151680 79906 151736 79962
rect 151634 78648 151690 78704
rect 151956 79872 152012 79928
rect 152324 79906 152380 79962
rect 152600 79906 152656 79962
rect 153428 79906 153484 79962
rect 151726 78376 151782 78432
rect 152094 79600 152150 79656
rect 152738 79736 152794 79792
rect 153980 79872 154036 79928
rect 154440 79872 154496 79928
rect 154624 79872 154680 79928
rect 154992 79906 155048 79962
rect 155176 79906 155232 79962
rect 155360 79872 155416 79928
rect 155636 79906 155692 79962
rect 155820 79906 155876 79962
rect 156096 79906 156152 79962
rect 153796 79736 153852 79792
rect 152186 77152 152242 77208
rect 152830 78648 152886 78704
rect 152738 78376 152794 78432
rect 152738 77424 152794 77480
rect 152922 77152 152978 77208
rect 153566 79600 153622 79656
rect 155130 79756 155186 79792
rect 155130 79736 155132 79756
rect 155132 79736 155184 79756
rect 155184 79736 155186 79756
rect 154762 79600 154818 79656
rect 154578 78104 154634 78160
rect 154302 77968 154358 78024
rect 155774 79736 155830 79792
rect 156556 79906 156612 79962
rect 157384 79906 157440 79962
rect 157108 79838 157164 79894
rect 155314 77832 155370 77888
rect 155682 77832 155738 77888
rect 156280 79736 156336 79792
rect 156142 79600 156198 79656
rect 155222 44784 155278 44840
rect 156326 78648 156382 78704
rect 156786 79736 156842 79792
rect 157430 79600 157486 79656
rect 157154 78648 157210 78704
rect 157062 77832 157118 77888
rect 156878 75384 156934 75440
rect 158120 79736 158176 79792
rect 158396 79906 158452 79962
rect 158672 79906 158728 79962
rect 158580 79736 158636 79792
rect 158718 79756 158774 79792
rect 158718 79736 158720 79756
rect 158720 79736 158772 79756
rect 158772 79736 158774 79756
rect 157890 78376 157946 78432
rect 158350 79600 158406 79656
rect 159224 79872 159280 79928
rect 159960 79872 160016 79928
rect 158994 77152 159050 77208
rect 158994 76472 159050 76528
rect 159362 79636 159364 79656
rect 159364 79636 159416 79656
rect 159416 79636 159418 79656
rect 159362 79600 159418 79636
rect 159362 78648 159418 78704
rect 159454 78104 159510 78160
rect 159362 75112 159418 75168
rect 160098 79736 160154 79792
rect 159730 78240 159786 78296
rect 160512 79872 160568 79928
rect 161064 79906 161120 79962
rect 161248 79872 161304 79928
rect 161524 79906 161580 79962
rect 161708 79906 161764 79962
rect 159914 75248 159970 75304
rect 160190 78376 160246 78432
rect 160834 75112 160890 75168
rect 161110 77424 161166 77480
rect 161202 77152 161258 77208
rect 161386 76336 161442 76392
rect 161570 75928 161626 75984
rect 161478 75248 161534 75304
rect 160742 50224 160798 50280
rect 158902 4800 158958 4856
rect 162720 79736 162776 79792
rect 162904 79872 162960 79928
rect 162398 79056 162454 79112
rect 162674 74976 162730 75032
rect 162950 79736 163006 79792
rect 164008 79872 164064 79928
rect 163042 79600 163098 79656
rect 162950 75656 163006 75712
rect 163686 79600 163742 79656
rect 163594 78376 163650 78432
rect 164100 79736 164156 79792
rect 164652 79838 164708 79894
rect 164238 79600 164294 79656
rect 164422 79636 164424 79656
rect 164424 79636 164476 79656
rect 164476 79636 164478 79656
rect 164422 79600 164478 79636
rect 164422 77560 164478 77616
rect 165572 79872 165628 79928
rect 165756 79906 165812 79962
rect 165480 79772 165482 79792
rect 165482 79772 165534 79792
rect 165534 79772 165536 79792
rect 164790 78648 164846 78704
rect 164974 79620 165030 79656
rect 164974 79600 164976 79620
rect 164976 79600 165028 79620
rect 165028 79600 165030 79620
rect 165480 79736 165536 79772
rect 164974 78648 165030 78704
rect 165158 78648 165214 78704
rect 165434 75928 165490 75984
rect 165618 79328 165674 79384
rect 165618 79056 165674 79112
rect 166400 79872 166456 79928
rect 166584 79872 166640 79928
rect 166078 79600 166134 79656
rect 166078 79328 166134 79384
rect 165986 79192 166042 79248
rect 165986 78512 166042 78568
rect 165986 77832 166042 77888
rect 165986 77560 166042 77616
rect 166262 79192 166318 79248
rect 166262 78104 166318 78160
rect 166952 79872 167008 79928
rect 166722 79600 166778 79656
rect 166630 77424 166686 77480
rect 166998 78648 167054 78704
rect 166906 77832 166962 77888
rect 166814 77288 166870 77344
rect 167182 79600 167238 79656
rect 167688 79872 167744 79928
rect 167182 78648 167238 78704
rect 167182 75928 167238 75984
rect 164882 3304 164938 3360
rect 167550 79328 167606 79384
rect 168148 79872 168204 79928
rect 168424 79906 168480 79962
rect 168010 79328 168066 79384
rect 168010 78648 168066 78704
rect 168010 78104 168066 78160
rect 168332 79736 168388 79792
rect 168976 79906 169032 79962
rect 168194 75928 168250 75984
rect 168654 79328 168710 79384
rect 169712 79872 169768 79928
rect 169896 79906 169952 79962
rect 170448 79906 170504 79962
rect 170816 79872 170872 79928
rect 168930 79328 168986 79384
rect 168746 78240 168802 78296
rect 169574 76472 169630 76528
rect 171184 79872 171240 79928
rect 169850 79328 169906 79384
rect 170402 79464 170458 79520
rect 170494 79328 170550 79384
rect 170586 78648 170642 78704
rect 170494 78240 170550 78296
rect 170310 77424 170366 77480
rect 170586 78104 170642 78160
rect 170954 75928 171010 75984
rect 171460 79906 171516 79962
rect 171736 79872 171792 79928
rect 171920 79872 171976 79928
rect 172196 79872 172252 79928
rect 171322 78648 171378 78704
rect 171230 77968 171286 78024
rect 171782 79364 171784 79384
rect 171784 79364 171836 79384
rect 171836 79364 171838 79384
rect 171782 79328 171838 79364
rect 172472 79872 172528 79928
rect 171966 78240 172022 78296
rect 172058 77832 172114 77888
rect 172426 79328 172482 79384
rect 172334 77152 172390 77208
rect 173208 79872 173264 79928
rect 172886 79192 172942 79248
rect 172794 77696 172850 77752
rect 173070 79600 173126 79656
rect 173760 79906 173816 79962
rect 173944 79906 174000 79962
rect 173070 79328 173126 79384
rect 173346 79328 173402 79384
rect 173346 79192 173402 79248
rect 173254 78784 173310 78840
rect 173438 79056 173494 79112
rect 173530 78920 173586 78976
rect 173162 76336 173218 76392
rect 173346 75656 173402 75712
rect 173622 3304 173678 3360
rect 174450 71032 174506 71088
rect 179418 78512 179474 78568
rect 176658 75520 176714 75576
rect 180890 122848 180946 122904
rect 180798 114688 180854 114744
rect 181074 128288 181130 128344
rect 180982 111968 181038 112024
rect 180062 80416 180118 80472
rect 182178 126928 182234 126984
rect 182270 124208 182326 124264
rect 182362 121488 182418 121544
rect 182178 109248 182234 109304
rect 182546 118768 182602 118824
rect 183006 129648 183062 129704
rect 182730 120128 182786 120184
rect 182638 117408 182694 117464
rect 182454 110608 182510 110664
rect 182270 107888 182326 107944
rect 182546 86128 182602 86184
rect 182730 84768 182786 84824
rect 182822 83408 182878 83464
rect 182822 82048 182878 82104
rect 182178 80688 182234 80744
rect 183282 106528 183338 106584
rect 183282 105168 183338 105224
rect 183282 103808 183338 103864
rect 183282 102448 183338 102504
rect 183282 101088 183338 101144
rect 183190 99728 183246 99784
rect 183190 98368 183246 98424
rect 183190 97008 183246 97064
rect 183190 95648 183246 95704
rect 183466 94288 183522 94344
rect 183466 92928 183522 92984
rect 183466 91568 183522 91624
rect 183466 90208 183522 90264
rect 183466 88848 183522 88904
rect 183466 87488 183522 87544
rect 184938 78240 184994 78296
rect 194598 74296 194654 74352
rect 193218 65456 193274 65512
rect 191838 40840 191894 40896
rect 193310 24384 193366 24440
rect 211158 77016 211214 77072
rect 212538 17312 212594 17368
rect 225142 3576 225198 3632
rect 230478 74160 230534 74216
rect 227718 58520 227774 58576
rect 227534 7792 227590 7848
rect 229374 13640 229430 13696
rect 247038 76880 247094 76936
rect 244278 74024 244334 74080
rect 242990 40704 243046 40760
rect 248418 19896 248474 19952
rect 246394 3440 246450 3496
rect 263598 57432 263654 57488
rect 266358 42064 266414 42120
rect 264978 13504 265034 13560
rect 282918 76744 282974 76800
rect 280710 12280 280766 12336
rect 279514 9152 279570 9208
rect 281906 6296 281962 6352
rect 284390 14728 284446 14784
rect 298098 73888 298154 73944
rect 299478 55800 299534 55856
rect 299570 25608 299626 25664
rect 301502 10648 301558 10704
rect 318798 76608 318854 76664
rect 316038 17176 316094 17232
rect 318062 12144 318118 12200
rect 317326 6160 317382 6216
rect 396906 80552 396962 80608
rect 397458 78648 397514 78704
rect 333978 62872 334034 62928
rect 336278 12008 336334 12064
rect 337014 10512 337070 10568
rect 351918 53352 351974 53408
rect 350538 21392 350594 21448
rect 354678 21256 354734 21312
rect 349250 15816 349306 15872
rect 369858 37848 369914 37904
rect 365810 14592 365866 14648
rect 372894 14456 372950 14512
rect 371238 13368 371294 13424
rect 402978 75384 403034 75440
rect 387798 44784 387854 44840
rect 386418 26832 386474 26888
rect 405738 29552 405794 29608
rect 407118 24248 407174 24304
rect 407210 24112 407266 24168
rect 423678 48864 423734 48920
rect 422298 22616 422354 22672
rect 462318 80008 462374 80064
rect 421378 4936 421434 4992
rect 424966 7656 425022 7712
rect 459558 75248 459614 75304
rect 440330 59880 440386 59936
rect 449898 57296 449954 57352
rect 442630 10376 442686 10432
rect 443366 10240 443422 10296
rect 458178 54440 458234 54496
rect 483018 77832 483074 77888
rect 456890 13232 456946 13288
rect 474094 11872 474150 11928
rect 478142 11736 478198 11792
rect 476946 9016 477002 9072
rect 496818 75112 496874 75168
rect 494058 57160 494114 57216
rect 495898 4800 495954 4856
rect 501786 3304 501842 3360
rect 511998 64096 512054 64152
rect 510618 40568 510674 40624
rect 513378 13096 513434 13152
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580262 644000 580318 644056
rect 579986 630808 580042 630864
rect 580170 577632 580226 577688
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580078 431568 580134 431624
rect 580078 418240 580134 418296
rect 580078 404912 580134 404968
rect 580078 378392 580134 378448
rect 579802 365064 579858 365120
rect 580078 351908 580080 351928
rect 580080 351908 580132 351928
rect 580132 351908 580134 351928
rect 580078 351872 580134 351908
rect 580078 312024 580134 312080
rect 580078 298696 580134 298752
rect 579802 272176 579858 272232
rect 579986 258848 580042 258904
rect 579986 245520 580042 245576
rect 580078 232328 580134 232384
rect 580170 219000 580226 219056
rect 580170 205692 580226 205728
rect 580170 205672 580172 205692
rect 580172 205672 580224 205692
rect 580224 205672 580226 205692
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 579986 152632 580042 152688
rect 580170 139304 580226 139360
rect 579802 125976 579858 126032
rect 580170 112784 580226 112840
rect 580170 99456 580226 99512
rect 579986 86128 580042 86184
rect 580722 617480 580778 617536
rect 580354 590960 580410 591016
rect 527178 77152 527234 77208
rect 514850 53216 514906 53272
rect 529938 69536 529994 69592
rect 528558 51720 528614 51776
rect 531318 39208 531374 39264
rect 531410 25472 531466 25528
rect 547878 62736 547934 62792
rect 546498 18536 546554 18592
rect 549258 46144 549314 46200
rect 549074 7520 549130 7576
rect 580538 564304 580594 564360
rect 580446 537784 580502 537840
rect 580630 484608 580686 484664
rect 580814 511264 580870 511320
rect 580906 325216 580962 325272
rect 580722 192480 580778 192536
rect 565818 76472 565874 76528
rect 578238 73752 578294 73808
rect 567566 12960 567622 13016
rect 575478 53080 575534 53136
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 19760 580226 19816
rect 577410 8880 577466 8936
rect 580262 6568 580318 6624
rect 583390 11600 583446 11656
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697234 584960 697324
rect 567150 697174 584960 697234
rect 396574 696900 396580 696964
rect 396644 696962 396650 696964
rect 567150 696962 567210 697174
rect 583520 697084 584960 697174
rect 396644 696902 567210 696962
rect 396644 696900 396650 696902
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580257 644058 580323 644061
rect 583520 644058 584960 644148
rect 580257 644056 584960 644058
rect 580257 644000 580262 644056
rect 580318 644000 584960 644056
rect 580257 643998 584960 644000
rect 580257 643995 580323 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3325 632090 3391 632093
rect -960 632088 3391 632090
rect -960 632032 3330 632088
rect 3386 632032 3391 632088
rect -960 632030 3391 632032
rect -960 631940 480 632030
rect 3325 632027 3391 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3693 619170 3759 619173
rect -960 619168 3759 619170
rect -960 619112 3698 619168
rect 3754 619112 3759 619168
rect -960 619110 3759 619112
rect -960 619020 480 619110
rect 3693 619107 3759 619110
rect 580717 617538 580783 617541
rect 583520 617538 584960 617628
rect 580717 617536 584960 617538
rect 580717 617480 580722 617536
rect 580778 617480 584960 617536
rect 580717 617478 584960 617480
rect 580717 617475 580783 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3601 606114 3667 606117
rect -960 606112 3667 606114
rect -960 606056 3606 606112
rect 3662 606056 3667 606112
rect -960 606054 3667 606056
rect -960 605964 480 606054
rect 3601 606051 3667 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580349 591018 580415 591021
rect 583520 591018 584960 591108
rect 580349 591016 584960 591018
rect 580349 590960 580354 591016
rect 580410 590960 584960 591016
rect 580349 590958 584960 590960
rect 580349 590955 580415 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3877 566946 3943 566949
rect -960 566944 3943 566946
rect -960 566888 3882 566944
rect 3938 566888 3943 566944
rect -960 566886 3943 566888
rect -960 566796 480 566886
rect 3877 566883 3943 566886
rect 580533 564362 580599 564365
rect 583520 564362 584960 564452
rect 580533 564360 584960 564362
rect 580533 564304 580538 564360
rect 580594 564304 584960 564360
rect 580533 564302 584960 564304
rect 580533 564299 580599 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3785 553890 3851 553893
rect -960 553888 3851 553890
rect -960 553832 3790 553888
rect 3846 553832 3851 553888
rect -960 553830 3851 553832
rect -960 553740 480 553830
rect 3785 553827 3851 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580441 537842 580507 537845
rect 583520 537842 584960 537932
rect 580441 537840 584960 537842
rect 580441 537784 580446 537840
rect 580502 537784 584960 537840
rect 580441 537782 584960 537784
rect 580441 537779 580507 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 580809 511322 580875 511325
rect 583520 511322 584960 511412
rect 580809 511320 584960 511322
rect 580809 511264 580814 511320
rect 580870 511264 584960 511320
rect 580809 511262 584960 511264
rect 580809 511259 580875 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3233 501802 3299 501805
rect -960 501800 3299 501802
rect -960 501744 3238 501800
rect 3294 501744 3299 501800
rect -960 501742 3299 501744
rect -960 501652 480 501742
rect 3233 501739 3299 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580625 484666 580691 484669
rect 583520 484666 584960 484756
rect 580625 484664 584960 484666
rect 580625 484608 580630 484664
rect 580686 484608 584960 484664
rect 580625 484606 584960 484608
rect 580625 484603 580691 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580073 431626 580139 431629
rect 583520 431626 584960 431716
rect 580073 431624 584960 431626
rect 580073 431568 580078 431624
rect 580134 431568 584960 431624
rect 580073 431566 584960 431568
rect 580073 431563 580139 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 2957 423602 3023 423605
rect -960 423600 3023 423602
rect -960 423544 2962 423600
rect 3018 423544 3023 423600
rect -960 423542 3023 423544
rect -960 423452 480 423542
rect 2957 423539 3023 423542
rect 580073 418298 580139 418301
rect 583520 418298 584960 418388
rect 580073 418296 584960 418298
rect 580073 418240 580078 418296
rect 580134 418240 584960 418296
rect 580073 418238 584960 418240
rect 580073 418235 580139 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580073 404970 580139 404973
rect 583520 404970 584960 405060
rect 580073 404968 584960 404970
rect 580073 404912 580078 404968
rect 580134 404912 584960 404968
rect 580073 404910 584960 404912
rect 580073 404907 580139 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580073 378450 580139 378453
rect 583520 378450 584960 378540
rect 580073 378448 584960 378450
rect 580073 378392 580078 378448
rect 580134 378392 584960 378448
rect 580073 378390 584960 378392
rect 580073 378387 580139 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 579797 365122 579863 365125
rect 583520 365122 584960 365212
rect 579797 365120 584960 365122
rect 579797 365064 579802 365120
rect 579858 365064 584960 365120
rect 579797 365062 584960 365064
rect 579797 365059 579863 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580073 351930 580139 351933
rect 583520 351930 584960 352020
rect 580073 351928 584960 351930
rect 580073 351872 580078 351928
rect 580134 351872 584960 351928
rect 580073 351870 584960 351872
rect 580073 351867 580139 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580901 325274 580967 325277
rect 583520 325274 584960 325364
rect 580901 325272 584960 325274
rect 580901 325216 580906 325272
rect 580962 325216 584960 325272
rect 580901 325214 584960 325216
rect 580901 325211 580967 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3141 319290 3207 319293
rect -960 319288 3207 319290
rect -960 319232 3146 319288
rect 3202 319232 3207 319288
rect -960 319230 3207 319232
rect -960 319140 480 319230
rect 3141 319227 3207 319230
rect 580073 312082 580139 312085
rect 583520 312082 584960 312172
rect 580073 312080 584960 312082
rect 580073 312024 580078 312080
rect 580134 312024 584960 312080
rect 580073 312022 584960 312024
rect 580073 312019 580139 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 4061 306234 4127 306237
rect -960 306232 4127 306234
rect -960 306176 4066 306232
rect 4122 306176 4127 306232
rect -960 306174 4127 306176
rect -960 306084 480 306174
rect 4061 306171 4127 306174
rect 580073 298754 580139 298757
rect 583520 298754 584960 298844
rect 580073 298752 584960 298754
rect 580073 298696 580078 298752
rect 580134 298696 584960 298752
rect 580073 298694 584960 298696
rect 580073 298691 580139 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3969 293178 4035 293181
rect -960 293176 4035 293178
rect -960 293120 3974 293176
rect 4030 293120 4035 293176
rect -960 293118 4035 293120
rect -960 293028 480 293118
rect 3969 293115 4035 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579797 272234 579863 272237
rect 583520 272234 584960 272324
rect 579797 272232 584960 272234
rect 579797 272176 579802 272232
rect 579858 272176 584960 272232
rect 579797 272174 584960 272176
rect 579797 272171 579863 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3233 267202 3299 267205
rect -960 267200 3299 267202
rect -960 267144 3238 267200
rect 3294 267144 3299 267200
rect -960 267142 3299 267144
rect -960 267052 480 267142
rect 3233 267139 3299 267142
rect 579981 258906 580047 258909
rect 583520 258906 584960 258996
rect 579981 258904 584960 258906
rect 579981 258848 579986 258904
rect 580042 258848 584960 258904
rect 579981 258846 584960 258848
rect 579981 258843 580047 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3325 254146 3391 254149
rect -960 254144 3391 254146
rect -960 254088 3330 254144
rect 3386 254088 3391 254144
rect -960 254086 3391 254088
rect -960 253996 480 254086
rect 3325 254083 3391 254086
rect 579981 245578 580047 245581
rect 583520 245578 584960 245668
rect 579981 245576 584960 245578
rect 579981 245520 579986 245576
rect 580042 245520 584960 245576
rect 579981 245518 584960 245520
rect 579981 245515 580047 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 580073 232386 580139 232389
rect 583520 232386 584960 232476
rect 580073 232384 584960 232386
rect 580073 232328 580078 232384
rect 580134 232328 584960 232384
rect 580073 232326 584960 232328
rect 580073 232323 580139 232326
rect 583520 232236 584960 232326
rect -960 228034 480 228124
rect 3049 228034 3115 228037
rect -960 228032 3115 228034
rect -960 227976 3054 228032
rect 3110 227976 3115 228032
rect -960 227974 3115 227976
rect -960 227884 480 227974
rect 3049 227971 3115 227974
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3693 201922 3759 201925
rect -960 201920 3759 201922
rect -960 201864 3698 201920
rect 3754 201864 3759 201920
rect -960 201862 3759 201864
rect -960 201772 480 201862
rect 3693 201859 3759 201862
rect 143533 200698 143599 200701
rect 144678 200698 144684 200700
rect 143533 200696 144684 200698
rect 143533 200640 143538 200696
rect 143594 200640 144684 200696
rect 143533 200638 144684 200640
rect 143533 200635 143599 200638
rect 144678 200636 144684 200638
rect 144748 200636 144754 200700
rect 147622 199276 147628 199340
rect 147692 199338 147698 199340
rect 163497 199338 163563 199341
rect 147692 199336 163563 199338
rect 147692 199280 163502 199336
rect 163558 199280 163563 199336
rect 147692 199278 163563 199280
rect 147692 199276 147698 199278
rect 163497 199275 163563 199278
rect 147489 196482 147555 196485
rect 147622 196482 147628 196484
rect 147489 196480 147628 196482
rect 147489 196424 147494 196480
rect 147550 196424 147628 196480
rect 147489 196422 147628 196424
rect 147489 196419 147555 196422
rect 147622 196420 147628 196422
rect 147692 196420 147698 196484
rect 153285 196210 153351 196213
rect 166073 196210 166139 196213
rect 153285 196208 166139 196210
rect 153285 196152 153290 196208
rect 153346 196152 166078 196208
rect 166134 196152 166139 196208
rect 153285 196150 166139 196152
rect 153285 196147 153351 196150
rect 166073 196147 166139 196150
rect 151302 196012 151308 196076
rect 151372 196074 151378 196076
rect 166165 196074 166231 196077
rect 151372 196072 166231 196074
rect 151372 196016 166170 196072
rect 166226 196016 166231 196072
rect 151372 196014 166231 196016
rect 151372 196012 151378 196014
rect 166165 196011 166231 196014
rect 139393 195938 139459 195941
rect 142337 195938 142403 195941
rect 153193 195938 153259 195941
rect 139393 195936 142403 195938
rect 139393 195880 139398 195936
rect 139454 195880 142342 195936
rect 142398 195880 142403 195936
rect 139393 195878 142403 195880
rect 139393 195875 139459 195878
rect 142337 195875 142403 195878
rect 151126 195936 153259 195938
rect 151126 195880 153198 195936
rect 153254 195880 153259 195936
rect 151126 195878 153259 195880
rect 138105 195802 138171 195805
rect 140773 195802 140839 195805
rect 138105 195800 140839 195802
rect 138105 195744 138110 195800
rect 138166 195744 140778 195800
rect 140834 195744 140839 195800
rect 138105 195742 140839 195744
rect 138105 195739 138171 195742
rect 140773 195739 140839 195742
rect 151126 195696 151186 195878
rect 153193 195875 153259 195878
rect 153929 195938 153995 195941
rect 155953 195938 156019 195941
rect 158253 195938 158319 195941
rect 153929 195936 156019 195938
rect 153929 195880 153934 195936
rect 153990 195880 155958 195936
rect 156014 195880 156019 195936
rect 153929 195878 156019 195880
rect 153929 195875 153995 195878
rect 155953 195875 156019 195878
rect 156278 195936 158319 195938
rect 156278 195880 158258 195936
rect 158314 195880 158319 195936
rect 156278 195878 158319 195880
rect 156278 195802 156338 195878
rect 158253 195875 158319 195878
rect 158897 195938 158963 195941
rect 161381 195938 161447 195941
rect 158897 195936 161447 195938
rect 158897 195880 158902 195936
rect 158958 195880 161386 195936
rect 161442 195880 161447 195936
rect 158897 195878 161447 195880
rect 158897 195875 158963 195878
rect 161381 195875 161447 195878
rect 159817 195802 159883 195805
rect 144678 195604 144684 195668
rect 144748 195604 144754 195668
rect 149830 195604 149836 195668
rect 149900 195666 149906 195668
rect 150341 195666 150407 195669
rect 149900 195664 150407 195666
rect 149900 195608 150346 195664
rect 150402 195608 150407 195664
rect 150604 195636 151186 195696
rect 155358 195742 156338 195802
rect 157750 195800 159883 195802
rect 157750 195744 159822 195800
rect 159878 195744 159883 195800
rect 157750 195742 159883 195744
rect 155358 195666 155418 195742
rect 157750 195696 157810 195742
rect 159817 195739 159883 195742
rect 157228 195636 157810 195696
rect 149900 195606 150407 195608
rect 149900 195604 149906 195606
rect 144686 195410 144746 195604
rect 150341 195603 150407 195606
rect 153929 194714 153995 194717
rect 155217 194714 155283 194717
rect 153929 194712 155283 194714
rect 153929 194656 153934 194712
rect 153990 194656 155222 194712
rect 155278 194656 155283 194712
rect 153929 194654 155283 194656
rect 153929 194651 153995 194654
rect 155217 194651 155283 194654
rect 151629 193626 151695 193629
rect 153285 193626 153351 193629
rect 151629 193624 153351 193626
rect 151629 193568 151634 193624
rect 151690 193568 153290 193624
rect 153346 193568 153351 193624
rect 151629 193566 153351 193568
rect 151629 193563 151695 193566
rect 153285 193563 153351 193566
rect 580717 192538 580783 192541
rect 583520 192538 584960 192628
rect 580717 192536 584960 192538
rect 580717 192480 580722 192536
rect 580778 192480 584960 192536
rect 580717 192478 584960 192480
rect 580717 192475 580783 192478
rect 583520 192388 584960 192478
rect 143574 191744 143580 191808
rect 143644 191806 143650 191808
rect 143644 191746 143796 191806
rect 143644 191744 143650 191746
rect 143536 191336 144164 191396
rect 141734 191252 141740 191316
rect 141804 191314 141810 191316
rect 143536 191314 143596 191336
rect 151302 191316 151308 191318
rect 141804 191254 143596 191314
rect 151156 191256 151308 191316
rect 151302 191254 151308 191256
rect 151372 191254 151378 191318
rect 141804 191252 141810 191254
rect 141918 190572 141924 190636
rect 141988 190634 141994 190636
rect 144134 190634 144194 191226
rect 141988 190574 144194 190634
rect 149789 190636 149855 190637
rect 149789 190632 149836 190636
rect 149900 190634 149906 190636
rect 149789 190576 149794 190632
rect 141988 190572 141994 190574
rect 149789 190572 149836 190576
rect 149900 190574 149946 190634
rect 149900 190572 149906 190574
rect 149789 190571 149855 190572
rect -960 188866 480 188956
rect 2957 188866 3023 188869
rect -960 188864 3023 188866
rect -960 188808 2962 188864
rect 3018 188808 3023 188864
rect -960 188806 3023 188808
rect -960 188716 480 188806
rect 2957 188803 3023 188806
rect 140630 186900 140636 186964
rect 140700 186962 140706 186964
rect 144637 186962 144703 186965
rect 140700 186960 144703 186962
rect 140700 186904 144642 186960
rect 144698 186904 144703 186960
rect 140700 186902 144703 186904
rect 140700 186900 140706 186902
rect 144637 186899 144703 186902
rect 146109 180708 146175 180709
rect 146109 180704 146156 180708
rect 146220 180706 146226 180708
rect 146109 180648 146114 180704
rect 146109 180644 146156 180648
rect 146220 180646 146266 180706
rect 146220 180644 146226 180646
rect 146109 180643 146175 180644
rect 140446 179148 140452 179212
rect 140516 179210 140522 179212
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 140516 179150 148058 179210
rect 140516 179148 140522 179150
rect 147998 179077 148058 179150
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 147998 179072 148107 179077
rect 147998 179016 148046 179072
rect 148102 179016 148107 179072
rect 583520 179060 584960 179150
rect 147998 179014 148107 179016
rect 148041 179011 148107 179014
rect 142661 178804 142727 178805
rect 142654 178740 142660 178804
rect 142724 178802 142730 178804
rect 142724 178742 142816 178802
rect 142724 178740 142730 178742
rect 142661 178739 142727 178740
rect 142061 176762 142127 176765
rect 142654 176762 142660 176764
rect 142061 176760 142660 176762
rect 142061 176704 142066 176760
rect 142122 176704 142660 176760
rect 142061 176702 142660 176704
rect 142061 176699 142127 176702
rect 142654 176700 142660 176702
rect 142724 176700 142730 176764
rect -960 175946 480 176036
rect 3325 175946 3391 175949
rect -960 175944 3391 175946
rect -960 175888 3330 175944
rect 3386 175888 3391 175944
rect -960 175886 3391 175888
rect -960 175796 480 175886
rect 3325 175883 3391 175886
rect 144177 174586 144243 174589
rect 156045 174586 156111 174589
rect 144177 174584 156111 174586
rect 144177 174528 144182 174584
rect 144238 174528 156050 174584
rect 156106 174528 156111 174584
rect 144177 174526 156111 174528
rect 144177 174523 144243 174526
rect 156045 174523 156111 174526
rect 135253 174042 135319 174045
rect 137829 174042 137895 174045
rect 135253 174040 137895 174042
rect 135253 173984 135258 174040
rect 135314 173984 137834 174040
rect 137890 173984 137895 174040
rect 135253 173982 137895 173984
rect 135253 173979 135319 173982
rect 137829 173979 137895 173982
rect 142470 173844 142476 173908
rect 142540 173906 142546 173908
rect 145649 173906 145715 173909
rect 142540 173904 145715 173906
rect 142540 173848 145654 173904
rect 145710 173848 145715 173904
rect 142540 173846 145715 173848
rect 142540 173844 142546 173846
rect 145649 173843 145715 173846
rect 142286 173708 142292 173772
rect 142356 173770 142362 173772
rect 142613 173770 142679 173773
rect 142356 173768 142679 173770
rect 142356 173712 142618 173768
rect 142674 173712 142679 173768
rect 142356 173710 142679 173712
rect 142356 173708 142362 173710
rect 142613 173707 142679 173710
rect 144126 173708 144132 173772
rect 144196 173770 144202 173772
rect 148685 173770 148751 173773
rect 144196 173768 148751 173770
rect 144196 173712 148690 173768
rect 148746 173712 148751 173768
rect 144196 173710 148751 173712
rect 144196 173708 144202 173710
rect 148685 173707 148751 173710
rect 142654 173572 142660 173636
rect 142724 173634 142730 173636
rect 146753 173634 146819 173637
rect 142724 173632 146819 173634
rect 142724 173576 146758 173632
rect 146814 173576 146819 173632
rect 142724 173574 146819 173576
rect 142724 173572 142730 173574
rect 146753 173571 146819 173574
rect 142102 171260 142108 171324
rect 142172 171260 142178 171324
rect 142110 171189 142170 171260
rect 142061 171186 142170 171189
rect 142016 171184 142170 171186
rect 142016 171128 142066 171184
rect 142122 171128 142170 171184
rect 142016 171126 142170 171128
rect 142061 171123 142127 171126
rect 142061 171050 142127 171053
rect 142016 171048 142170 171050
rect 142016 170992 142066 171048
rect 142122 170992 142170 171048
rect 142016 170990 142170 170992
rect 142061 170987 142170 170990
rect 142110 170916 142170 170987
rect 142102 170852 142108 170916
rect 142172 170852 142178 170916
rect 141734 166364 141740 166428
rect 141804 166426 141810 166428
rect 164325 166426 164391 166429
rect 141804 166424 164391 166426
rect 141804 166368 164330 166424
rect 164386 166368 164391 166424
rect 141804 166366 164391 166368
rect 141804 166364 141810 166366
rect 164325 166363 164391 166366
rect 141918 166228 141924 166292
rect 141988 166290 141994 166292
rect 166993 166290 167059 166293
rect 141988 166288 167059 166290
rect 141988 166232 166998 166288
rect 167054 166232 167059 166288
rect 141988 166230 167059 166232
rect 141988 166228 141994 166230
rect 166993 166227 167059 166230
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 142061 161532 142127 161533
rect 142061 161530 142108 161532
rect 142016 161528 142108 161530
rect 142172 161530 142178 161532
rect 142016 161472 142066 161528
rect 142016 161470 142108 161472
rect 142061 161468 142108 161470
rect 142172 161470 142254 161530
rect 142172 161468 142178 161470
rect 142061 161467 142127 161468
rect 579981 152690 580047 152693
rect 583520 152690 584960 152780
rect 579981 152688 584960 152690
rect 579981 152632 579986 152688
rect 580042 152632 584960 152688
rect 579981 152630 584960 152632
rect 579981 152627 580047 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 142470 143380 142476 143444
rect 142540 143442 142546 143444
rect 146477 143442 146543 143445
rect 142540 143440 146543 143442
rect 142540 143384 146482 143440
rect 146538 143384 146543 143440
rect 142540 143382 146543 143384
rect 142540 143380 142546 143382
rect 146477 143379 146543 143382
rect 142654 143244 142660 143308
rect 142724 143306 142730 143308
rect 148041 143306 148107 143309
rect 142724 143304 148107 143306
rect 142724 143248 148046 143304
rect 148102 143248 148107 143304
rect 142724 143246 148107 143248
rect 142724 143244 142730 143246
rect 148041 143243 148107 143246
rect 140446 143108 140452 143172
rect 140516 143170 140522 143172
rect 149605 143170 149671 143173
rect 140516 143168 149671 143170
rect 140516 143112 149610 143168
rect 149666 143112 149671 143168
rect 140516 143110 149671 143112
rect 140516 143108 140522 143110
rect 149605 143107 149671 143110
rect 144126 142972 144132 143036
rect 144196 143034 144202 143036
rect 151169 143034 151235 143037
rect 144196 143032 151235 143034
rect 144196 142976 151174 143032
rect 151230 142976 151235 143032
rect 144196 142974 151235 142976
rect 144196 142972 144202 142974
rect 151169 142971 151235 142974
rect 151353 143034 151419 143037
rect 160553 143034 160619 143037
rect 151353 143032 160619 143034
rect 151353 142976 151358 143032
rect 151414 142976 160558 143032
rect 160614 142976 160619 143032
rect 151353 142974 160619 142976
rect 151353 142971 151419 142974
rect 160553 142971 160619 142974
rect 146150 142836 146156 142900
rect 146220 142898 146226 142900
rect 171501 142898 171567 142901
rect 146220 142896 171567 142898
rect 146220 142840 171506 142896
rect 171562 142840 171567 142896
rect 146220 142838 171567 142840
rect 146220 142836 146226 142838
rect 171501 142835 171567 142838
rect 140630 142700 140636 142764
rect 140700 142762 140706 142764
rect 173065 142762 173131 142765
rect 140700 142760 173131 142762
rect 140700 142704 173070 142760
rect 173126 142704 173131 142760
rect 140700 142702 173131 142704
rect 140700 142700 140706 142702
rect 173065 142699 173131 142702
rect 143574 142564 143580 142628
rect 143644 142626 143650 142628
rect 151353 142626 151419 142629
rect 143644 142624 151419 142626
rect 143644 142568 151358 142624
rect 151414 142568 151419 142624
rect 143644 142566 151419 142568
rect 143644 142564 143650 142566
rect 151353 142563 151419 142566
rect 142102 142428 142108 142492
rect 142172 142490 142178 142492
rect 143533 142490 143599 142493
rect 142172 142488 143599 142490
rect 142172 142432 143538 142488
rect 143594 142432 143599 142488
rect 142172 142430 143599 142432
rect 142172 142428 142178 142430
rect 143533 142427 143599 142430
rect 142061 142218 142127 142221
rect 142286 142218 142292 142220
rect 142061 142216 142292 142218
rect 142061 142160 142066 142216
rect 142122 142160 142292 142216
rect 142061 142158 142292 142160
rect 142061 142155 142127 142158
rect 142286 142156 142292 142158
rect 142356 142156 142362 142220
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 117313 137594 117379 137597
rect 117313 137592 120060 137594
rect 117313 137536 117318 137592
rect 117374 137536 120060 137592
rect 117313 137534 120060 137536
rect 117313 137531 117379 137534
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 117313 136098 117379 136101
rect 117313 136096 120060 136098
rect 117313 136040 117318 136096
rect 117374 136040 120060 136096
rect 117313 136038 120060 136040
rect 117313 136035 117379 136038
rect 117313 134602 117379 134605
rect 117313 134600 120060 134602
rect 117313 134544 117318 134600
rect 117374 134544 120060 134600
rect 117313 134542 120060 134544
rect 117313 134539 117379 134542
rect 117405 133106 117471 133109
rect 117405 133104 120060 133106
rect 117405 133048 117410 133104
rect 117466 133048 120060 133104
rect 117405 133046 120060 133048
rect 117405 133043 117471 133046
rect 117313 131610 117379 131613
rect 117313 131608 120060 131610
rect 117313 131552 117318 131608
rect 117374 131552 120060 131608
rect 117313 131550 120060 131552
rect 117313 131547 117379 131550
rect 179646 130525 179706 131036
rect 179646 130520 179755 130525
rect 179646 130464 179694 130520
rect 179750 130464 179755 130520
rect 179646 130462 179755 130464
rect 179689 130459 179755 130462
rect 117313 130114 117379 130117
rect 117313 130112 120060 130114
rect 117313 130056 117318 130112
rect 117374 130056 120060 130112
rect 117313 130054 120060 130056
rect 117313 130051 117379 130054
rect 183001 129706 183067 129709
rect 179860 129704 183067 129706
rect 179860 129648 183006 129704
rect 183062 129648 183067 129704
rect 179860 129646 183067 129648
rect 183001 129643 183067 129646
rect 117313 128618 117379 128621
rect 117313 128616 120060 128618
rect 117313 128560 117318 128616
rect 117374 128560 120060 128616
rect 117313 128558 120060 128560
rect 117313 128555 117379 128558
rect 181069 128346 181135 128349
rect 179860 128344 181135 128346
rect 179860 128288 181074 128344
rect 181130 128288 181135 128344
rect 179860 128286 181135 128288
rect 181069 128283 181135 128286
rect 117313 127122 117379 127125
rect 117313 127120 120060 127122
rect 117313 127064 117318 127120
rect 117374 127064 120060 127120
rect 117313 127062 120060 127064
rect 117313 127059 117379 127062
rect 182173 126986 182239 126989
rect 179860 126984 182239 126986
rect 179860 126928 182178 126984
rect 182234 126928 182239 126984
rect 179860 126926 182239 126928
rect 182173 126923 182239 126926
rect 179413 126170 179479 126173
rect 179413 126168 179522 126170
rect 179413 126112 179418 126168
rect 179474 126112 179522 126168
rect 179413 126107 179522 126112
rect 117313 125626 117379 125629
rect 117313 125624 120060 125626
rect 117313 125568 117318 125624
rect 117374 125568 120060 125624
rect 179462 125596 179522 126107
rect 579797 126034 579863 126037
rect 583520 126034 584960 126124
rect 579797 126032 584960 126034
rect 579797 125976 579802 126032
rect 579858 125976 584960 126032
rect 579797 125974 584960 125976
rect 579797 125971 579863 125974
rect 583520 125884 584960 125974
rect 117313 125566 120060 125568
rect 117313 125563 117379 125566
rect 182265 124266 182331 124269
rect 179860 124264 182331 124266
rect 179860 124208 182270 124264
rect 182326 124208 182331 124264
rect 179860 124206 182331 124208
rect 182265 124203 182331 124206
rect 117313 124130 117379 124133
rect 117313 124128 120060 124130
rect 117313 124072 117318 124128
rect 117374 124072 120060 124128
rect 117313 124070 120060 124072
rect 117313 124067 117379 124070
rect -960 123572 480 123812
rect 180885 122906 180951 122909
rect 179860 122904 180951 122906
rect 179860 122848 180890 122904
rect 180946 122848 180951 122904
rect 179860 122846 180951 122848
rect 180885 122843 180951 122846
rect 117313 122634 117379 122637
rect 117313 122632 120060 122634
rect 117313 122576 117318 122632
rect 117374 122576 120060 122632
rect 117313 122574 120060 122576
rect 117313 122571 117379 122574
rect 182357 121546 182423 121549
rect 179860 121544 182423 121546
rect 179860 121488 182362 121544
rect 182418 121488 182423 121544
rect 179860 121486 182423 121488
rect 182357 121483 182423 121486
rect 117313 121138 117379 121141
rect 117313 121136 120060 121138
rect 117313 121080 117318 121136
rect 117374 121080 120060 121136
rect 117313 121078 120060 121080
rect 117313 121075 117379 121078
rect 182725 120186 182791 120189
rect 179860 120184 182791 120186
rect 179860 120128 182730 120184
rect 182786 120128 182791 120184
rect 179860 120126 182791 120128
rect 182725 120123 182791 120126
rect 117313 119642 117379 119645
rect 117313 119640 120060 119642
rect 117313 119584 117318 119640
rect 117374 119584 120060 119640
rect 117313 119582 120060 119584
rect 117313 119579 117379 119582
rect 182541 118826 182607 118829
rect 179860 118824 182607 118826
rect 179860 118768 182546 118824
rect 182602 118768 182607 118824
rect 179860 118766 182607 118768
rect 182541 118763 182607 118766
rect 117313 118146 117379 118149
rect 117313 118144 120060 118146
rect 117313 118088 117318 118144
rect 117374 118088 120060 118144
rect 117313 118086 120060 118088
rect 117313 118083 117379 118086
rect 182633 117466 182699 117469
rect 179860 117464 182699 117466
rect 179860 117408 182638 117464
rect 182694 117408 182699 117464
rect 179860 117406 182699 117408
rect 182633 117403 182699 117406
rect 117313 116650 117379 116653
rect 179505 116650 179571 116653
rect 117313 116648 120060 116650
rect 117313 116592 117318 116648
rect 117374 116592 120060 116648
rect 117313 116590 120060 116592
rect 179462 116648 179571 116650
rect 179462 116592 179510 116648
rect 179566 116592 179571 116648
rect 117313 116587 117379 116590
rect 179462 116587 179571 116592
rect 179462 116076 179522 116587
rect 117313 115154 117379 115157
rect 117313 115152 120060 115154
rect 117313 115096 117318 115152
rect 117374 115096 120060 115152
rect 117313 115094 120060 115096
rect 117313 115091 117379 115094
rect 180793 114746 180859 114749
rect 179860 114744 180859 114746
rect 179860 114688 180798 114744
rect 180854 114688 180859 114744
rect 179860 114686 180859 114688
rect 180793 114683 180859 114686
rect 179597 113930 179663 113933
rect 179597 113928 179706 113930
rect 179597 113872 179602 113928
rect 179658 113872 179706 113928
rect 179597 113867 179706 113872
rect 117313 113658 117379 113661
rect 117313 113656 120060 113658
rect 117313 113600 117318 113656
rect 117374 113600 120060 113656
rect 117313 113598 120060 113600
rect 117313 113595 117379 113598
rect 179646 113356 179706 113867
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect 117313 112162 117379 112165
rect 117313 112160 120060 112162
rect 117313 112104 117318 112160
rect 117374 112104 120060 112160
rect 117313 112102 120060 112104
rect 117313 112099 117379 112102
rect 180977 112026 181043 112029
rect 179860 112024 181043 112026
rect 179860 111968 180982 112024
rect 181038 111968 181043 112024
rect 179860 111966 181043 111968
rect 180977 111963 181043 111966
rect -960 110666 480 110756
rect 2957 110666 3023 110669
rect -960 110664 3023 110666
rect -960 110608 2962 110664
rect 3018 110608 3023 110664
rect -960 110606 3023 110608
rect -960 110516 480 110606
rect 2957 110603 3023 110606
rect 117313 110666 117379 110669
rect 182449 110666 182515 110669
rect 117313 110664 120060 110666
rect 117313 110608 117318 110664
rect 117374 110608 120060 110664
rect 117313 110606 120060 110608
rect 179860 110664 182515 110666
rect 179860 110608 182454 110664
rect 182510 110608 182515 110664
rect 179860 110606 182515 110608
rect 117313 110603 117379 110606
rect 182449 110603 182515 110606
rect 182173 109306 182239 109309
rect 179860 109304 182239 109306
rect 179860 109248 182178 109304
rect 182234 109248 182239 109304
rect 179860 109246 182239 109248
rect 182173 109243 182239 109246
rect 118601 109170 118667 109173
rect 118601 109168 120060 109170
rect 118601 109112 118606 109168
rect 118662 109112 120060 109168
rect 118601 109110 120060 109112
rect 118601 109107 118667 109110
rect 120625 108354 120691 108357
rect 121085 108354 121151 108357
rect 120625 108352 121151 108354
rect 120625 108296 120630 108352
rect 120686 108296 121090 108352
rect 121146 108296 121151 108352
rect 120625 108294 121151 108296
rect 120625 108291 120691 108294
rect 121085 108291 121151 108294
rect 182265 107946 182331 107949
rect 179860 107944 182331 107946
rect 179860 107888 182270 107944
rect 182326 107888 182331 107944
rect 179860 107886 182331 107888
rect 182265 107883 182331 107886
rect 120993 107674 121059 107677
rect 120612 107672 121059 107674
rect 120612 107616 120998 107672
rect 121054 107616 121059 107672
rect 120612 107614 121059 107616
rect 120993 107611 121059 107614
rect 183277 106586 183343 106589
rect 179860 106584 183343 106586
rect 179860 106528 183282 106584
rect 183338 106528 183343 106584
rect 179860 106526 183343 106528
rect 183277 106523 183343 106526
rect 118969 106178 119035 106181
rect 118969 106176 120060 106178
rect 118969 106120 118974 106176
rect 119030 106120 120060 106176
rect 118969 106118 120060 106120
rect 118969 106115 119035 106118
rect 183277 105226 183343 105229
rect 179860 105224 183343 105226
rect 179860 105168 183282 105224
rect 183338 105168 183343 105224
rect 179860 105166 183343 105168
rect 183277 105163 183343 105166
rect 118877 104682 118943 104685
rect 118877 104680 120060 104682
rect 118877 104624 118882 104680
rect 118938 104624 120060 104680
rect 118877 104622 120060 104624
rect 118877 104619 118943 104622
rect 183277 103866 183343 103869
rect 179860 103864 183343 103866
rect 179860 103808 183282 103864
rect 183338 103808 183343 103864
rect 179860 103806 183343 103808
rect 183277 103803 183343 103806
rect 117957 103186 118023 103189
rect 117957 103184 120060 103186
rect 117957 103128 117962 103184
rect 118018 103128 120060 103184
rect 117957 103126 120060 103128
rect 117957 103123 118023 103126
rect 183277 102506 183343 102509
rect 179860 102504 183343 102506
rect 179860 102448 183282 102504
rect 183338 102448 183343 102504
rect 179860 102446 183343 102448
rect 183277 102443 183343 102446
rect 120809 102098 120875 102101
rect 120582 102096 120875 102098
rect 120582 102040 120814 102096
rect 120870 102040 120875 102096
rect 120582 102038 120875 102040
rect 120582 101660 120642 102038
rect 120809 102035 120875 102038
rect 183277 101146 183343 101149
rect 179860 101144 183343 101146
rect 179860 101088 183282 101144
rect 183338 101088 183343 101144
rect 179860 101086 183343 101088
rect 183277 101083 183343 101086
rect 118785 100194 118851 100197
rect 118785 100192 120060 100194
rect 118785 100136 118790 100192
rect 118846 100136 120060 100192
rect 118785 100134 120060 100136
rect 118785 100131 118851 100134
rect 183185 99786 183251 99789
rect 179860 99784 183251 99786
rect 179860 99728 183190 99784
rect 183246 99728 183251 99784
rect 179860 99726 183251 99728
rect 183185 99723 183251 99726
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 118693 98698 118759 98701
rect 118693 98696 120060 98698
rect 118693 98640 118698 98696
rect 118754 98640 120060 98696
rect 118693 98638 120060 98640
rect 118693 98635 118759 98638
rect 183185 98426 183251 98429
rect 179860 98424 183251 98426
rect 179860 98368 183190 98424
rect 183246 98368 183251 98424
rect 179860 98366 183251 98368
rect 183185 98363 183251 98366
rect 120717 97746 120783 97749
rect 120582 97744 120783 97746
rect -960 97610 480 97700
rect 120582 97688 120722 97744
rect 120778 97688 120783 97744
rect 120582 97686 120783 97688
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 120582 97172 120642 97686
rect 120717 97683 120783 97686
rect 183185 97066 183251 97069
rect 179860 97064 183251 97066
rect 179860 97008 183190 97064
rect 183246 97008 183251 97064
rect 179860 97006 183251 97008
rect 183185 97003 183251 97006
rect 118233 95706 118299 95709
rect 183185 95706 183251 95709
rect 118233 95704 120060 95706
rect 118233 95648 118238 95704
rect 118294 95648 120060 95704
rect 118233 95646 120060 95648
rect 179860 95704 183251 95706
rect 179860 95648 183190 95704
rect 183246 95648 183251 95704
rect 179860 95646 183251 95648
rect 118233 95643 118299 95646
rect 183185 95643 183251 95646
rect 183461 94346 183527 94349
rect 179860 94344 183527 94346
rect 179860 94288 183466 94344
rect 183522 94288 183527 94344
rect 179860 94286 183527 94288
rect 183461 94283 183527 94286
rect 118325 94210 118391 94213
rect 118325 94208 120060 94210
rect 118325 94152 118330 94208
rect 118386 94152 120060 94208
rect 118325 94150 120060 94152
rect 118325 94147 118391 94150
rect 183461 92986 183527 92989
rect 179860 92984 183527 92986
rect 179860 92928 183466 92984
rect 183522 92928 183527 92984
rect 179860 92926 183527 92928
rect 183461 92923 183527 92926
rect 118509 92714 118575 92717
rect 118509 92712 120060 92714
rect 118509 92656 118514 92712
rect 118570 92656 120060 92712
rect 118509 92654 120060 92656
rect 118509 92651 118575 92654
rect 183461 91626 183527 91629
rect 179860 91624 183527 91626
rect 179860 91568 183466 91624
rect 183522 91568 183527 91624
rect 179860 91566 183527 91568
rect 183461 91563 183527 91566
rect 118417 91218 118483 91221
rect 118417 91216 120060 91218
rect 118417 91160 118422 91216
rect 118478 91160 120060 91216
rect 118417 91158 120060 91160
rect 118417 91155 118483 91158
rect 183461 90266 183527 90269
rect 179860 90264 183527 90266
rect 179860 90208 183466 90264
rect 183522 90208 183527 90264
rect 179860 90206 183527 90208
rect 183461 90203 183527 90206
rect 118049 89722 118115 89725
rect 118049 89720 120060 89722
rect 118049 89664 118054 89720
rect 118110 89664 120060 89720
rect 118049 89662 120060 89664
rect 118049 89659 118115 89662
rect 183461 88906 183527 88909
rect 179860 88904 183527 88906
rect 179860 88848 183466 88904
rect 183522 88848 183527 88904
rect 179860 88846 183527 88848
rect 183461 88843 183527 88846
rect 118141 88226 118207 88229
rect 118141 88224 120060 88226
rect 118141 88168 118146 88224
rect 118202 88168 120060 88224
rect 118141 88166 120060 88168
rect 118141 88163 118207 88166
rect 183461 87546 183527 87549
rect 179860 87544 183527 87546
rect 179860 87488 183466 87544
rect 183522 87488 183527 87544
rect 179860 87486 183527 87488
rect 183461 87483 183527 87486
rect 118509 86730 118575 86733
rect 118509 86728 120060 86730
rect 118509 86672 118514 86728
rect 118570 86672 120060 86728
rect 118509 86670 120060 86672
rect 118509 86667 118575 86670
rect 182541 86186 182607 86189
rect 179860 86184 182607 86186
rect 179860 86128 182546 86184
rect 182602 86128 182607 86184
rect 179860 86126 182607 86128
rect 182541 86123 182607 86126
rect 579981 86186 580047 86189
rect 583520 86186 584960 86276
rect 579981 86184 584960 86186
rect 579981 86128 579986 86184
rect 580042 86128 584960 86184
rect 579981 86126 584960 86128
rect 579981 86123 580047 86126
rect 583520 86036 584960 86126
rect 118601 85234 118667 85237
rect 118601 85232 120060 85234
rect 118601 85176 118606 85232
rect 118662 85176 120060 85232
rect 118601 85174 120060 85176
rect 118601 85171 118667 85174
rect 182725 84826 182791 84829
rect 179860 84824 182791 84826
rect -960 84690 480 84780
rect 179860 84768 182730 84824
rect 182786 84768 182791 84824
rect 179860 84766 182791 84768
rect 182725 84763 182791 84766
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 118417 83738 118483 83741
rect 118417 83736 120060 83738
rect 118417 83680 118422 83736
rect 118478 83680 120060 83736
rect 118417 83678 120060 83680
rect 118417 83675 118483 83678
rect 182817 83466 182883 83469
rect 179860 83464 182883 83466
rect 179860 83408 182822 83464
rect 182878 83408 182883 83464
rect 179860 83406 182883 83408
rect 182817 83403 182883 83406
rect 118325 82242 118391 82245
rect 118325 82240 120060 82242
rect 118325 82184 118330 82240
rect 118386 82184 120060 82240
rect 118325 82182 120060 82184
rect 118325 82179 118391 82182
rect 182817 82106 182883 82109
rect 179860 82104 182883 82106
rect 179860 82048 182822 82104
rect 182878 82048 182883 82104
rect 179860 82046 182883 82048
rect 182817 82043 182883 82046
rect 182173 80746 182239 80749
rect 179860 80744 182239 80746
rect 179860 80688 182178 80744
rect 182234 80688 182239 80744
rect 179860 80686 182239 80688
rect 182173 80683 182239 80686
rect 168046 80548 168052 80612
rect 168116 80610 168122 80612
rect 174905 80610 174971 80613
rect 396901 80610 396967 80613
rect 168116 80608 174971 80610
rect 168116 80552 174910 80608
rect 174966 80552 174971 80608
rect 168116 80550 174971 80552
rect 168116 80548 168122 80550
rect 174905 80547 174971 80550
rect 180750 80608 396967 80610
rect 180750 80552 396906 80608
rect 396962 80552 396967 80608
rect 180750 80550 396967 80552
rect 118509 80474 118575 80477
rect 180057 80474 180123 80477
rect 118509 80472 180123 80474
rect 118509 80416 118514 80472
rect 118570 80416 180062 80472
rect 180118 80416 180123 80472
rect 118509 80414 180123 80416
rect 118509 80411 118575 80414
rect 180057 80411 180123 80414
rect 172278 80276 172284 80340
rect 172348 80338 172354 80340
rect 174537 80338 174603 80341
rect 172348 80336 174603 80338
rect 172348 80280 174542 80336
rect 174598 80280 174603 80336
rect 172348 80278 174603 80280
rect 172348 80276 172354 80278
rect 174537 80275 174603 80278
rect 123477 80202 123543 80205
rect 123477 80200 131360 80202
rect 123477 80144 123482 80200
rect 123538 80144 131360 80200
rect 123477 80142 131360 80144
rect 123477 80139 123543 80142
rect 125823 79962 125889 79967
rect 125542 79868 125548 79932
rect 125612 79930 125618 79932
rect 125823 79930 125828 79962
rect 125612 79906 125828 79930
rect 125884 79906 125889 79962
rect 129503 79964 129569 79967
rect 131159 79964 131225 79967
rect 129503 79962 129704 79964
rect 128031 79930 128097 79933
rect 125612 79901 125889 79906
rect 126148 79928 128097 79930
rect 125612 79870 125886 79901
rect 126148 79872 128036 79928
rect 128092 79872 128097 79928
rect 126148 79870 128097 79872
rect 125612 79868 125618 79870
rect 122373 79794 122439 79797
rect 126148 79794 126208 79870
rect 128031 79867 128097 79870
rect 128399 79928 128465 79933
rect 128675 79932 128741 79933
rect 129043 79932 129109 79933
rect 128670 79930 128676 79932
rect 128399 79872 128404 79928
rect 128460 79872 128465 79928
rect 128399 79867 128465 79872
rect 128584 79870 128676 79930
rect 128670 79868 128676 79870
rect 128740 79868 128746 79932
rect 129038 79930 129044 79932
rect 128952 79870 129044 79930
rect 129038 79868 129044 79870
rect 129108 79868 129114 79932
rect 129503 79906 129508 79962
rect 129564 79906 129704 79962
rect 130886 79962 131225 79964
rect 129503 79904 129704 79906
rect 129503 79901 129569 79904
rect 128675 79867 128741 79868
rect 129043 79867 129109 79868
rect 127019 79796 127085 79797
rect 127014 79794 127020 79796
rect 122373 79792 126208 79794
rect 122373 79736 122378 79792
rect 122434 79736 126208 79792
rect 122373 79734 126208 79736
rect 126928 79734 127020 79794
rect 122373 79731 122439 79734
rect 127014 79732 127020 79734
rect 127084 79732 127090 79796
rect 128402 79794 128462 79867
rect 128670 79794 128676 79796
rect 128402 79734 128676 79794
rect 128670 79732 128676 79734
rect 128740 79732 128746 79796
rect 129457 79794 129523 79797
rect 129644 79794 129704 79904
rect 129774 79868 129780 79932
rect 129844 79930 129850 79932
rect 129963 79930 130029 79933
rect 130699 79930 130765 79933
rect 130886 79932 131164 79962
rect 129844 79928 130029 79930
rect 129844 79872 129968 79928
rect 130024 79872 130029 79928
rect 129844 79870 130029 79872
rect 129844 79868 129850 79870
rect 129963 79867 130029 79870
rect 130518 79928 130765 79930
rect 130518 79872 130704 79928
rect 130760 79872 130765 79928
rect 130518 79870 130765 79872
rect 130285 79794 130351 79797
rect 129457 79792 129704 79794
rect 129457 79736 129462 79792
rect 129518 79736 129704 79792
rect 129457 79734 129704 79736
rect 129920 79792 130351 79794
rect 129920 79736 130290 79792
rect 130346 79736 130351 79792
rect 129920 79734 130351 79736
rect 127019 79731 127085 79732
rect 129457 79731 129523 79734
rect 129920 79661 129980 79734
rect 130285 79731 130351 79734
rect 129917 79656 129983 79661
rect 129917 79600 129922 79656
rect 129978 79600 129983 79656
rect 129917 79595 129983 79600
rect 130285 79658 130351 79661
rect 130518 79658 130578 79870
rect 130699 79867 130765 79870
rect 130878 79868 130884 79932
rect 130948 79906 131164 79932
rect 131220 79906 131225 79962
rect 130948 79904 131225 79906
rect 130948 79868 130954 79904
rect 131159 79901 131225 79904
rect 131300 79930 131360 80142
rect 161974 80140 161980 80204
rect 162044 80202 162050 80204
rect 180750 80202 180810 80550
rect 396901 80547 396967 80550
rect 162044 80142 168712 80202
rect 162044 80140 162050 80142
rect 160134 80066 160140 80068
rect 158854 80006 160140 80066
rect 131711 79964 131777 79967
rect 131668 79962 131777 79964
rect 131527 79930 131593 79933
rect 131300 79928 131593 79930
rect 131300 79872 131532 79928
rect 131588 79872 131593 79928
rect 131300 79870 131593 79872
rect 131527 79867 131593 79870
rect 131668 79906 131716 79962
rect 131772 79906 131777 79962
rect 132815 79964 132881 79967
rect 132815 79962 132924 79964
rect 131668 79901 131777 79906
rect 132539 79928 132605 79933
rect 131251 79796 131317 79797
rect 131246 79794 131252 79796
rect 131160 79734 131252 79794
rect 131246 79732 131252 79734
rect 131316 79732 131322 79796
rect 131668 79794 131728 79901
rect 132171 79894 132237 79899
rect 132171 79838 132176 79894
rect 132232 79838 132237 79894
rect 132539 79872 132544 79928
rect 132600 79872 132605 79928
rect 132815 79906 132820 79962
rect 132876 79930 132924 79962
rect 133643 79962 133709 79967
rect 133086 79930 133092 79932
rect 132876 79906 133092 79930
rect 132815 79901 133092 79906
rect 132539 79867 132605 79872
rect 132864 79870 133092 79901
rect 133086 79868 133092 79870
rect 133156 79868 133162 79932
rect 133270 79868 133276 79932
rect 133340 79930 133346 79932
rect 133643 79930 133648 79962
rect 133340 79906 133648 79930
rect 133704 79906 133709 79962
rect 134011 79962 134077 79967
rect 133340 79901 133709 79906
rect 133340 79870 133706 79901
rect 133340 79868 133346 79870
rect 133822 79868 133828 79932
rect 133892 79930 133898 79932
rect 134011 79930 134016 79962
rect 133892 79906 134016 79930
rect 134072 79906 134077 79962
rect 133892 79901 134077 79906
rect 134195 79962 134261 79967
rect 134195 79906 134200 79962
rect 134256 79906 134261 79962
rect 134195 79901 134261 79906
rect 134655 79962 134721 79967
rect 134655 79906 134660 79962
rect 134716 79906 134721 79962
rect 135483 79962 135549 79967
rect 135483 79932 135488 79962
rect 135544 79932 135549 79962
rect 136587 79962 136653 79967
rect 134655 79901 134721 79906
rect 133892 79870 134074 79901
rect 133892 79868 133898 79870
rect 132171 79833 132237 79838
rect 131392 79734 131728 79794
rect 131251 79731 131317 79732
rect 130285 79656 130578 79658
rect 130285 79600 130290 79656
rect 130346 79600 130578 79656
rect 130285 79598 130578 79600
rect 131205 79658 131271 79661
rect 131392 79658 131452 79734
rect 131205 79656 131452 79658
rect 131205 79600 131210 79656
rect 131266 79600 131452 79656
rect 131205 79598 131452 79600
rect 131573 79658 131639 79661
rect 132174 79658 132234 79833
rect 132542 79661 132602 79867
rect 134198 79794 134258 79901
rect 134658 79797 134718 79901
rect 135478 79868 135484 79932
rect 135548 79930 135554 79932
rect 135943 79930 136009 79933
rect 135548 79870 135606 79930
rect 135943 79928 136052 79930
rect 135943 79872 135948 79928
rect 136004 79872 136052 79928
rect 135548 79868 135554 79870
rect 135943 79867 136052 79872
rect 136214 79868 136220 79932
rect 136284 79930 136290 79932
rect 136587 79930 136592 79962
rect 136284 79906 136592 79930
rect 136648 79906 136653 79962
rect 137967 79962 138033 79967
rect 137047 79930 137113 79933
rect 136284 79901 136653 79906
rect 137004 79928 137113 79930
rect 136284 79870 136650 79901
rect 137004 79872 137052 79928
rect 137108 79872 137113 79928
rect 136284 79868 136290 79870
rect 135115 79826 135181 79831
rect 134333 79794 134399 79797
rect 134198 79792 134399 79794
rect 134198 79736 134338 79792
rect 134394 79736 134399 79792
rect 134198 79734 134399 79736
rect 134333 79731 134399 79734
rect 134655 79792 134721 79797
rect 134655 79736 134660 79792
rect 134716 79736 134721 79792
rect 135115 79770 135120 79826
rect 135176 79770 135181 79826
rect 135115 79765 135181 79770
rect 134655 79731 134721 79736
rect 135118 79661 135178 79765
rect 135992 79661 136052 79867
rect 137004 79867 137113 79872
rect 137686 79868 137692 79932
rect 137756 79930 137762 79932
rect 137967 79930 137972 79962
rect 137756 79906 137972 79930
rect 138028 79906 138033 79962
rect 138795 79962 138861 79967
rect 137756 79901 138033 79906
rect 138151 79930 138217 79933
rect 138151 79928 138352 79930
rect 137756 79870 138030 79901
rect 138151 79872 138156 79928
rect 138212 79872 138352 79928
rect 138151 79870 138352 79872
rect 137756 79868 137762 79870
rect 138151 79867 138217 79870
rect 137004 79796 137064 79867
rect 137921 79796 137987 79797
rect 136950 79732 136956 79796
rect 137020 79734 137064 79796
rect 137870 79794 137876 79796
rect 137830 79734 137876 79794
rect 137940 79792 137987 79796
rect 137982 79736 137987 79792
rect 137020 79732 137026 79734
rect 137870 79732 137876 79734
rect 137940 79732 137987 79736
rect 138054 79732 138060 79796
rect 138124 79794 138130 79796
rect 138292 79794 138352 79870
rect 138611 79928 138677 79933
rect 138611 79872 138616 79928
rect 138672 79872 138677 79928
rect 138795 79906 138800 79962
rect 138856 79930 138861 79962
rect 140819 79962 140885 79967
rect 139347 79932 139413 79933
rect 138974 79930 138980 79932
rect 138856 79906 138980 79930
rect 138795 79901 138980 79906
rect 138611 79867 138677 79872
rect 138798 79870 138980 79901
rect 138974 79868 138980 79870
rect 139044 79868 139050 79932
rect 139342 79930 139348 79932
rect 139256 79870 139348 79930
rect 139342 79868 139348 79870
rect 139412 79868 139418 79932
rect 140819 79906 140824 79962
rect 140880 79906 140885 79962
rect 142015 79962 142081 79967
rect 141463 79930 141529 79933
rect 140819 79901 140885 79906
rect 141328 79928 141529 79930
rect 139531 79894 139597 79899
rect 139347 79867 139413 79868
rect 138614 79797 138674 79867
rect 139531 79838 139536 79894
rect 139592 79838 139597 79894
rect 139531 79833 139597 79838
rect 138124 79734 138352 79794
rect 138565 79792 138674 79797
rect 138565 79736 138570 79792
rect 138626 79736 138674 79792
rect 138565 79734 138674 79736
rect 138124 79732 138130 79734
rect 137921 79731 137987 79732
rect 138565 79731 138631 79734
rect 138790 79732 138796 79796
rect 138860 79794 138866 79796
rect 139163 79794 139229 79797
rect 138860 79792 139229 79794
rect 138860 79736 139168 79792
rect 139224 79736 139229 79792
rect 138860 79734 139229 79736
rect 138860 79732 138866 79734
rect 139163 79731 139229 79734
rect 131573 79656 132234 79658
rect 131573 79600 131578 79656
rect 131634 79600 132234 79656
rect 131573 79598 132234 79600
rect 132493 79656 132602 79661
rect 132493 79600 132498 79656
rect 132554 79600 132602 79656
rect 132493 79598 132602 79600
rect 130285 79595 130351 79598
rect 131205 79595 131271 79598
rect 131573 79595 131639 79598
rect 132493 79595 132559 79598
rect 133638 79596 133644 79660
rect 133708 79658 133714 79660
rect 133965 79658 134031 79661
rect 133708 79656 134031 79658
rect 133708 79600 133970 79656
rect 134026 79600 134031 79656
rect 133708 79598 134031 79600
rect 133708 79596 133714 79598
rect 133965 79595 134031 79598
rect 135069 79656 135178 79661
rect 135069 79600 135074 79656
rect 135130 79600 135178 79656
rect 135069 79598 135178 79600
rect 135989 79656 136055 79661
rect 135989 79600 135994 79656
rect 136050 79600 136055 79656
rect 135069 79595 135135 79598
rect 135989 79595 136055 79600
rect 139393 79658 139459 79661
rect 139534 79658 139594 79833
rect 139393 79656 139594 79658
rect 139393 79600 139398 79656
rect 139454 79600 139594 79656
rect 139393 79598 139594 79600
rect 139393 79595 139459 79598
rect 140078 79596 140084 79660
rect 140148 79658 140154 79660
rect 140313 79658 140379 79661
rect 140148 79656 140379 79658
rect 140148 79600 140318 79656
rect 140374 79600 140379 79656
rect 140148 79598 140379 79600
rect 140148 79596 140154 79598
rect 140313 79595 140379 79598
rect 140681 79658 140747 79661
rect 140822 79658 140882 79901
rect 141328 79872 141468 79928
rect 141524 79872 141529 79928
rect 142015 79906 142020 79962
rect 142076 79930 142081 79962
rect 142475 79962 142541 79967
rect 142751 79964 142817 79967
rect 142286 79930 142292 79932
rect 142076 79906 142292 79930
rect 142015 79901 142292 79906
rect 141328 79870 141529 79872
rect 142018 79870 142292 79901
rect 141328 79794 141388 79870
rect 141463 79867 141529 79870
rect 142286 79868 142292 79870
rect 142356 79868 142362 79932
rect 142475 79906 142480 79962
rect 142536 79906 142541 79962
rect 142475 79901 142541 79906
rect 142708 79962 142817 79964
rect 142708 79906 142756 79962
rect 142812 79906 142817 79962
rect 143763 79962 143829 79967
rect 143395 79930 143461 79933
rect 142708 79901 142817 79906
rect 143352 79928 143461 79930
rect 141509 79794 141575 79797
rect 141328 79792 141575 79794
rect 141328 79736 141514 79792
rect 141570 79736 141575 79792
rect 141328 79734 141575 79736
rect 141509 79731 141575 79734
rect 141918 79732 141924 79796
rect 141988 79794 141994 79796
rect 142061 79794 142127 79797
rect 141988 79792 142127 79794
rect 141988 79736 142066 79792
rect 142122 79736 142127 79792
rect 141988 79734 142127 79736
rect 141988 79732 141994 79734
rect 142061 79731 142127 79734
rect 140681 79656 140882 79658
rect 140681 79600 140686 79656
rect 140742 79600 140882 79656
rect 140681 79598 140882 79600
rect 142061 79658 142127 79661
rect 142478 79658 142538 79901
rect 142708 79797 142768 79901
rect 143352 79872 143400 79928
rect 143456 79872 143461 79928
rect 143352 79867 143461 79872
rect 143579 79928 143645 79933
rect 143579 79872 143584 79928
rect 143640 79872 143645 79928
rect 143763 79906 143768 79962
rect 143824 79906 143829 79962
rect 144315 79962 144381 79967
rect 144039 79930 144105 79933
rect 144315 79932 144320 79962
rect 144376 79932 144381 79962
rect 144867 79962 144933 79967
rect 143763 79901 143829 79906
rect 143996 79928 144105 79930
rect 143579 79867 143645 79872
rect 142705 79792 142771 79797
rect 142705 79736 142710 79792
rect 142766 79736 142771 79792
rect 142705 79731 142771 79736
rect 143206 79732 143212 79796
rect 143276 79794 143282 79796
rect 143352 79794 143412 79867
rect 143276 79734 143412 79794
rect 143276 79732 143282 79734
rect 143582 79661 143642 79867
rect 142061 79656 142538 79658
rect 142061 79600 142066 79656
rect 142122 79600 142538 79656
rect 142061 79598 142538 79600
rect 143533 79656 143642 79661
rect 143533 79600 143538 79656
rect 143594 79600 143642 79656
rect 143533 79598 143642 79600
rect 143766 79661 143826 79901
rect 143996 79872 144044 79928
rect 144100 79872 144105 79928
rect 143996 79867 144105 79872
rect 144310 79868 144316 79932
rect 144380 79930 144386 79932
rect 144380 79870 144438 79930
rect 144867 79906 144872 79962
rect 144928 79906 144933 79962
rect 145051 79962 145117 79967
rect 145051 79932 145056 79962
rect 145112 79932 145117 79962
rect 146707 79962 146773 79967
rect 145787 79932 145853 79933
rect 144867 79901 144933 79906
rect 144380 79868 144386 79870
rect 143996 79794 144056 79867
rect 144870 79797 144930 79901
rect 145046 79868 145052 79932
rect 145116 79930 145122 79932
rect 145782 79930 145788 79932
rect 145116 79870 145174 79930
rect 145696 79870 145788 79930
rect 145116 79868 145122 79870
rect 145782 79868 145788 79870
rect 145852 79868 145858 79932
rect 146150 79868 146156 79932
rect 146220 79930 146226 79932
rect 146431 79930 146497 79933
rect 146220 79928 146497 79930
rect 146220 79872 146436 79928
rect 146492 79872 146497 79928
rect 146707 79906 146712 79962
rect 146768 79906 146773 79962
rect 147443 79962 147509 79967
rect 147259 79932 147325 79933
rect 147254 79930 147260 79932
rect 146707 79901 146773 79906
rect 146220 79870 146497 79872
rect 146220 79868 146226 79870
rect 145787 79867 145853 79868
rect 146431 79867 146497 79870
rect 146710 79797 146770 79901
rect 147168 79870 147260 79930
rect 147254 79868 147260 79870
rect 147324 79868 147330 79932
rect 147443 79906 147448 79962
rect 147504 79906 147509 79962
rect 150663 79964 150729 79967
rect 150663 79962 151002 79964
rect 147443 79901 147509 79906
rect 148271 79930 148337 79933
rect 149559 79930 149625 79933
rect 149830 79930 149836 79932
rect 148271 79928 148610 79930
rect 147259 79867 147325 79868
rect 144269 79794 144335 79797
rect 144499 79796 144565 79797
rect 144494 79794 144500 79796
rect 143996 79792 144335 79794
rect 143996 79736 144274 79792
rect 144330 79736 144335 79792
rect 143996 79734 144335 79736
rect 144408 79734 144500 79794
rect 144269 79731 144335 79734
rect 144494 79732 144500 79734
rect 144564 79732 144570 79796
rect 144867 79792 144933 79797
rect 144867 79736 144872 79792
rect 144928 79736 144933 79792
rect 144499 79731 144565 79732
rect 144867 79731 144933 79736
rect 146710 79792 146819 79797
rect 146710 79736 146758 79792
rect 146814 79736 146819 79792
rect 146710 79734 146819 79736
rect 146753 79731 146819 79734
rect 147446 79661 147506 79901
rect 148271 79872 148276 79928
rect 148332 79872 148610 79928
rect 148271 79870 148610 79872
rect 148271 79867 148337 79870
rect 148225 79796 148291 79797
rect 148174 79732 148180 79796
rect 148244 79794 148291 79796
rect 148244 79792 148336 79794
rect 148286 79736 148336 79792
rect 148244 79734 148336 79736
rect 148244 79732 148291 79734
rect 148225 79731 148291 79732
rect 143766 79656 143875 79661
rect 143766 79600 143814 79656
rect 143870 79600 143875 79656
rect 143766 79598 143875 79600
rect 140681 79595 140747 79598
rect 142061 79595 142127 79598
rect 143533 79595 143599 79598
rect 143809 79595 143875 79598
rect 145598 79596 145604 79660
rect 145668 79658 145674 79660
rect 146017 79658 146083 79661
rect 145668 79656 146083 79658
rect 145668 79600 146022 79656
rect 146078 79600 146083 79656
rect 145668 79598 146083 79600
rect 145668 79596 145674 79598
rect 146017 79595 146083 79598
rect 146518 79596 146524 79660
rect 146588 79658 146594 79660
rect 146661 79658 146727 79661
rect 146588 79656 146727 79658
rect 146588 79600 146666 79656
rect 146722 79600 146727 79656
rect 146588 79598 146727 79600
rect 147446 79656 147555 79661
rect 147446 79600 147494 79656
rect 147550 79600 147555 79656
rect 147446 79598 147555 79600
rect 146588 79596 146594 79598
rect 146661 79595 146727 79598
rect 147489 79595 147555 79598
rect 148317 79658 148383 79661
rect 148550 79658 148610 79870
rect 149559 79928 149836 79930
rect 149559 79872 149564 79928
rect 149620 79872 149836 79928
rect 149559 79870 149836 79872
rect 149559 79867 149625 79870
rect 149830 79868 149836 79870
rect 149900 79868 149906 79932
rect 150111 79930 150177 79933
rect 150068 79928 150177 79930
rect 150068 79872 150116 79928
rect 150172 79872 150177 79928
rect 150663 79906 150668 79962
rect 150724 79932 151002 79962
rect 151675 79962 151741 79967
rect 150724 79906 150940 79932
rect 150663 79904 150940 79906
rect 150663 79901 150729 79904
rect 150068 79867 150177 79872
rect 150934 79868 150940 79904
rect 151004 79868 151010 79932
rect 151215 79930 151281 79933
rect 151080 79928 151281 79930
rect 151080 79872 151220 79928
rect 151276 79872 151281 79928
rect 151675 79906 151680 79962
rect 151736 79906 151741 79962
rect 152319 79962 152385 79967
rect 151675 79901 151741 79906
rect 151951 79930 152017 79933
rect 151951 79928 152152 79930
rect 151080 79870 151281 79872
rect 148726 79732 148732 79796
rect 148796 79794 148802 79796
rect 148915 79794 148981 79797
rect 148796 79792 148981 79794
rect 148796 79736 148920 79792
rect 148976 79736 148981 79792
rect 148796 79734 148981 79736
rect 148796 79732 148802 79734
rect 148915 79731 148981 79734
rect 149646 79732 149652 79796
rect 149716 79794 149722 79796
rect 150068 79794 150128 79867
rect 149716 79734 150128 79794
rect 150893 79794 150959 79797
rect 151080 79794 151140 79870
rect 151215 79867 151281 79870
rect 150893 79792 151140 79794
rect 150893 79736 150898 79792
rect 150954 79736 151140 79792
rect 150893 79734 151140 79736
rect 149716 79732 149722 79734
rect 150893 79731 150959 79734
rect 151486 79732 151492 79796
rect 151556 79794 151562 79796
rect 151678 79794 151738 79901
rect 151951 79872 151956 79928
rect 152012 79872 152152 79928
rect 152319 79906 152324 79962
rect 152380 79906 152385 79962
rect 152319 79901 152385 79906
rect 152595 79962 152661 79967
rect 153423 79964 153489 79967
rect 152595 79906 152600 79962
rect 152656 79930 152661 79962
rect 153380 79962 153489 79964
rect 152774 79930 152780 79932
rect 152656 79906 152780 79930
rect 152595 79901 152780 79906
rect 151951 79870 152152 79872
rect 151951 79867 152017 79870
rect 152092 79796 152152 79870
rect 151556 79734 151738 79794
rect 151556 79732 151562 79734
rect 152038 79732 152044 79796
rect 152108 79734 152152 79796
rect 152108 79732 152114 79734
rect 148317 79656 148610 79658
rect 148317 79600 148322 79656
rect 148378 79600 148610 79656
rect 148317 79598 148610 79600
rect 152089 79658 152155 79661
rect 152322 79658 152382 79901
rect 152598 79870 152780 79901
rect 152774 79868 152780 79870
rect 152844 79868 152850 79932
rect 153380 79906 153428 79962
rect 153484 79930 153489 79962
rect 154987 79962 155053 79967
rect 153694 79930 153700 79932
rect 153484 79906 153700 79930
rect 153380 79870 153700 79906
rect 153694 79868 153700 79870
rect 153764 79868 153770 79932
rect 153975 79930 154041 79933
rect 154435 79932 154501 79933
rect 154619 79932 154685 79933
rect 154430 79930 154436 79932
rect 153975 79928 154176 79930
rect 153975 79872 153980 79928
rect 154036 79872 154176 79928
rect 153975 79870 154176 79872
rect 154344 79870 154436 79930
rect 153975 79867 154041 79870
rect 152590 79732 152596 79796
rect 152660 79794 152666 79796
rect 152733 79794 152799 79797
rect 153791 79794 153857 79797
rect 152660 79792 152799 79794
rect 152660 79736 152738 79792
rect 152794 79736 152799 79792
rect 152660 79734 152799 79736
rect 152660 79732 152666 79734
rect 152733 79731 152799 79734
rect 153610 79792 153857 79794
rect 153610 79736 153796 79792
rect 153852 79736 153857 79792
rect 153610 79734 153857 79736
rect 154116 79794 154176 79870
rect 154430 79868 154436 79870
rect 154500 79868 154506 79932
rect 154614 79868 154620 79932
rect 154684 79930 154690 79932
rect 154684 79870 154776 79930
rect 154987 79906 154992 79962
rect 155048 79906 155053 79962
rect 154987 79901 155053 79906
rect 155171 79962 155237 79967
rect 155631 79964 155697 79967
rect 155171 79906 155176 79962
rect 155232 79906 155237 79962
rect 155588 79962 155697 79964
rect 155355 79932 155421 79933
rect 155171 79901 155237 79906
rect 154684 79868 154690 79870
rect 154435 79867 154501 79868
rect 154619 79867 154685 79868
rect 154246 79794 154252 79796
rect 154116 79734 154252 79794
rect 153610 79661 153670 79734
rect 153791 79731 153857 79734
rect 154246 79732 154252 79734
rect 154316 79732 154322 79796
rect 152089 79656 152382 79658
rect 152089 79600 152094 79656
rect 152150 79600 152382 79656
rect 152089 79598 152382 79600
rect 153561 79656 153670 79661
rect 153561 79600 153566 79656
rect 153622 79600 153670 79656
rect 153561 79598 153670 79600
rect 154757 79658 154823 79661
rect 154990 79658 155050 79901
rect 155174 79797 155234 79901
rect 155350 79868 155356 79932
rect 155420 79930 155426 79932
rect 155420 79870 155512 79930
rect 155588 79906 155636 79962
rect 155692 79906 155697 79962
rect 155588 79901 155697 79906
rect 155815 79962 155881 79967
rect 155815 79906 155820 79962
rect 155876 79906 155881 79962
rect 155815 79901 155881 79906
rect 156091 79962 156157 79967
rect 156091 79906 156096 79962
rect 156152 79906 156157 79962
rect 156091 79901 156157 79906
rect 156551 79964 156617 79967
rect 156551 79962 156844 79964
rect 156551 79906 156556 79962
rect 156612 79906 156844 79962
rect 157379 79962 157445 79967
rect 158391 79964 158457 79967
rect 157379 79932 157384 79962
rect 157440 79932 157445 79962
rect 158348 79962 158457 79964
rect 156551 79904 156844 79906
rect 156551 79901 156617 79904
rect 155420 79868 155426 79870
rect 155355 79867 155421 79868
rect 155125 79792 155234 79797
rect 155125 79736 155130 79792
rect 155186 79736 155234 79792
rect 155125 79734 155234 79736
rect 155125 79731 155191 79734
rect 154757 79656 155050 79658
rect 154757 79600 154762 79656
rect 154818 79600 155050 79656
rect 154757 79598 155050 79600
rect 155588 79658 155648 79901
rect 155818 79797 155878 79901
rect 155769 79792 155878 79797
rect 155769 79736 155774 79792
rect 155830 79736 155878 79792
rect 155769 79734 155878 79736
rect 155769 79731 155835 79734
rect 156094 79661 156154 79901
rect 156784 79797 156844 79904
rect 157103 79896 157169 79899
rect 157060 79894 157169 79896
rect 157060 79838 157108 79894
rect 157164 79838 157169 79894
rect 157374 79868 157380 79932
rect 157444 79930 157450 79932
rect 157444 79870 157502 79930
rect 157444 79868 157450 79870
rect 158110 79868 158116 79932
rect 158180 79930 158186 79932
rect 158348 79930 158396 79962
rect 158180 79906 158396 79930
rect 158452 79906 158457 79962
rect 158667 79962 158733 79967
rect 158667 79932 158672 79962
rect 158728 79932 158733 79962
rect 158180 79901 158457 79906
rect 158180 79870 158408 79901
rect 158180 79868 158186 79870
rect 158662 79868 158668 79932
rect 158732 79930 158738 79932
rect 158732 79870 158790 79930
rect 158732 79868 158738 79870
rect 157060 79833 157169 79838
rect 156275 79796 156341 79797
rect 156270 79732 156276 79796
rect 156340 79794 156346 79796
rect 156340 79734 156432 79794
rect 156781 79792 156847 79797
rect 156781 79736 156786 79792
rect 156842 79736 156847 79792
rect 156340 79732 156346 79734
rect 156275 79731 156341 79732
rect 156781 79731 156847 79736
rect 155718 79658 155724 79660
rect 155588 79598 155724 79658
rect 148317 79595 148383 79598
rect 152089 79595 152155 79598
rect 153561 79595 153627 79598
rect 154757 79595 154823 79598
rect 155718 79596 155724 79598
rect 155788 79596 155794 79660
rect 156094 79656 156203 79661
rect 156094 79600 156142 79656
rect 156198 79600 156203 79656
rect 156094 79598 156203 79600
rect 156137 79595 156203 79598
rect 156822 79596 156828 79660
rect 156892 79658 156898 79660
rect 157060 79658 157120 79833
rect 157926 79732 157932 79796
rect 157996 79794 158002 79796
rect 158115 79794 158181 79797
rect 157996 79792 158181 79794
rect 157996 79736 158120 79792
rect 158176 79736 158181 79792
rect 157996 79734 158181 79736
rect 157996 79732 158002 79734
rect 158115 79731 158181 79734
rect 158294 79732 158300 79796
rect 158364 79794 158370 79796
rect 158575 79794 158641 79797
rect 158364 79792 158641 79794
rect 158364 79736 158580 79792
rect 158636 79736 158641 79792
rect 158364 79734 158641 79736
rect 158364 79732 158370 79734
rect 158575 79731 158641 79734
rect 158713 79794 158779 79797
rect 158854 79794 158914 80006
rect 160134 80004 160140 80006
rect 160204 80004 160210 80068
rect 161059 79964 161125 79967
rect 161059 79962 161182 79964
rect 159219 79928 159285 79933
rect 159955 79932 160021 79933
rect 160507 79932 160573 79933
rect 161059 79932 161064 79962
rect 161120 79932 161182 79962
rect 161519 79962 161585 79967
rect 159950 79930 159956 79932
rect 159219 79872 159224 79928
rect 159280 79872 159285 79928
rect 159219 79867 159285 79872
rect 159864 79870 159956 79930
rect 159950 79868 159956 79870
rect 160020 79868 160026 79932
rect 160502 79930 160508 79932
rect 160416 79870 160508 79930
rect 160502 79868 160508 79870
rect 160572 79868 160578 79932
rect 161054 79868 161060 79932
rect 161124 79904 161182 79932
rect 161243 79928 161309 79933
rect 161124 79868 161130 79904
rect 161243 79872 161248 79928
rect 161304 79872 161309 79928
rect 161519 79906 161524 79962
rect 161580 79906 161585 79962
rect 161519 79901 161585 79906
rect 161703 79964 161769 79967
rect 161703 79962 162042 79964
rect 161703 79906 161708 79962
rect 161764 79930 162042 79962
rect 165751 79962 165817 79967
rect 162710 79930 162716 79932
rect 161764 79906 162716 79930
rect 161703 79904 162716 79906
rect 161703 79901 161769 79904
rect 159955 79867 160021 79868
rect 160507 79867 160573 79868
rect 161243 79867 161309 79872
rect 158713 79792 158914 79794
rect 158713 79736 158718 79792
rect 158774 79736 158914 79792
rect 158713 79734 158914 79736
rect 159222 79794 159282 79867
rect 160093 79794 160159 79797
rect 159222 79792 160159 79794
rect 159222 79736 160098 79792
rect 160154 79736 160159 79792
rect 159222 79734 160159 79736
rect 158713 79731 158779 79734
rect 160093 79731 160159 79734
rect 161054 79732 161060 79796
rect 161124 79794 161130 79796
rect 161246 79794 161306 79867
rect 161124 79734 161306 79794
rect 161522 79794 161582 79901
rect 161982 79870 162716 79904
rect 162710 79868 162716 79870
rect 162780 79868 162786 79932
rect 162899 79930 162965 79933
rect 162899 79928 163330 79930
rect 162899 79872 162904 79928
rect 162960 79872 163330 79928
rect 162899 79870 163330 79872
rect 162899 79867 162965 79870
rect 161790 79794 161796 79796
rect 161522 79734 161796 79794
rect 161124 79732 161130 79734
rect 161790 79732 161796 79734
rect 161860 79732 161866 79796
rect 162342 79732 162348 79796
rect 162412 79794 162418 79796
rect 162715 79794 162781 79797
rect 162945 79794 163011 79797
rect 162412 79792 162781 79794
rect 162412 79736 162720 79792
rect 162776 79736 162781 79792
rect 162412 79734 162781 79736
rect 162412 79732 162418 79734
rect 162715 79731 162781 79734
rect 162902 79792 163011 79794
rect 162902 79736 162950 79792
rect 163006 79736 163011 79792
rect 162902 79731 163011 79736
rect 156892 79598 157120 79658
rect 156892 79596 156898 79598
rect 157190 79596 157196 79660
rect 157260 79658 157266 79660
rect 157425 79658 157491 79661
rect 157260 79656 157491 79658
rect 157260 79600 157430 79656
rect 157486 79600 157491 79656
rect 157260 79598 157491 79600
rect 157260 79596 157266 79598
rect 157425 79595 157491 79598
rect 158345 79658 158411 79661
rect 158478 79658 158484 79660
rect 158345 79656 158484 79658
rect 158345 79600 158350 79656
rect 158406 79600 158484 79656
rect 158345 79598 158484 79600
rect 158345 79595 158411 79598
rect 158478 79596 158484 79598
rect 158548 79596 158554 79660
rect 159030 79596 159036 79660
rect 159100 79658 159106 79660
rect 159357 79658 159423 79661
rect 159100 79656 159423 79658
rect 159100 79600 159362 79656
rect 159418 79600 159423 79656
rect 159100 79598 159423 79600
rect 162902 79658 162962 79731
rect 163037 79658 163103 79661
rect 162902 79656 163103 79658
rect 162902 79600 163042 79656
rect 163098 79600 163103 79656
rect 162902 79598 163103 79600
rect 163270 79658 163330 79870
rect 163446 79868 163452 79932
rect 163516 79930 163522 79932
rect 164003 79930 164069 79933
rect 163516 79928 164069 79930
rect 163516 79872 164008 79928
rect 164064 79872 164069 79928
rect 163516 79870 164069 79872
rect 163516 79868 163522 79870
rect 164003 79867 164069 79870
rect 164236 79899 164710 79930
rect 164236 79894 164713 79899
rect 164236 79870 164652 79894
rect 163630 79732 163636 79796
rect 163700 79794 163706 79796
rect 164095 79794 164161 79797
rect 163700 79792 164161 79794
rect 163700 79736 164100 79792
rect 164156 79736 164161 79792
rect 163700 79734 164161 79736
rect 163700 79732 163706 79734
rect 164095 79731 164161 79734
rect 164236 79661 164296 79870
rect 164647 79838 164652 79870
rect 164708 79838 164713 79894
rect 165102 79868 165108 79932
rect 165172 79930 165178 79932
rect 165567 79930 165633 79933
rect 165172 79928 165633 79930
rect 165172 79872 165572 79928
rect 165628 79872 165633 79928
rect 165751 79906 165756 79962
rect 165812 79906 165817 79962
rect 168419 79962 168485 79967
rect 166395 79932 166461 79933
rect 166390 79930 166396 79932
rect 165751 79901 165817 79906
rect 165172 79870 165633 79872
rect 165172 79868 165178 79870
rect 165567 79867 165633 79870
rect 164647 79833 164713 79838
rect 165475 79796 165541 79797
rect 165470 79732 165476 79796
rect 165540 79794 165546 79796
rect 165540 79734 165632 79794
rect 165540 79732 165546 79734
rect 165475 79731 165541 79732
rect 163681 79658 163747 79661
rect 163270 79656 163747 79658
rect 163270 79600 163686 79656
rect 163742 79600 163747 79656
rect 163270 79598 163747 79600
rect 159100 79596 159106 79598
rect 159357 79595 159423 79598
rect 163037 79595 163103 79598
rect 163681 79595 163747 79598
rect 164233 79656 164299 79661
rect 164233 79600 164238 79656
rect 164294 79600 164299 79656
rect 164233 79595 164299 79600
rect 164417 79658 164483 79661
rect 164969 79660 165035 79661
rect 164734 79658 164740 79660
rect 164417 79656 164740 79658
rect 164417 79600 164422 79656
rect 164478 79600 164740 79656
rect 164417 79598 164740 79600
rect 164417 79595 164483 79598
rect 164734 79596 164740 79598
rect 164804 79596 164810 79660
rect 164918 79658 164924 79660
rect 164878 79598 164924 79658
rect 164988 79656 165035 79660
rect 165030 79600 165035 79656
rect 164918 79596 164924 79598
rect 164988 79596 165035 79600
rect 165754 79658 165814 79901
rect 166304 79870 166396 79930
rect 166390 79868 166396 79870
rect 166460 79868 166466 79932
rect 166579 79928 166645 79933
rect 166579 79872 166584 79928
rect 166640 79872 166645 79928
rect 166395 79867 166461 79868
rect 166579 79867 166645 79872
rect 166758 79868 166764 79932
rect 166828 79930 166834 79932
rect 166947 79930 167013 79933
rect 167683 79930 167749 79933
rect 166828 79928 167013 79930
rect 166828 79872 166952 79928
rect 167008 79872 167013 79928
rect 166828 79870 167013 79872
rect 166828 79868 166834 79870
rect 166947 79867 167013 79870
rect 167180 79928 167749 79930
rect 167180 79872 167688 79928
rect 167744 79872 167749 79928
rect 167180 79870 167749 79872
rect 166073 79658 166139 79661
rect 165754 79656 166139 79658
rect 165754 79600 166078 79656
rect 166134 79600 166139 79656
rect 165754 79598 166139 79600
rect 166582 79658 166642 79867
rect 167180 79661 167240 79870
rect 167683 79867 167749 79870
rect 167862 79868 167868 79932
rect 167932 79930 167938 79932
rect 168143 79930 168209 79933
rect 168419 79932 168424 79962
rect 168480 79932 168485 79962
rect 167932 79928 168209 79930
rect 167932 79872 168148 79928
rect 168204 79872 168209 79928
rect 167932 79870 168209 79872
rect 167932 79868 167938 79870
rect 168143 79867 168209 79870
rect 168414 79868 168420 79932
rect 168484 79930 168490 79932
rect 168484 79870 168542 79930
rect 168484 79868 168490 79870
rect 168327 79792 168393 79797
rect 168327 79736 168332 79792
rect 168388 79736 168393 79792
rect 168327 79731 168393 79736
rect 168652 79794 168712 80142
rect 171458 80142 180810 80202
rect 171458 79967 171518 80142
rect 462313 80066 462379 80069
rect 180750 80064 462379 80066
rect 180750 80008 462318 80064
rect 462374 80008 462379 80064
rect 180750 80006 462379 80008
rect 168971 79962 169037 79967
rect 168971 79932 168976 79962
rect 169032 79932 169037 79962
rect 169891 79962 169957 79967
rect 168966 79868 168972 79932
rect 169036 79930 169042 79932
rect 169036 79870 169094 79930
rect 169036 79868 169042 79870
rect 169518 79868 169524 79932
rect 169588 79930 169594 79932
rect 169707 79930 169773 79933
rect 169891 79932 169896 79962
rect 169952 79932 169957 79962
rect 170443 79962 170509 79967
rect 170443 79932 170448 79962
rect 170504 79932 170509 79962
rect 171455 79962 171521 79967
rect 170811 79932 170877 79933
rect 171179 79932 171245 79933
rect 169588 79928 169773 79930
rect 169588 79872 169712 79928
rect 169768 79872 169773 79928
rect 169588 79870 169773 79872
rect 169588 79868 169594 79870
rect 169707 79867 169773 79870
rect 169886 79868 169892 79932
rect 169956 79930 169962 79932
rect 169956 79870 170014 79930
rect 169956 79868 169962 79870
rect 170438 79868 170444 79932
rect 170508 79930 170514 79932
rect 170806 79930 170812 79932
rect 170508 79870 170566 79930
rect 170720 79870 170812 79930
rect 170508 79868 170514 79870
rect 170806 79868 170812 79870
rect 170876 79868 170882 79932
rect 171174 79930 171180 79932
rect 171088 79870 171180 79930
rect 171174 79868 171180 79870
rect 171244 79868 171250 79932
rect 171455 79906 171460 79962
rect 171516 79906 171521 79962
rect 173755 79962 173821 79967
rect 171731 79932 171797 79933
rect 171915 79932 171981 79933
rect 172191 79932 172257 79933
rect 172467 79932 172533 79933
rect 171726 79930 171732 79932
rect 171455 79901 171521 79906
rect 171640 79870 171732 79930
rect 171726 79868 171732 79870
rect 171796 79868 171802 79932
rect 171910 79868 171916 79932
rect 171980 79930 171986 79932
rect 171980 79870 172072 79930
rect 171980 79868 171986 79870
rect 172140 79868 172146 79932
rect 172210 79930 172257 79932
rect 172210 79928 172302 79930
rect 172252 79872 172302 79928
rect 172210 79870 172302 79872
rect 172210 79868 172257 79870
rect 172462 79868 172468 79932
rect 172532 79930 172538 79932
rect 172532 79870 172624 79930
rect 173203 79928 173269 79933
rect 173755 79932 173760 79962
rect 173816 79932 173821 79962
rect 173939 79962 174005 79967
rect 173203 79872 173208 79928
rect 173264 79872 173269 79928
rect 172532 79868 172538 79870
rect 170811 79867 170877 79868
rect 171179 79867 171245 79868
rect 171731 79867 171797 79868
rect 171915 79867 171981 79868
rect 172191 79867 172257 79868
rect 172467 79867 172533 79868
rect 173203 79867 173269 79872
rect 173750 79868 173756 79932
rect 173820 79930 173826 79932
rect 173820 79870 173878 79930
rect 173939 79906 173944 79962
rect 174000 79906 174005 79962
rect 173939 79901 174005 79906
rect 173820 79868 173826 79870
rect 173206 79794 173266 79867
rect 173942 79796 174002 79901
rect 168652 79734 173266 79794
rect 173934 79732 173940 79796
rect 174004 79732 174010 79796
rect 166717 79658 166783 79661
rect 166582 79656 166783 79658
rect 166582 79600 166722 79656
rect 166778 79600 166783 79656
rect 166582 79598 166783 79600
rect 164969 79595 165035 79596
rect 166073 79595 166139 79598
rect 166717 79595 166783 79598
rect 167177 79656 167243 79661
rect 167177 79600 167182 79656
rect 167238 79600 167243 79656
rect 167177 79595 167243 79600
rect 167678 79596 167684 79660
rect 167748 79658 167754 79660
rect 168330 79658 168390 79731
rect 172830 79658 172836 79660
rect 167748 79598 168390 79658
rect 168790 79598 172836 79658
rect 167748 79596 167754 79598
rect 43437 79522 43503 79525
rect 168790 79522 168850 79598
rect 172830 79596 172836 79598
rect 172900 79596 172906 79660
rect 173065 79658 173131 79661
rect 180750 79658 180810 80006
rect 462313 80003 462379 80006
rect 173065 79656 180810 79658
rect 173065 79600 173070 79656
rect 173126 79600 180810 79656
rect 173065 79598 180810 79600
rect 173065 79595 173131 79598
rect 43437 79520 168850 79522
rect 43437 79464 43442 79520
rect 43498 79464 168850 79520
rect 43437 79462 168850 79464
rect 170397 79522 170463 79525
rect 173934 79522 173940 79524
rect 170397 79520 173940 79522
rect 170397 79464 170402 79520
rect 170458 79464 173940 79520
rect 170397 79462 173940 79464
rect 43437 79459 43503 79462
rect 170397 79459 170463 79462
rect 173934 79460 173940 79462
rect 174004 79460 174010 79524
rect 37917 79386 37983 79389
rect 165613 79386 165679 79389
rect 37917 79384 165679 79386
rect 37917 79328 37922 79384
rect 37978 79328 165618 79384
rect 165674 79328 165679 79384
rect 37917 79326 165679 79328
rect 37917 79323 37983 79326
rect 165613 79323 165679 79326
rect 166073 79386 166139 79389
rect 166390 79386 166396 79388
rect 166073 79384 166396 79386
rect 166073 79328 166078 79384
rect 166134 79328 166396 79384
rect 166073 79326 166396 79328
rect 166073 79323 166139 79326
rect 166390 79324 166396 79326
rect 166460 79324 166466 79388
rect 167310 79324 167316 79388
rect 167380 79386 167386 79388
rect 167545 79386 167611 79389
rect 167380 79384 167611 79386
rect 167380 79328 167550 79384
rect 167606 79328 167611 79384
rect 167380 79326 167611 79328
rect 167380 79324 167386 79326
rect 167545 79323 167611 79326
rect 167862 79324 167868 79388
rect 167932 79386 167938 79388
rect 168005 79386 168071 79389
rect 167932 79384 168071 79386
rect 167932 79328 168010 79384
rect 168066 79328 168071 79384
rect 167932 79326 168071 79328
rect 167932 79324 167938 79326
rect 168005 79323 168071 79326
rect 168649 79386 168715 79389
rect 168925 79388 168991 79389
rect 169845 79388 169911 79389
rect 168782 79386 168788 79388
rect 168649 79384 168788 79386
rect 168649 79328 168654 79384
rect 168710 79328 168788 79384
rect 168649 79326 168788 79328
rect 168649 79323 168715 79326
rect 168782 79324 168788 79326
rect 168852 79324 168858 79388
rect 168925 79384 168972 79388
rect 169036 79386 169042 79388
rect 169845 79386 169892 79388
rect 168925 79328 168930 79384
rect 168925 79324 168972 79328
rect 169036 79326 169082 79386
rect 169800 79384 169892 79386
rect 169800 79328 169850 79384
rect 169800 79326 169892 79328
rect 169036 79324 169042 79326
rect 169845 79324 169892 79326
rect 169956 79324 169962 79388
rect 170254 79324 170260 79388
rect 170324 79386 170330 79388
rect 170489 79386 170555 79389
rect 170324 79384 170555 79386
rect 170324 79328 170494 79384
rect 170550 79328 170555 79384
rect 170324 79326 170555 79328
rect 170324 79324 170330 79326
rect 168925 79323 168991 79324
rect 169845 79323 169911 79324
rect 170489 79323 170555 79326
rect 171174 79324 171180 79388
rect 171244 79386 171250 79388
rect 171777 79386 171843 79389
rect 171244 79384 171843 79386
rect 171244 79328 171782 79384
rect 171838 79328 171843 79384
rect 171244 79326 171843 79328
rect 171244 79324 171250 79326
rect 171777 79323 171843 79326
rect 172421 79386 172487 79389
rect 173065 79386 173131 79389
rect 172421 79384 173131 79386
rect 172421 79328 172426 79384
rect 172482 79328 173070 79384
rect 173126 79328 173131 79384
rect 172421 79326 173131 79328
rect 172421 79323 172487 79326
rect 173065 79323 173131 79326
rect 173198 79324 173204 79388
rect 173268 79386 173274 79388
rect 173341 79386 173407 79389
rect 173268 79384 173407 79386
rect 173268 79328 173346 79384
rect 173402 79328 173407 79384
rect 173268 79326 173407 79328
rect 173268 79324 173274 79326
rect 173341 79323 173407 79326
rect 6913 79250 6979 79253
rect 165981 79250 166047 79253
rect 6913 79248 166047 79250
rect 6913 79192 6918 79248
rect 6974 79192 165986 79248
rect 166042 79192 166047 79248
rect 6913 79190 166047 79192
rect 6913 79187 6979 79190
rect 165981 79187 166047 79190
rect 166257 79250 166323 79253
rect 172881 79250 172947 79253
rect 166257 79248 172947 79250
rect 166257 79192 166262 79248
rect 166318 79192 172886 79248
rect 172942 79192 172947 79248
rect 166257 79190 172947 79192
rect 166257 79187 166323 79190
rect 172881 79187 172947 79190
rect 173341 79250 173407 79253
rect 173750 79250 173756 79252
rect 173341 79248 173756 79250
rect 173341 79192 173346 79248
rect 173402 79192 173756 79248
rect 173341 79190 173756 79192
rect 173341 79187 173407 79190
rect 173750 79188 173756 79190
rect 173820 79188 173826 79252
rect 3785 79114 3851 79117
rect 162393 79114 162459 79117
rect 162526 79114 162532 79116
rect 3785 79112 162226 79114
rect 3785 79056 3790 79112
rect 3846 79056 162226 79112
rect 3785 79054 162226 79056
rect 3785 79051 3851 79054
rect 3601 78978 3667 78981
rect 161974 78978 161980 78980
rect 3601 78976 161980 78978
rect 3601 78920 3606 78976
rect 3662 78920 161980 78976
rect 3601 78918 161980 78920
rect 3601 78915 3667 78918
rect 161974 78916 161980 78918
rect 162044 78916 162050 78980
rect 162166 78978 162226 79054
rect 162393 79112 162532 79114
rect 162393 79056 162398 79112
rect 162454 79056 162532 79112
rect 162393 79054 162532 79056
rect 162393 79051 162459 79054
rect 162526 79052 162532 79054
rect 162596 79052 162602 79116
rect 165613 79114 165679 79117
rect 173433 79114 173499 79117
rect 165613 79112 173499 79114
rect 165613 79056 165618 79112
rect 165674 79056 173438 79112
rect 173494 79056 173499 79112
rect 165613 79054 173499 79056
rect 165613 79051 165679 79054
rect 173433 79051 173499 79054
rect 173525 78978 173591 78981
rect 162166 78976 173591 78978
rect 162166 78920 173530 78976
rect 173586 78920 173591 78976
rect 162166 78918 173591 78920
rect 173525 78915 173591 78918
rect 3417 78842 3483 78845
rect 173249 78842 173315 78845
rect 3417 78840 173315 78842
rect 3417 78784 3422 78840
rect 3478 78784 173254 78840
rect 173310 78784 173315 78840
rect 3417 78782 173315 78784
rect 3417 78779 3483 78782
rect 173249 78779 173315 78782
rect 133270 78644 133276 78708
rect 133340 78706 133346 78708
rect 133597 78706 133663 78709
rect 133340 78704 133663 78706
rect 133340 78648 133602 78704
rect 133658 78648 133663 78704
rect 133340 78646 133663 78648
rect 133340 78644 133346 78646
rect 133597 78643 133663 78646
rect 134006 78644 134012 78708
rect 134076 78706 134082 78708
rect 134241 78706 134307 78709
rect 136909 78708 136975 78709
rect 138013 78708 138079 78709
rect 136909 78706 136956 78708
rect 134076 78704 134307 78706
rect 134076 78648 134246 78704
rect 134302 78648 134307 78704
rect 134076 78646 134307 78648
rect 136864 78704 136956 78706
rect 136864 78648 136914 78704
rect 136864 78646 136956 78648
rect 134076 78644 134082 78646
rect 134241 78643 134307 78646
rect 136909 78644 136956 78646
rect 137020 78644 137026 78708
rect 138013 78706 138060 78708
rect 137968 78704 138060 78706
rect 137968 78648 138018 78704
rect 137968 78646 138060 78648
rect 138013 78644 138060 78646
rect 138124 78644 138130 78708
rect 140446 78644 140452 78708
rect 140516 78706 140522 78708
rect 140773 78706 140839 78709
rect 140516 78704 140839 78706
rect 140516 78648 140778 78704
rect 140834 78648 140839 78704
rect 140516 78646 140839 78648
rect 140516 78644 140522 78646
rect 136909 78643 136975 78644
rect 138013 78643 138079 78644
rect 140773 78643 140839 78646
rect 143349 78708 143415 78709
rect 143349 78704 143396 78708
rect 143460 78706 143466 78708
rect 143901 78706 143967 78709
rect 144310 78706 144316 78708
rect 143349 78648 143354 78704
rect 143349 78644 143396 78648
rect 143460 78646 143506 78706
rect 143901 78704 144316 78706
rect 143901 78648 143906 78704
rect 143962 78648 144316 78704
rect 143901 78646 144316 78648
rect 143460 78644 143466 78646
rect 143349 78643 143415 78644
rect 143901 78643 143967 78646
rect 144310 78644 144316 78646
rect 144380 78644 144386 78708
rect 145097 78706 145163 78709
rect 145782 78706 145788 78708
rect 145097 78704 145788 78706
rect 145097 78648 145102 78704
rect 145158 78648 145788 78704
rect 145097 78646 145788 78648
rect 145097 78643 145163 78646
rect 145782 78644 145788 78646
rect 145852 78644 145858 78708
rect 146017 78706 146083 78709
rect 146150 78706 146156 78708
rect 146017 78704 146156 78706
rect 146017 78648 146022 78704
rect 146078 78648 146156 78704
rect 146017 78646 146156 78648
rect 146017 78643 146083 78646
rect 146150 78644 146156 78646
rect 146220 78644 146226 78708
rect 151302 78644 151308 78708
rect 151372 78706 151378 78708
rect 151629 78706 151695 78709
rect 151372 78704 151695 78706
rect 151372 78648 151634 78704
rect 151690 78648 151695 78704
rect 151372 78646 151695 78648
rect 151372 78644 151378 78646
rect 151629 78643 151695 78646
rect 152825 78706 152891 78709
rect 156321 78708 156387 78709
rect 152958 78706 152964 78708
rect 152825 78704 152964 78706
rect 152825 78648 152830 78704
rect 152886 78648 152964 78704
rect 152825 78646 152964 78648
rect 152825 78643 152891 78646
rect 152958 78644 152964 78646
rect 153028 78644 153034 78708
rect 156270 78644 156276 78708
rect 156340 78706 156387 78708
rect 156340 78704 156432 78706
rect 156382 78648 156432 78704
rect 156340 78646 156432 78648
rect 156340 78644 156387 78646
rect 156638 78644 156644 78708
rect 156708 78706 156714 78708
rect 157149 78706 157215 78709
rect 156708 78704 157215 78706
rect 156708 78648 157154 78704
rect 157210 78648 157215 78704
rect 156708 78646 157215 78648
rect 156708 78644 156714 78646
rect 156321 78643 156387 78644
rect 157149 78643 157215 78646
rect 159357 78706 159423 78709
rect 159950 78706 159956 78708
rect 159357 78704 159956 78706
rect 159357 78648 159362 78704
rect 159418 78648 159956 78704
rect 159357 78646 159956 78648
rect 159357 78643 159423 78646
rect 159950 78644 159956 78646
rect 160020 78644 160026 78708
rect 162710 78644 162716 78708
rect 162780 78706 162786 78708
rect 164785 78706 164851 78709
rect 162780 78704 164851 78706
rect 162780 78648 164790 78704
rect 164846 78648 164851 78704
rect 162780 78646 164851 78648
rect 162780 78644 162786 78646
rect 164785 78643 164851 78646
rect 164969 78706 165035 78709
rect 165153 78706 165219 78709
rect 164969 78704 165219 78706
rect 164969 78648 164974 78704
rect 165030 78648 165158 78704
rect 165214 78648 165219 78704
rect 164969 78646 165219 78648
rect 164969 78643 165035 78646
rect 165153 78643 165219 78646
rect 166993 78706 167059 78709
rect 167177 78706 167243 78709
rect 168005 78708 168071 78709
rect 168005 78706 168052 78708
rect 166993 78704 167243 78706
rect 166993 78648 166998 78704
rect 167054 78648 167182 78704
rect 167238 78648 167243 78704
rect 166993 78646 167243 78648
rect 167960 78704 168052 78706
rect 167960 78648 168010 78704
rect 167960 78646 168052 78648
rect 166993 78643 167059 78646
rect 167177 78643 167243 78646
rect 168005 78644 168052 78646
rect 168116 78644 168122 78708
rect 170581 78706 170647 78709
rect 170990 78706 170996 78708
rect 170581 78704 170996 78706
rect 170581 78648 170586 78704
rect 170642 78648 170996 78704
rect 170581 78646 170996 78648
rect 168005 78643 168071 78644
rect 170581 78643 170647 78646
rect 170990 78644 170996 78646
rect 171060 78644 171066 78708
rect 171317 78706 171383 78709
rect 172278 78706 172284 78708
rect 171317 78704 172284 78706
rect 171317 78648 171322 78704
rect 171378 78648 172284 78704
rect 171317 78646 172284 78648
rect 171317 78643 171383 78646
rect 172278 78644 172284 78646
rect 172348 78644 172354 78708
rect 172462 78644 172468 78708
rect 172532 78706 172538 78708
rect 397453 78706 397519 78709
rect 172532 78704 397519 78706
rect 172532 78648 397458 78704
rect 397514 78648 397519 78704
rect 172532 78646 397519 78648
rect 172532 78644 172538 78646
rect 397453 78643 397519 78646
rect 4889 78570 4955 78573
rect 165981 78570 166047 78573
rect 4889 78568 166047 78570
rect 4889 78512 4894 78568
rect 4950 78512 165986 78568
rect 166042 78512 166047 78568
rect 4889 78510 166047 78512
rect 4889 78507 4955 78510
rect 165981 78507 166047 78510
rect 166950 78510 171794 78570
rect 132585 78434 132651 78437
rect 151721 78436 151787 78437
rect 133270 78434 133276 78436
rect 132585 78432 133276 78434
rect 132585 78376 132590 78432
rect 132646 78376 133276 78432
rect 132585 78374 133276 78376
rect 132585 78371 132651 78374
rect 133270 78372 133276 78374
rect 133340 78372 133346 78436
rect 151670 78434 151676 78436
rect 151630 78374 151676 78434
rect 151740 78432 151787 78436
rect 151782 78376 151787 78432
rect 151670 78372 151676 78374
rect 151740 78372 151787 78376
rect 152406 78372 152412 78436
rect 152476 78434 152482 78436
rect 152733 78434 152799 78437
rect 152476 78432 152799 78434
rect 152476 78376 152738 78432
rect 152794 78376 152799 78432
rect 152476 78374 152799 78376
rect 152476 78372 152482 78374
rect 151721 78371 151787 78372
rect 152733 78371 152799 78374
rect 157374 78372 157380 78436
rect 157444 78434 157450 78436
rect 157885 78434 157951 78437
rect 157444 78432 157951 78434
rect 157444 78376 157890 78432
rect 157946 78376 157951 78432
rect 157444 78374 157951 78376
rect 157444 78372 157450 78374
rect 157885 78371 157951 78374
rect 160185 78434 160251 78437
rect 160502 78434 160508 78436
rect 160185 78432 160508 78434
rect 160185 78376 160190 78432
rect 160246 78376 160508 78432
rect 160185 78374 160508 78376
rect 160185 78371 160251 78374
rect 160502 78372 160508 78374
rect 160572 78372 160578 78436
rect 163589 78434 163655 78437
rect 166950 78434 167010 78510
rect 171542 78434 171548 78436
rect 163589 78432 167010 78434
rect 163589 78376 163594 78432
rect 163650 78376 167010 78432
rect 163589 78374 167010 78376
rect 168330 78374 171548 78434
rect 163589 78371 163655 78374
rect 126145 78298 126211 78301
rect 130878 78298 130884 78300
rect 126145 78296 130884 78298
rect 126145 78240 126150 78296
rect 126206 78240 130884 78296
rect 126145 78238 130884 78240
rect 126145 78235 126211 78238
rect 130878 78236 130884 78238
rect 130948 78236 130954 78300
rect 133086 78236 133092 78300
rect 133156 78298 133162 78300
rect 133229 78298 133295 78301
rect 133156 78296 133295 78298
rect 133156 78240 133234 78296
rect 133290 78240 133295 78296
rect 133156 78238 133295 78240
rect 133156 78236 133162 78238
rect 133229 78235 133295 78238
rect 134926 78236 134932 78300
rect 134996 78298 135002 78300
rect 138289 78298 138355 78301
rect 139209 78300 139275 78301
rect 139158 78298 139164 78300
rect 134996 78296 138355 78298
rect 134996 78240 138294 78296
rect 138350 78240 138355 78296
rect 134996 78238 138355 78240
rect 139118 78238 139164 78298
rect 139228 78296 139275 78300
rect 139270 78240 139275 78296
rect 134996 78236 135002 78238
rect 138289 78235 138355 78238
rect 139158 78236 139164 78238
rect 139228 78236 139275 78240
rect 140998 78236 141004 78300
rect 141068 78298 141074 78300
rect 141918 78298 141924 78300
rect 141068 78238 141924 78298
rect 141068 78236 141074 78238
rect 141918 78236 141924 78238
rect 141988 78236 141994 78300
rect 143022 78236 143028 78300
rect 143092 78298 143098 78300
rect 143257 78298 143323 78301
rect 143092 78296 143323 78298
rect 143092 78240 143262 78296
rect 143318 78240 143323 78296
rect 143092 78238 143323 78240
rect 143092 78236 143098 78238
rect 139209 78235 139275 78236
rect 143257 78235 143323 78238
rect 148542 78236 148548 78300
rect 148612 78298 148618 78300
rect 148777 78298 148843 78301
rect 148612 78296 148843 78298
rect 148612 78240 148782 78296
rect 148838 78240 148843 78296
rect 148612 78238 148843 78240
rect 148612 78236 148618 78238
rect 148777 78235 148843 78238
rect 159725 78298 159791 78301
rect 168330 78298 168390 78374
rect 171542 78372 171548 78374
rect 171612 78372 171618 78436
rect 168741 78300 168807 78301
rect 168741 78298 168788 78300
rect 159725 78296 168390 78298
rect 159725 78240 159730 78296
rect 159786 78240 168390 78296
rect 159725 78238 168390 78240
rect 168696 78296 168788 78298
rect 168696 78240 168746 78296
rect 168696 78238 168788 78240
rect 159725 78235 159791 78238
rect 168741 78236 168788 78238
rect 168852 78236 168858 78300
rect 170254 78236 170260 78300
rect 170324 78298 170330 78300
rect 170489 78298 170555 78301
rect 170324 78296 170555 78298
rect 170324 78240 170494 78296
rect 170550 78240 170555 78296
rect 170324 78238 170555 78240
rect 170324 78236 170330 78238
rect 168741 78235 168807 78236
rect 170489 78235 170555 78238
rect 113817 78162 113883 78165
rect 123293 78162 123359 78165
rect 113817 78160 123359 78162
rect 113817 78104 113822 78160
rect 113878 78104 123298 78160
rect 123354 78104 123359 78160
rect 113817 78102 123359 78104
rect 113817 78099 113883 78102
rect 123293 78099 123359 78102
rect 128486 78100 128492 78164
rect 128556 78162 128562 78164
rect 128721 78162 128787 78165
rect 128556 78160 128787 78162
rect 128556 78104 128726 78160
rect 128782 78104 128787 78160
rect 128556 78102 128787 78104
rect 128556 78100 128562 78102
rect 128721 78099 128787 78102
rect 132769 78162 132835 78165
rect 133086 78162 133092 78164
rect 132769 78160 133092 78162
rect 132769 78104 132774 78160
rect 132830 78104 133092 78160
rect 132769 78102 133092 78104
rect 132769 78099 132835 78102
rect 133086 78100 133092 78102
rect 133156 78100 133162 78164
rect 136398 78100 136404 78164
rect 136468 78162 136474 78164
rect 143073 78162 143139 78165
rect 136468 78160 143139 78162
rect 136468 78104 143078 78160
rect 143134 78104 143139 78160
rect 136468 78102 143139 78104
rect 136468 78100 136474 78102
rect 143073 78099 143139 78102
rect 145598 78100 145604 78164
rect 145668 78162 145674 78164
rect 146109 78162 146175 78165
rect 145668 78160 146175 78162
rect 145668 78104 146114 78160
rect 146170 78104 146175 78160
rect 145668 78102 146175 78104
rect 145668 78100 145674 78102
rect 146109 78099 146175 78102
rect 149697 78162 149763 78165
rect 149830 78162 149836 78164
rect 149697 78160 149836 78162
rect 149697 78104 149702 78160
rect 149758 78104 149836 78160
rect 149697 78102 149836 78104
rect 149697 78099 149763 78102
rect 149830 78100 149836 78102
rect 149900 78100 149906 78164
rect 150014 78100 150020 78164
rect 150084 78162 150090 78164
rect 150157 78162 150223 78165
rect 150985 78164 151051 78165
rect 150084 78160 150223 78162
rect 150084 78104 150162 78160
rect 150218 78104 150223 78160
rect 150084 78102 150223 78104
rect 150084 78100 150090 78102
rect 150157 78099 150223 78102
rect 150934 78100 150940 78164
rect 151004 78162 151051 78164
rect 151004 78160 151096 78162
rect 151046 78104 151096 78160
rect 151004 78102 151096 78104
rect 151004 78100 151051 78102
rect 154062 78100 154068 78164
rect 154132 78162 154138 78164
rect 154573 78162 154639 78165
rect 154132 78160 154639 78162
rect 154132 78104 154578 78160
rect 154634 78104 154639 78160
rect 154132 78102 154639 78104
rect 154132 78100 154138 78102
rect 150985 78099 151051 78100
rect 154573 78099 154639 78102
rect 155350 78100 155356 78164
rect 155420 78162 155426 78164
rect 159449 78162 159515 78165
rect 155420 78160 159515 78162
rect 155420 78104 159454 78160
rect 159510 78104 159515 78160
rect 155420 78102 159515 78104
rect 155420 78100 155426 78102
rect 159449 78099 159515 78102
rect 166257 78162 166323 78165
rect 168005 78162 168071 78165
rect 166257 78160 168071 78162
rect 166257 78104 166262 78160
rect 166318 78104 168010 78160
rect 168066 78104 168071 78160
rect 166257 78102 168071 78104
rect 166257 78099 166323 78102
rect 168005 78099 168071 78102
rect 168414 78100 168420 78164
rect 168484 78162 168490 78164
rect 170581 78162 170647 78165
rect 168484 78160 170647 78162
rect 168484 78104 170586 78160
rect 170642 78104 170647 78160
rect 168484 78102 170647 78104
rect 168484 78100 168490 78102
rect 170581 78099 170647 78102
rect 124121 78026 124187 78029
rect 149237 78026 149303 78029
rect 124121 78024 149303 78026
rect 124121 77968 124126 78024
rect 124182 77968 149242 78024
rect 149298 77968 149303 78024
rect 124121 77966 149303 77968
rect 124121 77963 124187 77966
rect 149237 77963 149303 77966
rect 153878 77964 153884 78028
rect 153948 78026 153954 78028
rect 154297 78026 154363 78029
rect 153948 78024 154363 78026
rect 153948 77968 154302 78024
rect 154358 77968 154363 78024
rect 153948 77966 154363 77968
rect 153948 77964 153954 77966
rect 154297 77963 154363 77966
rect 154614 77964 154620 78028
rect 154684 78026 154690 78028
rect 171225 78026 171291 78029
rect 154684 78024 171291 78026
rect 154684 77968 171230 78024
rect 171286 77968 171291 78024
rect 154684 77966 171291 77968
rect 171734 78026 171794 78510
rect 171910 78508 171916 78572
rect 171980 78570 171986 78572
rect 179413 78570 179479 78573
rect 171980 78568 179479 78570
rect 171980 78512 179418 78568
rect 179474 78512 179479 78568
rect 171980 78510 179479 78512
rect 171980 78508 171986 78510
rect 179413 78507 179479 78510
rect 171961 78298 172027 78301
rect 184933 78298 184999 78301
rect 171961 78296 184999 78298
rect 171961 78240 171966 78296
rect 172022 78240 184938 78296
rect 184994 78240 184999 78296
rect 171961 78238 184999 78240
rect 171961 78235 172027 78238
rect 184933 78235 184999 78238
rect 172094 78100 172100 78164
rect 172164 78162 172170 78164
rect 396574 78162 396580 78164
rect 172164 78102 396580 78162
rect 172164 78100 172170 78102
rect 396574 78100 396580 78102
rect 396644 78100 396650 78164
rect 171734 77966 176670 78026
rect 154684 77964 154690 77966
rect 171225 77963 171291 77966
rect 17217 77890 17283 77893
rect 126053 77890 126119 77893
rect 17217 77888 126119 77890
rect 17217 77832 17222 77888
rect 17278 77832 126058 77888
rect 126114 77832 126119 77888
rect 17217 77830 126119 77832
rect 17217 77827 17283 77830
rect 126053 77827 126119 77830
rect 131982 77828 131988 77892
rect 132052 77890 132058 77892
rect 136541 77890 136607 77893
rect 132052 77888 136607 77890
rect 132052 77832 136546 77888
rect 136602 77832 136607 77888
rect 132052 77830 136607 77832
rect 132052 77828 132058 77830
rect 136541 77827 136607 77830
rect 137277 77890 137343 77893
rect 146845 77890 146911 77893
rect 137277 77888 146911 77890
rect 137277 77832 137282 77888
rect 137338 77832 146850 77888
rect 146906 77832 146911 77888
rect 137277 77830 146911 77832
rect 137277 77827 137343 77830
rect 146845 77827 146911 77830
rect 148358 77828 148364 77892
rect 148428 77890 148434 77892
rect 148961 77890 149027 77893
rect 148428 77888 149027 77890
rect 148428 77832 148966 77888
rect 149022 77832 149027 77888
rect 148428 77830 149027 77832
rect 148428 77828 148434 77830
rect 148961 77827 149027 77830
rect 149830 77828 149836 77892
rect 149900 77890 149906 77892
rect 150249 77890 150315 77893
rect 149900 77888 150315 77890
rect 149900 77832 150254 77888
rect 150310 77832 150315 77888
rect 149900 77830 150315 77832
rect 149900 77828 149906 77830
rect 150249 77827 150315 77830
rect 153694 77828 153700 77892
rect 153764 77890 153770 77892
rect 155309 77890 155375 77893
rect 153764 77888 155375 77890
rect 153764 77832 155314 77888
rect 155370 77832 155375 77888
rect 153764 77830 155375 77832
rect 153764 77828 153770 77830
rect 155309 77827 155375 77830
rect 155534 77828 155540 77892
rect 155604 77890 155610 77892
rect 155677 77890 155743 77893
rect 155604 77888 155743 77890
rect 155604 77832 155682 77888
rect 155738 77832 155743 77888
rect 155604 77830 155743 77832
rect 155604 77828 155610 77830
rect 155677 77827 155743 77830
rect 157057 77890 157123 77893
rect 165981 77890 166047 77893
rect 157057 77888 166047 77890
rect 157057 77832 157062 77888
rect 157118 77832 165986 77888
rect 166042 77832 166047 77888
rect 157057 77830 166047 77832
rect 157057 77827 157123 77830
rect 165981 77827 166047 77830
rect 166206 77828 166212 77892
rect 166276 77890 166282 77892
rect 166901 77890 166967 77893
rect 172053 77890 172119 77893
rect 166276 77888 166967 77890
rect 166276 77832 166906 77888
rect 166962 77832 166967 77888
rect 166276 77830 166967 77832
rect 166276 77828 166282 77830
rect 166901 77827 166967 77830
rect 167318 77888 172119 77890
rect 167318 77832 172058 77888
rect 172114 77832 172119 77888
rect 167318 77830 172119 77832
rect 176610 77890 176670 77966
rect 483013 77890 483079 77893
rect 176610 77888 483079 77890
rect 176610 77832 483018 77888
rect 483074 77832 483079 77888
rect 176610 77830 483079 77832
rect 140262 77692 140268 77756
rect 140332 77754 140338 77756
rect 140497 77754 140563 77757
rect 140332 77752 140563 77754
rect 140332 77696 140502 77752
rect 140558 77696 140563 77752
rect 140332 77694 140563 77696
rect 140332 77692 140338 77694
rect 140497 77691 140563 77694
rect 120901 77618 120967 77621
rect 129038 77618 129044 77620
rect 120901 77616 129044 77618
rect 120901 77560 120906 77616
rect 120962 77560 129044 77616
rect 120901 77558 129044 77560
rect 120901 77555 120967 77558
rect 129038 77556 129044 77558
rect 129108 77556 129114 77620
rect 130878 77556 130884 77620
rect 130948 77618 130954 77620
rect 137277 77618 137343 77621
rect 130948 77616 137343 77618
rect 130948 77560 137282 77616
rect 137338 77560 137343 77616
rect 130948 77558 137343 77560
rect 130948 77556 130954 77558
rect 137277 77555 137343 77558
rect 158662 77556 158668 77620
rect 158732 77618 158738 77620
rect 164417 77618 164483 77621
rect 158732 77616 164483 77618
rect 158732 77560 164422 77616
rect 164478 77560 164483 77616
rect 158732 77558 164483 77560
rect 158732 77556 158738 77558
rect 164417 77555 164483 77558
rect 165981 77618 166047 77621
rect 167318 77618 167378 77830
rect 172053 77827 172119 77830
rect 483013 77827 483079 77830
rect 171726 77692 171732 77756
rect 171796 77754 171802 77756
rect 172789 77754 172855 77757
rect 171796 77752 172855 77754
rect 171796 77696 172794 77752
rect 172850 77696 172855 77752
rect 171796 77694 172855 77696
rect 171796 77692 171802 77694
rect 172789 77691 172855 77694
rect 172278 77618 172284 77620
rect 165981 77616 167378 77618
rect 165981 77560 165986 77616
rect 166042 77560 167378 77616
rect 165981 77558 167378 77560
rect 168422 77558 172284 77618
rect 165981 77555 166047 77558
rect 140589 77484 140655 77485
rect 152733 77484 152799 77485
rect 140589 77480 140636 77484
rect 140700 77482 140706 77484
rect 152733 77482 152780 77484
rect 140589 77424 140594 77480
rect 140589 77420 140636 77424
rect 140700 77422 140746 77482
rect 152688 77480 152780 77482
rect 152688 77424 152738 77480
rect 152688 77422 152780 77424
rect 140700 77420 140706 77422
rect 152733 77420 152780 77422
rect 152844 77420 152850 77484
rect 157926 77420 157932 77484
rect 157996 77482 158002 77484
rect 161105 77482 161171 77485
rect 157996 77480 161171 77482
rect 157996 77424 161110 77480
rect 161166 77424 161171 77480
rect 157996 77422 161171 77424
rect 157996 77420 158002 77422
rect 140589 77419 140655 77420
rect 152733 77419 152799 77420
rect 161105 77419 161171 77422
rect 166390 77420 166396 77484
rect 166460 77482 166466 77484
rect 166625 77482 166691 77485
rect 166460 77480 166691 77482
rect 166460 77424 166630 77480
rect 166686 77424 166691 77480
rect 166460 77422 166691 77424
rect 166460 77420 166466 77422
rect 166625 77419 166691 77422
rect 129641 77346 129707 77349
rect 131389 77348 131455 77349
rect 129958 77346 129964 77348
rect 129641 77344 129964 77346
rect 129641 77288 129646 77344
rect 129702 77288 129964 77344
rect 129641 77286 129964 77288
rect 129641 77283 129707 77286
rect 129958 77284 129964 77286
rect 130028 77284 130034 77348
rect 131389 77344 131436 77348
rect 131500 77346 131506 77348
rect 135253 77346 135319 77349
rect 135478 77346 135484 77348
rect 131389 77288 131394 77344
rect 131389 77284 131436 77288
rect 131500 77286 131546 77346
rect 135253 77344 135484 77346
rect 135253 77288 135258 77344
rect 135314 77288 135484 77344
rect 135253 77286 135484 77288
rect 131500 77284 131506 77286
rect 131389 77283 131455 77284
rect 135253 77283 135319 77286
rect 135478 77284 135484 77286
rect 135548 77284 135554 77348
rect 166574 77284 166580 77348
rect 166644 77346 166650 77348
rect 166809 77346 166875 77349
rect 166644 77344 166875 77346
rect 166644 77288 166814 77344
rect 166870 77288 166875 77344
rect 166644 77286 166875 77288
rect 166644 77284 166650 77286
rect 166809 77283 166875 77286
rect 131062 77148 131068 77212
rect 131132 77210 131138 77212
rect 131297 77210 131363 77213
rect 131132 77208 131363 77210
rect 131132 77152 131302 77208
rect 131358 77152 131363 77208
rect 131132 77150 131363 77152
rect 131132 77148 131138 77150
rect 131297 77147 131363 77150
rect 132861 77210 132927 77213
rect 133638 77210 133644 77212
rect 132861 77208 133644 77210
rect 132861 77152 132866 77208
rect 132922 77152 133644 77208
rect 132861 77150 133644 77152
rect 132861 77147 132927 77150
rect 133638 77148 133644 77150
rect 133708 77148 133714 77212
rect 152038 77148 152044 77212
rect 152108 77210 152114 77212
rect 152181 77210 152247 77213
rect 152108 77208 152247 77210
rect 152108 77152 152186 77208
rect 152242 77152 152247 77208
rect 152108 77150 152247 77152
rect 152108 77148 152114 77150
rect 152181 77147 152247 77150
rect 152774 77148 152780 77212
rect 152844 77210 152850 77212
rect 152917 77210 152983 77213
rect 152844 77208 152983 77210
rect 152844 77152 152922 77208
rect 152978 77152 152983 77208
rect 152844 77150 152983 77152
rect 152844 77148 152850 77150
rect 152917 77147 152983 77150
rect 157926 77148 157932 77212
rect 157996 77210 158002 77212
rect 158989 77210 159055 77213
rect 157996 77208 159055 77210
rect 157996 77152 158994 77208
rect 159050 77152 159055 77208
rect 157996 77150 159055 77152
rect 157996 77148 158002 77150
rect 158989 77147 159055 77150
rect 161197 77210 161263 77213
rect 168422 77210 168482 77558
rect 172278 77556 172284 77558
rect 172348 77556 172354 77620
rect 170305 77482 170371 77485
rect 170622 77482 170628 77484
rect 170305 77480 170628 77482
rect 170305 77424 170310 77480
rect 170366 77424 170628 77480
rect 170305 77422 170628 77424
rect 170305 77419 170371 77422
rect 170622 77420 170628 77422
rect 170692 77420 170698 77484
rect 161197 77208 168482 77210
rect 161197 77152 161202 77208
rect 161258 77152 168482 77208
rect 161197 77150 168482 77152
rect 172329 77210 172395 77213
rect 527173 77210 527239 77213
rect 172329 77208 527239 77210
rect 172329 77152 172334 77208
rect 172390 77152 527178 77208
rect 527234 77152 527239 77208
rect 172329 77150 527239 77152
rect 161197 77147 161263 77150
rect 172329 77147 172395 77150
rect 527173 77147 527239 77150
rect 142286 77012 142292 77076
rect 142356 77074 142362 77076
rect 211153 77074 211219 77077
rect 142356 77072 211219 77074
rect 142356 77016 211158 77072
rect 211214 77016 211219 77072
rect 142356 77014 211219 77016
rect 142356 77012 142362 77014
rect 211153 77011 211219 77014
rect 144729 76938 144795 76941
rect 247033 76938 247099 76941
rect 144729 76936 247099 76938
rect 144729 76880 144734 76936
rect 144790 76880 247038 76936
rect 247094 76880 247099 76936
rect 144729 76878 247099 76880
rect 144729 76875 144795 76878
rect 247033 76875 247099 76878
rect 111793 76802 111859 76805
rect 134149 76802 134215 76805
rect 111793 76800 134215 76802
rect 111793 76744 111798 76800
rect 111854 76744 134154 76800
rect 134210 76744 134215 76800
rect 111793 76742 134215 76744
rect 111793 76739 111859 76742
rect 134149 76739 134215 76742
rect 142337 76802 142403 76805
rect 142838 76802 142844 76804
rect 142337 76800 142844 76802
rect 142337 76744 142342 76800
rect 142398 76744 142844 76800
rect 142337 76742 142844 76744
rect 142337 76739 142403 76742
rect 142838 76740 142844 76742
rect 142908 76740 142914 76804
rect 147581 76802 147647 76805
rect 282913 76802 282979 76805
rect 147581 76800 282979 76802
rect 147581 76744 147586 76800
rect 147642 76744 282918 76800
rect 282974 76744 282979 76800
rect 147581 76742 282979 76744
rect 147581 76739 147647 76742
rect 282913 76739 282979 76742
rect 93853 76666 93919 76669
rect 132677 76666 132743 76669
rect 93853 76664 132743 76666
rect 93853 76608 93858 76664
rect 93914 76608 132682 76664
rect 132738 76608 132743 76664
rect 93853 76606 132743 76608
rect 93853 76603 93919 76606
rect 132677 76603 132743 76606
rect 146293 76666 146359 76669
rect 146518 76666 146524 76668
rect 146293 76664 146524 76666
rect 146293 76608 146298 76664
rect 146354 76608 146524 76664
rect 146293 76606 146524 76608
rect 146293 76603 146359 76606
rect 146518 76604 146524 76606
rect 146588 76604 146594 76668
rect 147070 76604 147076 76668
rect 147140 76666 147146 76668
rect 147397 76666 147463 76669
rect 147140 76664 147463 76666
rect 147140 76608 147402 76664
rect 147458 76608 147463 76664
rect 147140 76606 147463 76608
rect 147140 76604 147146 76606
rect 147397 76603 147463 76606
rect 150341 76666 150407 76669
rect 318793 76666 318859 76669
rect 150341 76664 318859 76666
rect 150341 76608 150346 76664
rect 150402 76608 318798 76664
rect 318854 76608 318859 76664
rect 150341 76606 318859 76608
rect 150341 76603 150407 76606
rect 318793 76603 318859 76606
rect 20713 76530 20779 76533
rect 126789 76530 126855 76533
rect 20713 76528 126855 76530
rect 20713 76472 20718 76528
rect 20774 76472 126794 76528
rect 126850 76472 126855 76528
rect 20713 76470 126855 76472
rect 20713 76467 20779 76470
rect 126789 76467 126855 76470
rect 145414 76468 145420 76532
rect 145484 76530 145490 76532
rect 146201 76530 146267 76533
rect 147489 76532 147555 76533
rect 147438 76530 147444 76532
rect 145484 76528 146267 76530
rect 145484 76472 146206 76528
rect 146262 76472 146267 76528
rect 145484 76470 146267 76472
rect 147398 76470 147444 76530
rect 147508 76528 147555 76532
rect 147550 76472 147555 76528
rect 145484 76468 145490 76470
rect 146201 76467 146267 76470
rect 147438 76468 147444 76470
rect 147508 76468 147555 76472
rect 147489 76467 147555 76468
rect 147857 76530 147923 76533
rect 158989 76532 159055 76533
rect 148174 76530 148180 76532
rect 147857 76528 148180 76530
rect 147857 76472 147862 76528
rect 147918 76472 148180 76528
rect 147857 76470 148180 76472
rect 147857 76467 147923 76470
rect 148174 76468 148180 76470
rect 148244 76468 148250 76532
rect 158989 76528 159036 76532
rect 159100 76530 159106 76532
rect 169569 76530 169635 76533
rect 565813 76530 565879 76533
rect 158989 76472 158994 76528
rect 158989 76468 159036 76472
rect 159100 76470 159146 76530
rect 169569 76528 565879 76530
rect 169569 76472 169574 76528
rect 169630 76472 565818 76528
rect 565874 76472 565879 76528
rect 169569 76470 565879 76472
rect 159100 76468 159106 76470
rect 158989 76467 159055 76468
rect 169569 76467 169635 76470
rect 565813 76467 565879 76470
rect 145046 76332 145052 76396
rect 145116 76394 145122 76396
rect 145189 76394 145255 76397
rect 145116 76392 145255 76394
rect 145116 76336 145194 76392
rect 145250 76336 145255 76392
rect 145116 76334 145255 76336
rect 145116 76332 145122 76334
rect 145189 76331 145255 76334
rect 161381 76394 161447 76397
rect 173157 76394 173223 76397
rect 161381 76392 173223 76394
rect 161381 76336 161386 76392
rect 161442 76336 173162 76392
rect 173218 76336 173223 76392
rect 161381 76334 173223 76336
rect 161381 76331 161447 76334
rect 173157 76331 173223 76334
rect 127065 75986 127131 75989
rect 161565 75988 161631 75989
rect 127198 75986 127204 75988
rect 127065 75984 127204 75986
rect 127065 75928 127070 75984
rect 127126 75928 127204 75984
rect 127065 75926 127204 75928
rect 127065 75923 127131 75926
rect 127198 75924 127204 75926
rect 127268 75924 127274 75988
rect 161565 75986 161612 75988
rect 161520 75984 161612 75986
rect 161520 75928 161570 75984
rect 161520 75926 161612 75928
rect 161565 75924 161612 75926
rect 161676 75924 161682 75988
rect 165286 75924 165292 75988
rect 165356 75986 165362 75988
rect 165429 75986 165495 75989
rect 165356 75984 165495 75986
rect 165356 75928 165434 75984
rect 165490 75928 165495 75984
rect 165356 75926 165495 75928
rect 165356 75924 165362 75926
rect 161565 75923 161631 75924
rect 165429 75923 165495 75926
rect 167177 75986 167243 75989
rect 167310 75986 167316 75988
rect 167177 75984 167316 75986
rect 167177 75928 167182 75984
rect 167238 75928 167316 75984
rect 167177 75926 167316 75928
rect 167177 75923 167243 75926
rect 167310 75924 167316 75926
rect 167380 75924 167386 75988
rect 168046 75924 168052 75988
rect 168116 75986 168122 75988
rect 168189 75986 168255 75989
rect 168116 75984 168255 75986
rect 168116 75928 168194 75984
rect 168250 75928 168255 75984
rect 168116 75926 168255 75928
rect 168116 75924 168122 75926
rect 168189 75923 168255 75926
rect 170949 75986 171015 75989
rect 171726 75986 171732 75988
rect 170949 75984 171732 75986
rect 170949 75928 170954 75984
rect 171010 75928 171732 75984
rect 170949 75926 171732 75928
rect 170949 75923 171015 75926
rect 171726 75924 171732 75926
rect 171796 75924 171802 75988
rect 162945 75714 163011 75717
rect 173341 75714 173407 75717
rect 162945 75712 173407 75714
rect 162945 75656 162950 75712
rect 163006 75656 173346 75712
rect 173402 75656 173407 75712
rect 162945 75654 173407 75656
rect 162945 75651 163011 75654
rect 173341 75651 173407 75654
rect 139342 75516 139348 75580
rect 139412 75578 139418 75580
rect 176653 75578 176719 75581
rect 139412 75576 176719 75578
rect 139412 75520 176658 75576
rect 176714 75520 176719 75576
rect 139412 75518 176719 75520
rect 139412 75516 139418 75518
rect 176653 75515 176719 75518
rect 156873 75442 156939 75445
rect 402973 75442 403039 75445
rect 156873 75440 403039 75442
rect 156873 75384 156878 75440
rect 156934 75384 402978 75440
rect 403034 75384 403039 75440
rect 156873 75382 403039 75384
rect 156873 75379 156939 75382
rect 402973 75379 403039 75382
rect 159030 75244 159036 75308
rect 159100 75306 159106 75308
rect 159909 75306 159975 75309
rect 159100 75304 159975 75306
rect 159100 75248 159914 75304
rect 159970 75248 159975 75304
rect 159100 75246 159975 75248
rect 159100 75244 159106 75246
rect 159909 75243 159975 75246
rect 161473 75306 161539 75309
rect 459553 75306 459619 75309
rect 161473 75304 459619 75306
rect 161473 75248 161478 75304
rect 161534 75248 459558 75304
rect 459614 75248 459619 75304
rect 161473 75246 459619 75248
rect 161473 75243 161539 75246
rect 459553 75243 459619 75246
rect 158846 75108 158852 75172
rect 158916 75170 158922 75172
rect 159357 75170 159423 75173
rect 158916 75168 159423 75170
rect 158916 75112 159362 75168
rect 159418 75112 159423 75168
rect 158916 75110 159423 75112
rect 158916 75108 158922 75110
rect 159357 75107 159423 75110
rect 160134 75108 160140 75172
rect 160204 75170 160210 75172
rect 160829 75170 160895 75173
rect 160204 75168 160895 75170
rect 160204 75112 160834 75168
rect 160890 75112 160895 75168
rect 160204 75110 160895 75112
rect 160204 75108 160210 75110
rect 160829 75107 160895 75110
rect 164734 75108 164740 75172
rect 164804 75170 164810 75172
rect 496813 75170 496879 75173
rect 164804 75168 496879 75170
rect 164804 75112 496818 75168
rect 496874 75112 496879 75168
rect 164804 75110 496879 75112
rect 164804 75108 164810 75110
rect 496813 75107 496879 75110
rect 162158 74972 162164 75036
rect 162228 75034 162234 75036
rect 162669 75034 162735 75037
rect 162228 75032 162735 75034
rect 162228 74976 162674 75032
rect 162730 74976 162735 75032
rect 162228 74974 162735 74976
rect 162228 74972 162234 74974
rect 162669 74971 162735 74974
rect 129089 74490 129155 74493
rect 135478 74490 135484 74492
rect 129089 74488 135484 74490
rect 129089 74432 129094 74488
rect 129150 74432 135484 74488
rect 129089 74430 135484 74432
rect 129089 74427 129155 74430
rect 135478 74428 135484 74430
rect 135548 74428 135554 74492
rect 140078 74292 140084 74356
rect 140148 74354 140154 74356
rect 194593 74354 194659 74357
rect 140148 74352 194659 74354
rect 140148 74296 194598 74352
rect 194654 74296 194659 74352
rect 140148 74294 194659 74296
rect 140148 74292 140154 74294
rect 194593 74291 194659 74294
rect 37273 74218 37339 74221
rect 128445 74218 128511 74221
rect 37273 74216 128511 74218
rect 37273 74160 37278 74216
rect 37334 74160 128450 74216
rect 128506 74160 128511 74216
rect 37273 74158 128511 74160
rect 37273 74155 37339 74158
rect 128445 74155 128511 74158
rect 143390 74156 143396 74220
rect 143460 74218 143466 74220
rect 230473 74218 230539 74221
rect 143460 74216 230539 74218
rect 143460 74160 230478 74216
rect 230534 74160 230539 74216
rect 143460 74158 230539 74160
rect 143460 74156 143466 74158
rect 230473 74155 230539 74158
rect 144637 74082 144703 74085
rect 244273 74082 244339 74085
rect 144637 74080 244339 74082
rect 144637 74024 144642 74080
rect 144698 74024 244278 74080
rect 244334 74024 244339 74080
rect 144637 74022 244339 74024
rect 144637 74019 144703 74022
rect 244273 74019 244339 74022
rect 57973 73946 58039 73949
rect 122925 73946 122991 73949
rect 57973 73944 122991 73946
rect 57973 73888 57978 73944
rect 58034 73888 122930 73944
rect 122986 73888 122991 73944
rect 57973 73886 122991 73888
rect 57973 73883 58039 73886
rect 122925 73883 122991 73886
rect 148685 73946 148751 73949
rect 298093 73946 298159 73949
rect 148685 73944 298159 73946
rect 148685 73888 148690 73944
rect 148746 73888 298098 73944
rect 298154 73888 298159 73944
rect 148685 73886 298159 73888
rect 148685 73883 148751 73886
rect 298093 73883 298159 73886
rect 170990 73748 170996 73812
rect 171060 73810 171066 73812
rect 578233 73810 578299 73813
rect 171060 73808 578299 73810
rect 171060 73752 578238 73808
rect 578294 73752 578299 73808
rect 171060 73750 578299 73752
rect 171060 73748 171066 73750
rect 578233 73747 578299 73750
rect 144310 73612 144316 73676
rect 144380 73674 144386 73676
rect 144821 73674 144887 73677
rect 144380 73672 144887 73674
rect 144380 73616 144826 73672
rect 144882 73616 144887 73672
rect 144380 73614 144887 73616
rect 144380 73612 144386 73614
rect 144821 73611 144887 73614
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect 75913 72450 75979 72453
rect 131430 72450 131436 72452
rect 75913 72448 131436 72450
rect 75913 72392 75918 72448
rect 75974 72392 131436 72448
rect 75913 72390 131436 72392
rect 75913 72387 75979 72390
rect 131430 72388 131436 72390
rect 131500 72388 131506 72452
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 40033 71226 40099 71229
rect 129038 71226 129044 71228
rect 40033 71224 129044 71226
rect 40033 71168 40038 71224
rect 40094 71168 129044 71224
rect 40033 71166 129044 71168
rect 40033 71163 40099 71166
rect 129038 71164 129044 71166
rect 129108 71164 129114 71228
rect 35985 71090 36051 71093
rect 128854 71090 128860 71092
rect 35985 71088 128860 71090
rect 35985 71032 35990 71088
rect 36046 71032 128860 71088
rect 35985 71030 128860 71032
rect 35985 71027 36051 71030
rect 128854 71028 128860 71030
rect 128924 71028 128930 71092
rect 138790 71028 138796 71092
rect 138860 71090 138866 71092
rect 174445 71090 174511 71093
rect 138860 71088 174511 71090
rect 138860 71032 174450 71088
rect 174506 71032 174511 71088
rect 138860 71030 174511 71032
rect 138860 71028 138866 71030
rect 174445 71027 174511 71030
rect 73153 69594 73219 69597
rect 131246 69594 131252 69596
rect 73153 69592 131252 69594
rect 73153 69536 73158 69592
rect 73214 69536 131252 69592
rect 73153 69534 131252 69536
rect 73153 69531 73219 69534
rect 131246 69532 131252 69534
rect 131316 69532 131322 69596
rect 131757 69594 131823 69597
rect 135294 69594 135300 69596
rect 131757 69592 135300 69594
rect 131757 69536 131762 69592
rect 131818 69536 135300 69592
rect 131757 69534 135300 69536
rect 131757 69531 131823 69534
rect 135294 69532 135300 69534
rect 135364 69532 135370 69596
rect 166206 69532 166212 69596
rect 166276 69594 166282 69596
rect 529933 69594 529999 69597
rect 166276 69592 529999 69594
rect 166276 69536 529938 69592
rect 529994 69536 529999 69592
rect 166276 69534 529999 69536
rect 166276 69532 166282 69534
rect 529933 69531 529999 69534
rect 91093 68370 91159 68373
rect 133270 68370 133276 68372
rect 91093 68368 133276 68370
rect 91093 68312 91098 68368
rect 91154 68312 133276 68368
rect 91093 68310 133276 68312
rect 91093 68307 91159 68310
rect 133270 68308 133276 68310
rect 133340 68308 133346 68372
rect 55213 68234 55279 68237
rect 129958 68234 129964 68236
rect 55213 68232 129964 68234
rect 55213 68176 55218 68232
rect 55274 68176 129964 68232
rect 55213 68174 129964 68176
rect 55213 68171 55279 68174
rect 129958 68172 129964 68174
rect 130028 68172 130034 68236
rect 138974 67492 138980 67556
rect 139044 67554 139050 67556
rect 140037 67554 140103 67557
rect 139044 67552 140103 67554
rect 139044 67496 140042 67552
rect 140098 67496 140103 67552
rect 139044 67494 140103 67496
rect 139044 67492 139050 67494
rect 140037 67491 140103 67494
rect 140262 65452 140268 65516
rect 140332 65514 140338 65516
rect 193213 65514 193279 65517
rect 140332 65512 193279 65514
rect 140332 65456 193218 65512
rect 193274 65456 193279 65512
rect 140332 65454 193279 65456
rect 140332 65452 140338 65454
rect 193213 65451 193279 65454
rect 164918 64092 164924 64156
rect 164988 64154 164994 64156
rect 511993 64154 512059 64157
rect 164988 64152 512059 64154
rect 164988 64096 511998 64152
rect 512054 64096 512059 64152
rect 164988 64094 512059 64096
rect 164988 64092 164994 64094
rect 511993 64091 512059 64094
rect 151302 62868 151308 62932
rect 151372 62930 151378 62932
rect 333973 62930 334039 62933
rect 151372 62928 334039 62930
rect 151372 62872 333978 62928
rect 334034 62872 334039 62928
rect 151372 62870 334039 62872
rect 151372 62868 151378 62870
rect 333973 62867 334039 62870
rect 167494 62732 167500 62796
rect 167564 62794 167570 62796
rect 547873 62794 547939 62797
rect 167564 62792 547939 62794
rect 167564 62736 547878 62792
rect 547934 62736 547939 62792
rect 167564 62734 547939 62736
rect 167564 62732 167570 62734
rect 547873 62731 547939 62734
rect 171542 59876 171548 59940
rect 171612 59938 171618 59940
rect 440325 59938 440391 59941
rect 171612 59936 440391 59938
rect 171612 59880 440330 59936
rect 440386 59880 440391 59936
rect 171612 59878 440391 59880
rect 171612 59876 171618 59878
rect 440325 59875 440391 59878
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 143022 58516 143028 58580
rect 143092 58578 143098 58580
rect 227713 58578 227779 58581
rect 143092 58576 227779 58578
rect 143092 58520 227718 58576
rect 227774 58520 227779 58576
rect 143092 58518 227779 58520
rect 143092 58516 143098 58518
rect 227713 58515 227779 58518
rect 145230 57428 145236 57492
rect 145300 57490 145306 57492
rect 263593 57490 263659 57493
rect 145300 57488 263659 57490
rect 145300 57432 263598 57488
rect 263654 57432 263659 57488
rect 145300 57430 263659 57432
rect 145300 57428 145306 57430
rect 263593 57427 263659 57430
rect 172278 57292 172284 57356
rect 172348 57354 172354 57356
rect 449893 57354 449959 57357
rect 172348 57352 449959 57354
rect 172348 57296 449898 57352
rect 449954 57296 449959 57352
rect 172348 57294 449959 57296
rect 172348 57292 172354 57294
rect 449893 57291 449959 57294
rect 163446 57156 163452 57220
rect 163516 57218 163522 57220
rect 494053 57218 494119 57221
rect 163516 57216 494119 57218
rect 163516 57160 494058 57216
rect 494114 57160 494119 57216
rect 163516 57158 494119 57160
rect 163516 57156 163522 57158
rect 494053 57155 494119 57158
rect 148542 55796 148548 55860
rect 148612 55858 148618 55860
rect 299473 55858 299539 55861
rect 148612 55856 299539 55858
rect 148612 55800 299478 55856
rect 299534 55800 299539 55856
rect 148612 55798 299539 55800
rect 148612 55796 148618 55798
rect 299473 55795 299539 55798
rect 161054 54436 161060 54500
rect 161124 54498 161130 54500
rect 458173 54498 458239 54501
rect 161124 54496 458239 54498
rect 161124 54440 458178 54496
rect 458234 54440 458239 54496
rect 161124 54438 458239 54440
rect 161124 54436 161130 54438
rect 458173 54435 458239 54438
rect 152406 53348 152412 53412
rect 152476 53410 152482 53412
rect 351913 53410 351979 53413
rect 152476 53408 351979 53410
rect 152476 53352 351918 53408
rect 351974 53352 351979 53408
rect 152476 53350 351979 53352
rect 152476 53348 152482 53350
rect 351913 53347 351979 53350
rect 165102 53212 165108 53276
rect 165172 53274 165178 53276
rect 514845 53274 514911 53277
rect 165172 53272 514911 53274
rect 165172 53216 514850 53272
rect 514906 53216 514911 53272
rect 165172 53214 514911 53216
rect 165172 53212 165178 53214
rect 514845 53211 514911 53214
rect 170622 53076 170628 53140
rect 170692 53138 170698 53140
rect 575473 53138 575539 53141
rect 170692 53136 575539 53138
rect 170692 53080 575478 53136
rect 575534 53080 575539 53136
rect 170692 53078 575539 53080
rect 170692 53076 170698 53078
rect 575473 53075 575539 53078
rect 166390 51716 166396 51780
rect 166460 51778 166466 51780
rect 528553 51778 528619 51781
rect 166460 51776 528619 51778
rect 166460 51720 528558 51776
rect 528614 51720 528619 51776
rect 166460 51718 528619 51720
rect 166460 51716 166466 51718
rect 528553 51715 528619 51718
rect 139158 50220 139164 50284
rect 139228 50282 139234 50284
rect 160737 50282 160803 50285
rect 139228 50280 160803 50282
rect 139228 50224 160742 50280
rect 160798 50224 160803 50280
rect 139228 50222 160803 50224
rect 139228 50220 139234 50222
rect 160737 50219 160803 50222
rect 157926 48860 157932 48924
rect 157996 48922 158002 48924
rect 423673 48922 423739 48925
rect 157996 48920 423739 48922
rect 157996 48864 423678 48920
rect 423734 48864 423739 48920
rect 157996 48862 423739 48864
rect 157996 48860 158002 48862
rect 423673 48859 423739 48862
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 167678 46140 167684 46204
rect 167748 46202 167754 46204
rect 549253 46202 549319 46205
rect 167748 46200 549319 46202
rect 167748 46144 549258 46200
rect 549314 46144 549319 46200
rect 583520 46188 584960 46278
rect 167748 46142 549319 46144
rect 167748 46140 167754 46142
rect 549253 46139 549319 46142
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 137686 44780 137692 44844
rect 137756 44842 137762 44844
rect 155217 44842 155283 44845
rect 137756 44840 155283 44842
rect 137756 44784 155222 44840
rect 155278 44784 155283 44840
rect 137756 44782 155283 44784
rect 137756 44780 137762 44782
rect 155217 44779 155283 44782
rect 155534 44780 155540 44844
rect 155604 44842 155610 44844
rect 387793 44842 387859 44845
rect 155604 44840 387859 44842
rect 155604 44784 387798 44840
rect 387854 44784 387859 44840
rect 155604 44782 387859 44784
rect 155604 44780 155610 44782
rect 387793 44779 387859 44782
rect 145414 42060 145420 42124
rect 145484 42122 145490 42124
rect 266353 42122 266419 42125
rect 145484 42120 266419 42122
rect 145484 42064 266358 42120
rect 266414 42064 266419 42120
rect 145484 42062 266419 42064
rect 145484 42060 145490 42062
rect 266353 42059 266419 42062
rect 140446 40836 140452 40900
rect 140516 40898 140522 40900
rect 191833 40898 191899 40901
rect 140516 40896 191899 40898
rect 140516 40840 191838 40896
rect 191894 40840 191899 40896
rect 140516 40838 191899 40840
rect 140516 40836 140522 40838
rect 191833 40835 191899 40838
rect 144494 40700 144500 40764
rect 144564 40762 144570 40764
rect 242985 40762 243051 40765
rect 144564 40760 243051 40762
rect 144564 40704 242990 40760
rect 243046 40704 243051 40760
rect 144564 40702 243051 40704
rect 144564 40700 144570 40702
rect 242985 40699 243051 40702
rect 165286 40564 165292 40628
rect 165356 40626 165362 40628
rect 510613 40626 510679 40629
rect 165356 40624 510679 40626
rect 165356 40568 510618 40624
rect 510674 40568 510679 40624
rect 165356 40566 510679 40568
rect 165356 40564 165362 40566
rect 510613 40563 510679 40566
rect 166574 39204 166580 39268
rect 166644 39266 166650 39268
rect 531313 39266 531379 39269
rect 166644 39264 531379 39266
rect 166644 39208 531318 39264
rect 531374 39208 531379 39264
rect 166644 39206 531379 39208
rect 166644 39204 166650 39206
rect 531313 39203 531379 39206
rect 153878 37844 153884 37908
rect 153948 37906 153954 37908
rect 369853 37906 369919 37909
rect 153948 37904 369919 37906
rect 153948 37848 369858 37904
rect 369914 37848 369919 37904
rect 153948 37846 369919 37848
rect 153948 37844 153954 37846
rect 369853 37843 369919 37846
rect 19333 35186 19399 35189
rect 127198 35186 127204 35188
rect 19333 35184 127204 35186
rect 19333 35128 19338 35184
rect 19394 35128 127204 35184
rect 19333 35126 127204 35128
rect 19333 35123 19399 35126
rect 127198 35124 127204 35126
rect 127268 35124 127274 35188
rect 583520 33146 584960 33236
rect 583342 33086 584960 33146
rect 583342 33010 583402 33086
rect 583520 33010 584960 33086
rect 583342 32996 584960 33010
rect 583342 32950 583586 32996
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 171726 31724 171732 31788
rect 171796 31786 171802 31788
rect 583526 31786 583586 32950
rect 171796 31726 583586 31786
rect 171796 31724 171802 31726
rect 156822 29548 156828 29612
rect 156892 29610 156898 29612
rect 405733 29610 405799 29613
rect 156892 29608 405799 29610
rect 156892 29552 405738 29608
rect 405794 29552 405799 29608
rect 156892 29550 405799 29552
rect 156892 29548 156898 29550
rect 405733 29547 405799 29550
rect 155718 26828 155724 26892
rect 155788 26890 155794 26892
rect 386413 26890 386479 26893
rect 155788 26888 386479 26890
rect 155788 26832 386418 26888
rect 386474 26832 386479 26888
rect 155788 26830 386479 26832
rect 155788 26828 155794 26830
rect 386413 26827 386479 26830
rect 148726 25604 148732 25668
rect 148796 25666 148802 25668
rect 299565 25666 299631 25669
rect 148796 25664 299631 25666
rect 148796 25608 299570 25664
rect 299626 25608 299631 25664
rect 148796 25606 299631 25608
rect 148796 25604 148802 25606
rect 299565 25603 299631 25606
rect 166758 25468 166764 25532
rect 166828 25530 166834 25532
rect 531405 25530 531471 25533
rect 166828 25528 531471 25530
rect 166828 25472 531410 25528
rect 531466 25472 531471 25528
rect 166828 25470 531471 25472
rect 166828 25468 166834 25470
rect 531405 25467 531471 25470
rect 140630 24380 140636 24444
rect 140700 24442 140706 24444
rect 193305 24442 193371 24445
rect 140700 24440 193371 24442
rect 140700 24384 193310 24440
rect 193366 24384 193371 24440
rect 140700 24382 193371 24384
rect 140700 24380 140706 24382
rect 193305 24379 193371 24382
rect 156638 24244 156644 24308
rect 156708 24306 156714 24308
rect 407113 24306 407179 24309
rect 156708 24304 407179 24306
rect 156708 24248 407118 24304
rect 407174 24248 407179 24304
rect 156708 24246 407179 24248
rect 156708 24244 156714 24246
rect 407113 24243 407179 24246
rect 157006 24108 157012 24172
rect 157076 24170 157082 24172
rect 407205 24170 407271 24173
rect 157076 24168 407271 24170
rect 157076 24112 407210 24168
rect 407266 24112 407271 24168
rect 157076 24110 407271 24112
rect 157076 24108 157082 24110
rect 407205 24107 407271 24110
rect 158110 22612 158116 22676
rect 158180 22674 158186 22676
rect 422293 22674 422359 22677
rect 158180 22672 422359 22674
rect 158180 22616 422298 22672
rect 422354 22616 422359 22672
rect 158180 22614 422359 22616
rect 158180 22612 158186 22614
rect 422293 22611 422359 22614
rect 152590 21388 152596 21452
rect 152660 21450 152666 21452
rect 350533 21450 350599 21453
rect 152660 21448 350599 21450
rect 152660 21392 350538 21448
rect 350594 21392 350599 21448
rect 152660 21390 350599 21392
rect 152660 21388 152666 21390
rect 350533 21387 350599 21390
rect 2773 21314 2839 21317
rect 125726 21314 125732 21316
rect 2773 21312 125732 21314
rect 2773 21256 2778 21312
rect 2834 21256 125732 21312
rect 2773 21254 125732 21256
rect 2773 21251 2839 21254
rect 125726 21252 125732 21254
rect 125796 21252 125802 21316
rect 152774 21252 152780 21316
rect 152844 21314 152850 21316
rect 354673 21314 354739 21317
rect 152844 21312 354739 21314
rect 152844 21256 354678 21312
rect 354734 21256 354739 21312
rect 152844 21254 354739 21256
rect 152844 21252 152850 21254
rect 354673 21251 354739 21254
rect 144310 19892 144316 19956
rect 144380 19954 144386 19956
rect 248413 19954 248479 19957
rect 144380 19952 248479 19954
rect 144380 19896 248418 19952
rect 248474 19896 248479 19952
rect 144380 19894 248479 19896
rect 144380 19892 144386 19894
rect 248413 19891 248479 19894
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 167862 18532 167868 18596
rect 167932 18594 167938 18596
rect 546493 18594 546559 18597
rect 167932 18592 546559 18594
rect 167932 18536 546498 18592
rect 546554 18536 546559 18592
rect 167932 18534 546559 18536
rect 167932 18532 167938 18534
rect 546493 18531 546559 18534
rect 140998 17308 141004 17372
rect 141068 17370 141074 17372
rect 212533 17370 212599 17373
rect 141068 17368 212599 17370
rect 141068 17312 212538 17368
rect 212594 17312 212599 17368
rect 141068 17310 212599 17312
rect 141068 17308 141074 17310
rect 212533 17307 212599 17310
rect 149646 17172 149652 17236
rect 149716 17234 149722 17236
rect 316033 17234 316099 17237
rect 149716 17232 316099 17234
rect 149716 17176 316038 17232
rect 316094 17176 316099 17232
rect 149716 17174 316099 17176
rect 149716 17172 149722 17174
rect 316033 17171 316099 17174
rect 152958 15812 152964 15876
rect 153028 15874 153034 15876
rect 349245 15874 349311 15877
rect 153028 15872 349311 15874
rect 153028 15816 349250 15872
rect 349306 15816 349311 15872
rect 153028 15814 349311 15816
rect 153028 15812 153034 15814
rect 349245 15811 349311 15814
rect 130878 14724 130884 14788
rect 130948 14786 130954 14788
rect 284385 14786 284451 14789
rect 130948 14784 284451 14786
rect 130948 14728 284390 14784
rect 284446 14728 284451 14784
rect 130948 14726 284451 14728
rect 130948 14724 130954 14726
rect 284385 14723 284451 14726
rect 154246 14588 154252 14652
rect 154316 14650 154322 14652
rect 365805 14650 365871 14653
rect 154316 14648 365871 14650
rect 154316 14592 365810 14648
rect 365866 14592 365871 14648
rect 154316 14590 365871 14592
rect 154316 14588 154322 14590
rect 365805 14587 365871 14590
rect 154062 14452 154068 14516
rect 154132 14514 154138 14516
rect 372889 14514 372955 14517
rect 154132 14512 372955 14514
rect 154132 14456 372894 14512
rect 372950 14456 372955 14512
rect 154132 14454 372955 14456
rect 154132 14452 154138 14454
rect 372889 14451 372955 14454
rect 143206 13636 143212 13700
rect 143276 13698 143282 13700
rect 229369 13698 229435 13701
rect 143276 13696 229435 13698
rect 143276 13640 229374 13696
rect 229430 13640 229435 13696
rect 143276 13638 229435 13640
rect 143276 13636 143282 13638
rect 229369 13635 229435 13638
rect 145598 13500 145604 13564
rect 145668 13562 145674 13564
rect 264973 13562 265039 13565
rect 145668 13560 265039 13562
rect 145668 13504 264978 13560
rect 265034 13504 265039 13560
rect 145668 13502 265039 13504
rect 145668 13500 145674 13502
rect 264973 13499 265039 13502
rect 154430 13364 154436 13428
rect 154500 13426 154506 13428
rect 371233 13426 371299 13429
rect 154500 13424 371299 13426
rect 154500 13368 371238 13424
rect 371294 13368 371299 13424
rect 154500 13366 371299 13368
rect 154500 13364 154506 13366
rect 371233 13363 371299 13366
rect 160870 13228 160876 13292
rect 160940 13290 160946 13292
rect 456885 13290 456951 13293
rect 160940 13288 456951 13290
rect 160940 13232 456890 13288
rect 456946 13232 456951 13288
rect 160940 13230 456951 13232
rect 160940 13228 160946 13230
rect 456885 13227 456951 13230
rect 165470 13092 165476 13156
rect 165540 13154 165546 13156
rect 513373 13154 513439 13157
rect 165540 13152 513439 13154
rect 165540 13096 513378 13152
rect 513434 13096 513439 13152
rect 165540 13094 513439 13096
rect 165540 13092 165546 13094
rect 513373 13091 513439 13094
rect 169334 12956 169340 13020
rect 169404 13018 169410 13020
rect 567561 13018 567627 13021
rect 169404 13016 567627 13018
rect 169404 12960 567566 13016
rect 567622 12960 567627 13016
rect 169404 12958 567627 12960
rect 169404 12956 169410 12958
rect 567561 12955 567627 12958
rect 147070 12276 147076 12340
rect 147140 12338 147146 12340
rect 280705 12338 280771 12341
rect 147140 12336 280771 12338
rect 147140 12280 280710 12336
rect 280766 12280 280771 12336
rect 147140 12278 280771 12280
rect 147140 12276 147146 12278
rect 280705 12275 280771 12278
rect 149830 12140 149836 12204
rect 149900 12202 149906 12204
rect 318057 12202 318123 12205
rect 149900 12200 318123 12202
rect 149900 12144 318062 12200
rect 318118 12144 318123 12200
rect 149900 12142 318123 12144
rect 149900 12140 149906 12142
rect 318057 12139 318123 12142
rect 151486 12004 151492 12068
rect 151556 12066 151562 12068
rect 336273 12066 336339 12069
rect 151556 12064 336339 12066
rect 151556 12008 336278 12064
rect 336334 12008 336339 12064
rect 151556 12006 336339 12008
rect 151556 12004 151562 12006
rect 336273 12003 336339 12006
rect 162526 11868 162532 11932
rect 162596 11930 162602 11932
rect 474089 11930 474155 11933
rect 162596 11928 474155 11930
rect 162596 11872 474094 11928
rect 474150 11872 474155 11928
rect 162596 11870 474155 11872
rect 162596 11868 162602 11870
rect 474089 11867 474155 11870
rect 162342 11732 162348 11796
rect 162412 11794 162418 11796
rect 478137 11794 478203 11797
rect 162412 11792 478203 11794
rect 162412 11736 478142 11792
rect 478198 11736 478203 11792
rect 162412 11734 478203 11736
rect 162412 11732 162418 11734
rect 478137 11731 478203 11734
rect 170806 11596 170812 11660
rect 170876 11658 170882 11660
rect 583385 11658 583451 11661
rect 170876 11656 583451 11658
rect 170876 11600 583390 11656
rect 583446 11600 583451 11656
rect 170876 11598 583451 11600
rect 170876 11596 170882 11598
rect 583385 11595 583451 11598
rect 136214 10916 136220 10980
rect 136284 10978 136290 10980
rect 142429 10978 142495 10981
rect 136284 10976 142495 10978
rect 136284 10920 142434 10976
rect 142490 10920 142495 10976
rect 136284 10918 142495 10920
rect 136284 10916 136290 10918
rect 142429 10915 142495 10918
rect 148358 10644 148364 10708
rect 148428 10706 148434 10708
rect 301497 10706 301563 10709
rect 148428 10704 301563 10706
rect 148428 10648 301502 10704
rect 301558 10648 301563 10704
rect 148428 10646 301563 10648
rect 148428 10644 148434 10646
rect 301497 10643 301563 10646
rect 151670 10508 151676 10572
rect 151740 10570 151746 10572
rect 337009 10570 337075 10573
rect 151740 10568 337075 10570
rect 151740 10512 337014 10568
rect 337070 10512 337075 10568
rect 151740 10510 337075 10512
rect 151740 10508 151746 10510
rect 337009 10507 337075 10510
rect 114001 10434 114067 10437
rect 134006 10434 134012 10436
rect 114001 10432 134012 10434
rect 114001 10376 114006 10432
rect 114062 10376 134012 10432
rect 114001 10374 134012 10376
rect 114001 10371 114067 10374
rect 134006 10372 134012 10374
rect 134076 10372 134082 10436
rect 158846 10372 158852 10436
rect 158916 10434 158922 10436
rect 442625 10434 442691 10437
rect 158916 10432 442691 10434
rect 158916 10376 442630 10432
rect 442686 10376 442691 10432
rect 158916 10374 442691 10376
rect 158916 10372 158922 10374
rect 442625 10371 442691 10374
rect 92473 10298 92539 10301
rect 133086 10298 133092 10300
rect 92473 10296 133092 10298
rect 92473 10240 92478 10296
rect 92534 10240 133092 10296
rect 92473 10238 133092 10240
rect 92473 10235 92539 10238
rect 133086 10236 133092 10238
rect 133156 10236 133162 10300
rect 159030 10236 159036 10300
rect 159100 10298 159106 10300
rect 443361 10298 443427 10301
rect 159100 10296 443427 10298
rect 159100 10240 443366 10296
rect 443422 10240 443427 10296
rect 159100 10238 443427 10240
rect 159100 10236 159106 10238
rect 443361 10235 443427 10238
rect 74993 9210 75059 9213
rect 131062 9210 131068 9212
rect 74993 9208 131068 9210
rect 74993 9152 74998 9208
rect 75054 9152 131068 9208
rect 74993 9150 131068 9152
rect 74993 9147 75059 9150
rect 131062 9148 131068 9150
rect 131132 9148 131138 9212
rect 147254 9148 147260 9212
rect 147324 9210 147330 9212
rect 279509 9210 279575 9213
rect 147324 9208 279575 9210
rect 147324 9152 279514 9208
rect 279570 9152 279575 9208
rect 147324 9150 279575 9152
rect 147324 9148 147330 9150
rect 279509 9147 279575 9150
rect 57237 9074 57303 9077
rect 129774 9074 129780 9076
rect 57237 9072 129780 9074
rect 57237 9016 57242 9072
rect 57298 9016 129780 9072
rect 57237 9014 129780 9016
rect 57237 9011 57303 9014
rect 129774 9012 129780 9014
rect 129844 9012 129850 9076
rect 162158 9012 162164 9076
rect 162228 9074 162234 9076
rect 476941 9074 477007 9077
rect 162228 9072 477007 9074
rect 162228 9016 476946 9072
rect 477002 9016 477007 9072
rect 162228 9014 477007 9016
rect 162228 9012 162234 9014
rect 476941 9011 477007 9014
rect 41873 8938 41939 8941
rect 128670 8938 128676 8940
rect 41873 8936 128676 8938
rect 41873 8880 41878 8936
rect 41934 8880 128676 8936
rect 41873 8878 128676 8880
rect 41873 8875 41939 8878
rect 128670 8876 128676 8878
rect 128740 8876 128746 8940
rect 170438 8876 170444 8940
rect 170508 8938 170514 8940
rect 577405 8938 577471 8941
rect 170508 8936 577471 8938
rect 170508 8880 577410 8936
rect 577466 8880 577471 8936
rect 170508 8878 577471 8880
rect 170508 8876 170514 8878
rect 577405 8875 577471 8878
rect 142838 7788 142844 7852
rect 142908 7850 142914 7852
rect 227529 7850 227595 7853
rect 142908 7848 227595 7850
rect 142908 7792 227534 7848
rect 227590 7792 227595 7848
rect 142908 7790 227595 7792
rect 142908 7788 142914 7790
rect 227529 7787 227595 7790
rect 109309 7714 109375 7717
rect 133822 7714 133828 7716
rect 109309 7712 133828 7714
rect 109309 7656 109314 7712
rect 109370 7656 133828 7712
rect 109309 7654 133828 7656
rect 109309 7651 109375 7654
rect 133822 7652 133828 7654
rect 133892 7652 133898 7716
rect 158294 7652 158300 7716
rect 158364 7714 158370 7716
rect 424961 7714 425027 7717
rect 158364 7712 425027 7714
rect 158364 7656 424966 7712
rect 425022 7656 425027 7712
rect 158364 7654 425027 7656
rect 158364 7652 158370 7654
rect 424961 7651 425027 7654
rect 19425 7578 19491 7581
rect 127014 7578 127020 7580
rect 19425 7576 127020 7578
rect 19425 7520 19430 7576
rect 19486 7520 127020 7576
rect 19425 7518 127020 7520
rect 19425 7515 19491 7518
rect 127014 7516 127020 7518
rect 127084 7516 127090 7580
rect 168046 7516 168052 7580
rect 168116 7578 168122 7580
rect 549069 7578 549135 7581
rect 168116 7576 549135 7578
rect 168116 7520 549074 7576
rect 549130 7520 549135 7576
rect 168116 7518 549135 7520
rect 168116 7516 168122 7518
rect 549069 7515 549135 7518
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 147438 6292 147444 6356
rect 147508 6354 147514 6356
rect 281901 6354 281967 6357
rect 147508 6352 281967 6354
rect 147508 6296 281906 6352
rect 281962 6296 281967 6352
rect 147508 6294 281967 6296
rect 147508 6292 147514 6294
rect 281901 6291 281967 6294
rect 150014 6156 150020 6220
rect 150084 6218 150090 6220
rect 317321 6218 317387 6221
rect 150084 6216 317387 6218
rect 150084 6160 317326 6216
rect 317382 6160 317387 6216
rect 150084 6158 317387 6160
rect 150084 6156 150090 6158
rect 317321 6155 317387 6158
rect 158478 4932 158484 4996
rect 158548 4994 158554 4996
rect 421373 4994 421439 4997
rect 158548 4992 421439 4994
rect 158548 4936 421378 4992
rect 421434 4936 421439 4992
rect 158548 4934 421439 4936
rect 158548 4932 158554 4934
rect 421373 4931 421439 4934
rect 137870 4796 137876 4860
rect 137940 4858 137946 4860
rect 158897 4858 158963 4861
rect 137940 4856 158963 4858
rect 137940 4800 158902 4856
rect 158958 4800 158963 4856
rect 137940 4798 158963 4800
rect 137940 4796 137946 4798
rect 158897 4795 158963 4798
rect 163630 4796 163636 4860
rect 163700 4858 163706 4860
rect 495893 4858 495959 4861
rect 163700 4856 495959 4858
rect 163700 4800 495898 4856
rect 495954 4800 495959 4856
rect 163700 4798 495959 4800
rect 163700 4796 163706 4798
rect 495893 4795 495959 4798
rect 136398 3572 136404 3636
rect 136468 3634 136474 3636
rect 225137 3634 225203 3637
rect 136468 3632 225203 3634
rect 136468 3576 225142 3632
rect 225198 3576 225203 3632
rect 136468 3574 225203 3576
rect 136468 3572 136474 3574
rect 225137 3571 225203 3574
rect 131982 3436 131988 3500
rect 132052 3498 132058 3500
rect 246389 3498 246455 3501
rect 132052 3496 246455 3498
rect 132052 3440 246394 3496
rect 246450 3440 246455 3496
rect 132052 3438 246455 3440
rect 132052 3436 132058 3438
rect 246389 3435 246455 3438
rect 134926 3300 134932 3364
rect 134996 3362 135002 3364
rect 164877 3362 164943 3365
rect 134996 3360 164943 3362
rect 134996 3304 164882 3360
rect 164938 3304 164943 3360
rect 134996 3302 164943 3304
rect 134996 3300 135002 3302
rect 164877 3299 164943 3302
rect 173617 3362 173683 3365
rect 501781 3362 501847 3365
rect 173617 3360 501847 3362
rect 173617 3304 173622 3360
rect 173678 3304 501786 3360
rect 501842 3304 501847 3360
rect 173617 3302 501847 3304
rect 173617 3299 173683 3302
rect 501781 3299 501847 3302
<< via3 >>
rect 396580 696900 396644 696964
rect 144684 200636 144748 200700
rect 147628 199276 147692 199340
rect 147628 196420 147692 196484
rect 151308 196012 151372 196076
rect 144684 195604 144748 195668
rect 149836 195604 149900 195668
rect 143580 191744 143644 191808
rect 141740 191252 141804 191316
rect 151308 191254 151372 191318
rect 141924 190572 141988 190636
rect 149836 190632 149900 190636
rect 149836 190576 149850 190632
rect 149850 190576 149900 190632
rect 149836 190572 149900 190576
rect 140636 186900 140700 186964
rect 146156 180704 146220 180708
rect 146156 180648 146170 180704
rect 146170 180648 146220 180704
rect 146156 180644 146220 180648
rect 140452 179148 140516 179212
rect 142660 178800 142724 178804
rect 142660 178744 142666 178800
rect 142666 178744 142722 178800
rect 142722 178744 142724 178800
rect 142660 178740 142724 178744
rect 142660 176700 142724 176764
rect 142476 173844 142540 173908
rect 142292 173708 142356 173772
rect 144132 173708 144196 173772
rect 142660 173572 142724 173636
rect 142108 171260 142172 171324
rect 142108 170852 142172 170916
rect 141740 166364 141804 166428
rect 141924 166228 141988 166292
rect 142108 161528 142172 161532
rect 142108 161472 142122 161528
rect 142122 161472 142172 161528
rect 142108 161468 142172 161472
rect 142476 143380 142540 143444
rect 142660 143244 142724 143308
rect 140452 143108 140516 143172
rect 144132 142972 144196 143036
rect 146156 142836 146220 142900
rect 140636 142700 140700 142764
rect 143580 142564 143644 142628
rect 142108 142428 142172 142492
rect 142292 142156 142356 142220
rect 168052 80548 168116 80612
rect 172284 80276 172348 80340
rect 125548 79868 125612 79932
rect 128676 79928 128740 79932
rect 128676 79872 128680 79928
rect 128680 79872 128736 79928
rect 128736 79872 128740 79928
rect 128676 79868 128740 79872
rect 129044 79928 129108 79932
rect 129044 79872 129048 79928
rect 129048 79872 129104 79928
rect 129104 79872 129108 79928
rect 129044 79868 129108 79872
rect 127020 79792 127084 79796
rect 127020 79736 127024 79792
rect 127024 79736 127080 79792
rect 127080 79736 127084 79792
rect 127020 79732 127084 79736
rect 128676 79732 128740 79796
rect 129780 79868 129844 79932
rect 130884 79868 130948 79932
rect 161980 80140 162044 80204
rect 131252 79792 131316 79796
rect 131252 79736 131256 79792
rect 131256 79736 131312 79792
rect 131312 79736 131316 79792
rect 131252 79732 131316 79736
rect 133092 79868 133156 79932
rect 133276 79868 133340 79932
rect 133828 79868 133892 79932
rect 135484 79906 135488 79932
rect 135488 79906 135544 79932
rect 135544 79906 135548 79932
rect 135484 79868 135548 79906
rect 136220 79868 136284 79932
rect 137692 79868 137756 79932
rect 136956 79732 137020 79796
rect 137876 79792 137940 79796
rect 137876 79736 137926 79792
rect 137926 79736 137940 79792
rect 137876 79732 137940 79736
rect 138060 79732 138124 79796
rect 138980 79868 139044 79932
rect 139348 79928 139412 79932
rect 139348 79872 139352 79928
rect 139352 79872 139408 79928
rect 139408 79872 139412 79928
rect 139348 79868 139412 79872
rect 138796 79732 138860 79796
rect 133644 79596 133708 79660
rect 140084 79596 140148 79660
rect 142292 79868 142356 79932
rect 141924 79732 141988 79796
rect 143212 79732 143276 79796
rect 144316 79906 144320 79932
rect 144320 79906 144376 79932
rect 144376 79906 144380 79932
rect 144316 79868 144380 79906
rect 145052 79906 145056 79932
rect 145056 79906 145112 79932
rect 145112 79906 145116 79932
rect 145052 79868 145116 79906
rect 145788 79928 145852 79932
rect 145788 79872 145792 79928
rect 145792 79872 145848 79928
rect 145848 79872 145852 79928
rect 145788 79868 145852 79872
rect 146156 79868 146220 79932
rect 147260 79928 147324 79932
rect 147260 79872 147264 79928
rect 147264 79872 147320 79928
rect 147320 79872 147324 79928
rect 147260 79868 147324 79872
rect 144500 79792 144564 79796
rect 144500 79736 144504 79792
rect 144504 79736 144560 79792
rect 144560 79736 144564 79792
rect 144500 79732 144564 79736
rect 148180 79792 148244 79796
rect 148180 79736 148230 79792
rect 148230 79736 148244 79792
rect 148180 79732 148244 79736
rect 145604 79596 145668 79660
rect 146524 79596 146588 79660
rect 149836 79868 149900 79932
rect 150940 79868 151004 79932
rect 148732 79732 148796 79796
rect 149652 79732 149716 79796
rect 151492 79732 151556 79796
rect 152044 79732 152108 79796
rect 152780 79868 152844 79932
rect 153700 79868 153764 79932
rect 154436 79928 154500 79932
rect 154436 79872 154440 79928
rect 154440 79872 154496 79928
rect 154496 79872 154500 79928
rect 152596 79732 152660 79796
rect 154436 79868 154500 79872
rect 154620 79928 154684 79932
rect 154620 79872 154624 79928
rect 154624 79872 154680 79928
rect 154680 79872 154684 79928
rect 154620 79868 154684 79872
rect 154252 79732 154316 79796
rect 155356 79928 155420 79932
rect 155356 79872 155360 79928
rect 155360 79872 155416 79928
rect 155416 79872 155420 79928
rect 155356 79868 155420 79872
rect 157380 79906 157384 79932
rect 157384 79906 157440 79932
rect 157440 79906 157444 79932
rect 157380 79868 157444 79906
rect 158116 79868 158180 79932
rect 158668 79906 158672 79932
rect 158672 79906 158728 79932
rect 158728 79906 158732 79932
rect 158668 79868 158732 79906
rect 156276 79792 156340 79796
rect 156276 79736 156280 79792
rect 156280 79736 156336 79792
rect 156336 79736 156340 79792
rect 156276 79732 156340 79736
rect 155724 79596 155788 79660
rect 156828 79596 156892 79660
rect 157932 79732 157996 79796
rect 158300 79732 158364 79796
rect 160140 80004 160204 80068
rect 159956 79928 160020 79932
rect 159956 79872 159960 79928
rect 159960 79872 160016 79928
rect 160016 79872 160020 79928
rect 159956 79868 160020 79872
rect 160508 79928 160572 79932
rect 160508 79872 160512 79928
rect 160512 79872 160568 79928
rect 160568 79872 160572 79928
rect 160508 79868 160572 79872
rect 161060 79906 161064 79932
rect 161064 79906 161120 79932
rect 161120 79906 161124 79932
rect 161060 79868 161124 79906
rect 161060 79732 161124 79796
rect 162716 79868 162780 79932
rect 161796 79732 161860 79796
rect 162348 79732 162412 79796
rect 157196 79596 157260 79660
rect 158484 79596 158548 79660
rect 159036 79596 159100 79660
rect 163452 79868 163516 79932
rect 163636 79732 163700 79796
rect 165108 79868 165172 79932
rect 165476 79792 165540 79796
rect 165476 79736 165480 79792
rect 165480 79736 165536 79792
rect 165536 79736 165540 79792
rect 165476 79732 165540 79736
rect 164740 79596 164804 79660
rect 164924 79656 164988 79660
rect 164924 79600 164974 79656
rect 164974 79600 164988 79656
rect 164924 79596 164988 79600
rect 166396 79928 166460 79932
rect 166396 79872 166400 79928
rect 166400 79872 166456 79928
rect 166456 79872 166460 79928
rect 166396 79868 166460 79872
rect 166764 79868 166828 79932
rect 167868 79868 167932 79932
rect 168420 79906 168424 79932
rect 168424 79906 168480 79932
rect 168480 79906 168484 79932
rect 168420 79868 168484 79906
rect 168972 79906 168976 79932
rect 168976 79906 169032 79932
rect 169032 79906 169036 79932
rect 168972 79868 169036 79906
rect 169524 79868 169588 79932
rect 169892 79906 169896 79932
rect 169896 79906 169952 79932
rect 169952 79906 169956 79932
rect 169892 79868 169956 79906
rect 170444 79906 170448 79932
rect 170448 79906 170504 79932
rect 170504 79906 170508 79932
rect 170444 79868 170508 79906
rect 170812 79928 170876 79932
rect 170812 79872 170816 79928
rect 170816 79872 170872 79928
rect 170872 79872 170876 79928
rect 170812 79868 170876 79872
rect 171180 79928 171244 79932
rect 171180 79872 171184 79928
rect 171184 79872 171240 79928
rect 171240 79872 171244 79928
rect 171180 79868 171244 79872
rect 171732 79928 171796 79932
rect 171732 79872 171736 79928
rect 171736 79872 171792 79928
rect 171792 79872 171796 79928
rect 171732 79868 171796 79872
rect 171916 79928 171980 79932
rect 171916 79872 171920 79928
rect 171920 79872 171976 79928
rect 171976 79872 171980 79928
rect 171916 79868 171980 79872
rect 172146 79928 172210 79932
rect 172146 79872 172196 79928
rect 172196 79872 172210 79928
rect 172146 79868 172210 79872
rect 172468 79928 172532 79932
rect 172468 79872 172472 79928
rect 172472 79872 172528 79928
rect 172528 79872 172532 79928
rect 172468 79868 172532 79872
rect 173756 79906 173760 79932
rect 173760 79906 173816 79932
rect 173816 79906 173820 79932
rect 173756 79868 173820 79906
rect 173940 79732 174004 79796
rect 167684 79596 167748 79660
rect 172836 79596 172900 79660
rect 173940 79460 174004 79524
rect 166396 79324 166460 79388
rect 167316 79324 167380 79388
rect 167868 79324 167932 79388
rect 168788 79324 168852 79388
rect 168972 79384 169036 79388
rect 168972 79328 168986 79384
rect 168986 79328 169036 79384
rect 168972 79324 169036 79328
rect 169892 79384 169956 79388
rect 169892 79328 169906 79384
rect 169906 79328 169956 79384
rect 169892 79324 169956 79328
rect 170260 79324 170324 79388
rect 171180 79324 171244 79388
rect 173204 79324 173268 79388
rect 173756 79188 173820 79252
rect 161980 78916 162044 78980
rect 162532 79052 162596 79116
rect 133276 78644 133340 78708
rect 134012 78644 134076 78708
rect 136956 78704 137020 78708
rect 136956 78648 136970 78704
rect 136970 78648 137020 78704
rect 136956 78644 137020 78648
rect 138060 78704 138124 78708
rect 138060 78648 138074 78704
rect 138074 78648 138124 78704
rect 138060 78644 138124 78648
rect 140452 78644 140516 78708
rect 143396 78704 143460 78708
rect 143396 78648 143410 78704
rect 143410 78648 143460 78704
rect 143396 78644 143460 78648
rect 144316 78644 144380 78708
rect 145788 78644 145852 78708
rect 146156 78644 146220 78708
rect 151308 78644 151372 78708
rect 152964 78644 153028 78708
rect 156276 78704 156340 78708
rect 156276 78648 156326 78704
rect 156326 78648 156340 78704
rect 156276 78644 156340 78648
rect 156644 78644 156708 78708
rect 159956 78644 160020 78708
rect 162716 78644 162780 78708
rect 168052 78704 168116 78708
rect 168052 78648 168066 78704
rect 168066 78648 168116 78704
rect 168052 78644 168116 78648
rect 170996 78644 171060 78708
rect 172284 78644 172348 78708
rect 172468 78644 172532 78708
rect 133276 78372 133340 78436
rect 151676 78432 151740 78436
rect 151676 78376 151726 78432
rect 151726 78376 151740 78432
rect 151676 78372 151740 78376
rect 152412 78372 152476 78436
rect 157380 78372 157444 78436
rect 160508 78372 160572 78436
rect 130884 78236 130948 78300
rect 133092 78236 133156 78300
rect 134932 78236 134996 78300
rect 139164 78296 139228 78300
rect 139164 78240 139214 78296
rect 139214 78240 139228 78296
rect 139164 78236 139228 78240
rect 141004 78236 141068 78300
rect 141924 78236 141988 78300
rect 143028 78236 143092 78300
rect 148548 78236 148612 78300
rect 171548 78372 171612 78436
rect 168788 78296 168852 78300
rect 168788 78240 168802 78296
rect 168802 78240 168852 78296
rect 168788 78236 168852 78240
rect 170260 78236 170324 78300
rect 128492 78100 128556 78164
rect 133092 78100 133156 78164
rect 136404 78100 136468 78164
rect 145604 78100 145668 78164
rect 149836 78100 149900 78164
rect 150020 78100 150084 78164
rect 150940 78160 151004 78164
rect 150940 78104 150990 78160
rect 150990 78104 151004 78160
rect 150940 78100 151004 78104
rect 154068 78100 154132 78164
rect 155356 78100 155420 78164
rect 168420 78100 168484 78164
rect 153884 77964 153948 78028
rect 154620 77964 154684 78028
rect 171916 78508 171980 78572
rect 172100 78100 172164 78164
rect 396580 78100 396644 78164
rect 131988 77828 132052 77892
rect 148364 77828 148428 77892
rect 149836 77828 149900 77892
rect 153700 77828 153764 77892
rect 155540 77828 155604 77892
rect 166212 77828 166276 77892
rect 140268 77692 140332 77756
rect 129044 77556 129108 77620
rect 130884 77556 130948 77620
rect 158668 77556 158732 77620
rect 171732 77692 171796 77756
rect 140636 77480 140700 77484
rect 140636 77424 140650 77480
rect 140650 77424 140700 77480
rect 140636 77420 140700 77424
rect 152780 77480 152844 77484
rect 152780 77424 152794 77480
rect 152794 77424 152844 77480
rect 152780 77420 152844 77424
rect 157932 77420 157996 77484
rect 166396 77420 166460 77484
rect 129964 77284 130028 77348
rect 131436 77344 131500 77348
rect 131436 77288 131450 77344
rect 131450 77288 131500 77344
rect 131436 77284 131500 77288
rect 135484 77284 135548 77348
rect 166580 77284 166644 77348
rect 131068 77148 131132 77212
rect 133644 77148 133708 77212
rect 152044 77148 152108 77212
rect 152780 77148 152844 77212
rect 157932 77148 157996 77212
rect 172284 77556 172348 77620
rect 170628 77420 170692 77484
rect 142292 77012 142356 77076
rect 142844 76740 142908 76804
rect 146524 76604 146588 76668
rect 147076 76604 147140 76668
rect 145420 76468 145484 76532
rect 147444 76528 147508 76532
rect 147444 76472 147494 76528
rect 147494 76472 147508 76528
rect 147444 76468 147508 76472
rect 148180 76468 148244 76532
rect 159036 76528 159100 76532
rect 159036 76472 159050 76528
rect 159050 76472 159100 76528
rect 159036 76468 159100 76472
rect 145052 76332 145116 76396
rect 127204 75924 127268 75988
rect 161612 75984 161676 75988
rect 161612 75928 161626 75984
rect 161626 75928 161676 75984
rect 161612 75924 161676 75928
rect 165292 75924 165356 75988
rect 167316 75924 167380 75988
rect 168052 75924 168116 75988
rect 171732 75924 171796 75988
rect 139348 75516 139412 75580
rect 159036 75244 159100 75308
rect 158852 75108 158916 75172
rect 160140 75108 160204 75172
rect 164740 75108 164804 75172
rect 162164 74972 162228 75036
rect 135484 74428 135548 74492
rect 140084 74292 140148 74356
rect 143396 74156 143460 74220
rect 170996 73748 171060 73812
rect 144316 73612 144380 73676
rect 131436 72388 131500 72452
rect 129044 71164 129108 71228
rect 128860 71028 128924 71092
rect 138796 71028 138860 71092
rect 131252 69532 131316 69596
rect 135300 69532 135364 69596
rect 166212 69532 166276 69596
rect 133276 68308 133340 68372
rect 129964 68172 130028 68236
rect 138980 67492 139044 67556
rect 140268 65452 140332 65516
rect 164924 64092 164988 64156
rect 151308 62868 151372 62932
rect 167500 62732 167564 62796
rect 171548 59876 171612 59940
rect 143028 58516 143092 58580
rect 145236 57428 145300 57492
rect 172284 57292 172348 57356
rect 163452 57156 163516 57220
rect 148548 55796 148612 55860
rect 161060 54436 161124 54500
rect 152412 53348 152476 53412
rect 165108 53212 165172 53276
rect 170628 53076 170692 53140
rect 166396 51716 166460 51780
rect 139164 50220 139228 50284
rect 157932 48860 157996 48924
rect 167684 46140 167748 46204
rect 137692 44780 137756 44844
rect 155540 44780 155604 44844
rect 145420 42060 145484 42124
rect 140452 40836 140516 40900
rect 144500 40700 144564 40764
rect 165292 40564 165356 40628
rect 166580 39204 166644 39268
rect 153884 37844 153948 37908
rect 127204 35124 127268 35188
rect 171732 31724 171796 31788
rect 156828 29548 156892 29612
rect 155724 26828 155788 26892
rect 148732 25604 148796 25668
rect 166764 25468 166828 25532
rect 140636 24380 140700 24444
rect 156644 24244 156708 24308
rect 157012 24108 157076 24172
rect 158116 22612 158180 22676
rect 152596 21388 152660 21452
rect 125732 21252 125796 21316
rect 152780 21252 152844 21316
rect 144316 19892 144380 19956
rect 167868 18532 167932 18596
rect 141004 17308 141068 17372
rect 149652 17172 149716 17236
rect 152964 15812 153028 15876
rect 130884 14724 130948 14788
rect 154252 14588 154316 14652
rect 154068 14452 154132 14516
rect 143212 13636 143276 13700
rect 145604 13500 145668 13564
rect 154436 13364 154500 13428
rect 160876 13228 160940 13292
rect 165476 13092 165540 13156
rect 169340 12956 169404 13020
rect 147076 12276 147140 12340
rect 149836 12140 149900 12204
rect 151492 12004 151556 12068
rect 162532 11868 162596 11932
rect 162348 11732 162412 11796
rect 170812 11596 170876 11660
rect 136220 10916 136284 10980
rect 148364 10644 148428 10708
rect 151676 10508 151740 10572
rect 134012 10372 134076 10436
rect 158852 10372 158916 10436
rect 133092 10236 133156 10300
rect 159036 10236 159100 10300
rect 131068 9148 131132 9212
rect 147260 9148 147324 9212
rect 129780 9012 129844 9076
rect 162164 9012 162228 9076
rect 128676 8876 128740 8940
rect 170444 8876 170508 8940
rect 142844 7788 142908 7852
rect 133828 7652 133892 7716
rect 158300 7652 158364 7716
rect 127020 7516 127084 7580
rect 168052 7516 168116 7580
rect 147444 6292 147508 6356
rect 150020 6156 150084 6220
rect 158484 4932 158548 4996
rect 137876 4796 137940 4860
rect 163636 4796 163700 4860
rect 136404 3572 136468 3636
rect 131988 3436 132052 3500
rect 134932 3300 134996 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 248684 47414 263898
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 248684 51914 268398
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 248684 56414 272898
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 248684 60914 277398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 248684 65414 281898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 248684 69914 250398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 248684 74414 254898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 248684 78914 259398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 248684 83414 263898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 248684 87914 268398
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 248684 92414 272898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 248684 96914 277398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 248684 101414 281898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 248684 105914 250398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 248684 110414 254898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 248684 114914 259398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 248684 119414 263898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 248684 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 248684 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 248684 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 248684 137414 281898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 248684 141914 250398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 248684 146414 254898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 248684 150914 259398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 248684 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 248684 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 248684 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 248684 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 248684 173414 281898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 248684 177914 250398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 248684 182414 254898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 248684 186914 259398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 248684 191414 263898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 248684 195914 268398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 248684 200414 272898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 248684 204914 277398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 248684 209414 281898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 248684 213914 250398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 248684 218414 254898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 248684 222914 259398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 248684 227414 263898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 248684 231914 268398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 248684 236414 272898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 248684 240914 277398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 248684 245414 281898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 248684 249914 250398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 248684 254414 254898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 248684 258914 259398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 248684 263414 263898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 248684 267914 268398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 248684 272414 272898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 248684 276914 277398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 248684 281414 281898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 248684 285914 250398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 248684 290414 254898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 248684 294914 259398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 248684 299414 263898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 248684 303914 268398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 248684 308414 272898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 248684 312914 277398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 248684 317414 281898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 248684 321914 250398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 248684 326414 254898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 248684 330914 259398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 248684 335414 263898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 248684 339914 268398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 248684 344414 272898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 248684 348914 277398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 248684 353414 281898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 248684 357914 250398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 248684 362414 254898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 248684 366914 259398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 248684 371414 263898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 248684 375914 268398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 248684 380414 272898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 248684 384914 277398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 248684 389414 281898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 396579 696964 396645 696965
rect 396579 696900 396580 696964
rect 396644 696900 396645 696964
rect 396579 696899 396645 696900
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 248684 393914 250398
rect 65300 246303 70100 246486
rect 65300 246067 65342 246303
rect 65578 246067 65662 246303
rect 65898 246067 65982 246303
rect 66218 246067 66302 246303
rect 66538 246067 66622 246303
rect 66858 246067 66942 246303
rect 67178 246067 67262 246303
rect 67498 246067 67582 246303
rect 67818 246067 67902 246303
rect 68138 246067 68222 246303
rect 68458 246067 68542 246303
rect 68778 246067 68862 246303
rect 69098 246067 69182 246303
rect 69418 246067 69502 246303
rect 69738 246067 69822 246303
rect 70058 246067 70100 246303
rect 65300 245884 70100 246067
rect 65300 241953 71300 241984
rect 65300 241717 65462 241953
rect 65698 241717 65782 241953
rect 66018 241717 66102 241953
rect 66338 241717 66422 241953
rect 66658 241717 66742 241953
rect 66978 241717 67062 241953
rect 67298 241717 67382 241953
rect 67618 241717 67702 241953
rect 67938 241717 68022 241953
rect 68258 241717 68342 241953
rect 68578 241717 68662 241953
rect 68898 241717 68982 241953
rect 69218 241717 69302 241953
rect 69538 241717 69622 241953
rect 69858 241717 69942 241953
rect 70178 241717 70262 241953
rect 70498 241717 70582 241953
rect 70818 241717 70902 241953
rect 71138 241717 71300 241953
rect 65300 241633 71300 241717
rect 65300 241397 65462 241633
rect 65698 241397 65782 241633
rect 66018 241397 66102 241633
rect 66338 241397 66422 241633
rect 66658 241397 66742 241633
rect 66978 241397 67062 241633
rect 67298 241397 67382 241633
rect 67618 241397 67702 241633
rect 67938 241397 68022 241633
rect 68258 241397 68342 241633
rect 68578 241397 68662 241633
rect 68898 241397 68982 241633
rect 69218 241397 69302 241633
rect 69538 241397 69622 241633
rect 69858 241397 69942 241633
rect 70178 241397 70262 241633
rect 70498 241397 70582 241633
rect 70818 241397 70902 241633
rect 71138 241397 71300 241633
rect 65300 241366 71300 241397
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 228453 47414 228484
rect 46794 228217 46826 228453
rect 47062 228217 47146 228453
rect 47382 228217 47414 228453
rect 46794 228133 47414 228217
rect 46794 227897 46826 228133
rect 47062 227897 47146 228133
rect 47382 227897 47414 228133
rect 46794 192454 47414 227897
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 196954 51914 228484
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 201454 56414 228484
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 205954 60914 228484
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 210454 65414 228484
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 214954 69914 228484
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 219454 74414 228484
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 223954 78914 228484
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 228453 83414 228484
rect 82794 228217 82826 228453
rect 83062 228217 83146 228453
rect 83382 228217 83414 228453
rect 82794 228133 83414 228217
rect 82794 227897 82826 228133
rect 83062 227897 83146 228133
rect 83382 227897 83414 228133
rect 82794 192454 83414 227897
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 196954 87914 228484
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 201454 92414 228484
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 205954 96914 228484
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 210454 101414 228484
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 214954 105914 228484
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 219454 110414 228484
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 223954 114914 228484
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 118794 228453 119414 228484
rect 118794 228217 118826 228453
rect 119062 228217 119146 228453
rect 119382 228217 119414 228453
rect 118794 228133 119414 228217
rect 118794 227897 118826 228133
rect 119062 227897 119146 228133
rect 119382 227897 119414 228133
rect 118794 192454 119414 227897
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 142000 119414 155898
rect 123294 196954 123914 228484
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 142000 123914 160398
rect 127794 201454 128414 228484
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 142000 128414 164898
rect 132294 205954 132914 228484
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 135914 205954 165514 205986
rect 135914 205718 136036 205954
rect 136272 205718 136356 205954
rect 136592 205718 136676 205954
rect 136912 205718 136996 205954
rect 137232 205718 137316 205954
rect 137552 205718 137636 205954
rect 137872 205718 137956 205954
rect 138192 205718 138276 205954
rect 138512 205718 138596 205954
rect 138832 205718 138916 205954
rect 139152 205718 139236 205954
rect 139472 205718 139556 205954
rect 139792 205718 139876 205954
rect 140112 205718 140196 205954
rect 140432 205718 140516 205954
rect 140752 205718 140836 205954
rect 141072 205718 141156 205954
rect 141392 205718 141476 205954
rect 141712 205718 141796 205954
rect 142032 205718 142116 205954
rect 142352 205718 142436 205954
rect 142672 205718 142756 205954
rect 142992 205718 143076 205954
rect 143312 205718 143396 205954
rect 143632 205718 143716 205954
rect 143952 205718 144036 205954
rect 144272 205718 144356 205954
rect 144592 205718 144676 205954
rect 144912 205718 144996 205954
rect 145232 205718 145316 205954
rect 145552 205718 145636 205954
rect 145872 205718 145956 205954
rect 146192 205718 146276 205954
rect 146512 205718 146596 205954
rect 146832 205718 146916 205954
rect 147152 205718 147236 205954
rect 147472 205718 147556 205954
rect 147792 205718 147876 205954
rect 148112 205718 148196 205954
rect 148432 205718 148516 205954
rect 148752 205718 148836 205954
rect 149072 205718 149156 205954
rect 149392 205718 149476 205954
rect 149712 205718 149796 205954
rect 150032 205718 150116 205954
rect 150352 205718 150436 205954
rect 150672 205718 150756 205954
rect 150992 205718 151076 205954
rect 151312 205718 151396 205954
rect 151632 205718 151716 205954
rect 151952 205718 152036 205954
rect 152272 205718 152356 205954
rect 152592 205718 152676 205954
rect 152912 205718 152996 205954
rect 153232 205718 153316 205954
rect 153552 205718 153636 205954
rect 153872 205718 153956 205954
rect 154192 205718 154276 205954
rect 154512 205718 154596 205954
rect 154832 205718 154916 205954
rect 155152 205718 155236 205954
rect 155472 205718 155556 205954
rect 155792 205718 155876 205954
rect 156112 205718 156196 205954
rect 156432 205718 156516 205954
rect 156752 205718 156836 205954
rect 157072 205718 157156 205954
rect 157392 205718 157476 205954
rect 157712 205718 157796 205954
rect 158032 205718 158116 205954
rect 158352 205718 158436 205954
rect 158672 205718 158756 205954
rect 158992 205718 159076 205954
rect 159312 205718 159396 205954
rect 159632 205718 159716 205954
rect 159952 205718 160036 205954
rect 160272 205718 160356 205954
rect 160592 205718 160676 205954
rect 160912 205718 160996 205954
rect 161232 205718 161316 205954
rect 161552 205718 161636 205954
rect 161872 205718 161956 205954
rect 162192 205718 162276 205954
rect 162512 205718 162596 205954
rect 162832 205718 162916 205954
rect 163152 205718 163236 205954
rect 163472 205718 163556 205954
rect 163792 205718 163876 205954
rect 164112 205718 164196 205954
rect 164432 205718 164516 205954
rect 164752 205718 164836 205954
rect 165072 205718 165156 205954
rect 165392 205718 165514 205954
rect 135914 205634 165514 205718
rect 135914 205398 136036 205634
rect 136272 205398 136356 205634
rect 136592 205398 136676 205634
rect 136912 205398 136996 205634
rect 137232 205398 137316 205634
rect 137552 205398 137636 205634
rect 137872 205398 137956 205634
rect 138192 205398 138276 205634
rect 138512 205398 138596 205634
rect 138832 205398 138916 205634
rect 139152 205398 139236 205634
rect 139472 205398 139556 205634
rect 139792 205398 139876 205634
rect 140112 205398 140196 205634
rect 140432 205398 140516 205634
rect 140752 205398 140836 205634
rect 141072 205398 141156 205634
rect 141392 205398 141476 205634
rect 141712 205398 141796 205634
rect 142032 205398 142116 205634
rect 142352 205398 142436 205634
rect 142672 205398 142756 205634
rect 142992 205398 143076 205634
rect 143312 205398 143396 205634
rect 143632 205398 143716 205634
rect 143952 205398 144036 205634
rect 144272 205398 144356 205634
rect 144592 205398 144676 205634
rect 144912 205398 144996 205634
rect 145232 205398 145316 205634
rect 145552 205398 145636 205634
rect 145872 205398 145956 205634
rect 146192 205398 146276 205634
rect 146512 205398 146596 205634
rect 146832 205398 146916 205634
rect 147152 205398 147236 205634
rect 147472 205398 147556 205634
rect 147792 205398 147876 205634
rect 148112 205398 148196 205634
rect 148432 205398 148516 205634
rect 148752 205398 148836 205634
rect 149072 205398 149156 205634
rect 149392 205398 149476 205634
rect 149712 205398 149796 205634
rect 150032 205398 150116 205634
rect 150352 205398 150436 205634
rect 150672 205398 150756 205634
rect 150992 205398 151076 205634
rect 151312 205398 151396 205634
rect 151632 205398 151716 205634
rect 151952 205398 152036 205634
rect 152272 205398 152356 205634
rect 152592 205398 152676 205634
rect 152912 205398 152996 205634
rect 153232 205398 153316 205634
rect 153552 205398 153636 205634
rect 153872 205398 153956 205634
rect 154192 205398 154276 205634
rect 154512 205398 154596 205634
rect 154832 205398 154916 205634
rect 155152 205398 155236 205634
rect 155472 205398 155556 205634
rect 155792 205398 155876 205634
rect 156112 205398 156196 205634
rect 156432 205398 156516 205634
rect 156752 205398 156836 205634
rect 157072 205398 157156 205634
rect 157392 205398 157476 205634
rect 157712 205398 157796 205634
rect 158032 205398 158116 205634
rect 158352 205398 158436 205634
rect 158672 205398 158756 205634
rect 158992 205398 159076 205634
rect 159312 205398 159396 205634
rect 159632 205398 159716 205634
rect 159952 205398 160036 205634
rect 160272 205398 160356 205634
rect 160592 205398 160676 205634
rect 160912 205398 160996 205634
rect 161232 205398 161316 205634
rect 161552 205398 161636 205634
rect 161872 205398 161956 205634
rect 162192 205398 162276 205634
rect 162512 205398 162596 205634
rect 162832 205398 162916 205634
rect 163152 205398 163236 205634
rect 163472 205398 163556 205634
rect 163792 205398 163876 205634
rect 164112 205398 164196 205634
rect 164432 205398 164516 205634
rect 164752 205398 164836 205634
rect 165072 205398 165156 205634
rect 165392 205398 165514 205634
rect 135914 205366 165514 205398
rect 168294 205954 168914 228484
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 137314 201454 165514 201486
rect 137314 201218 137376 201454
rect 137612 201218 137696 201454
rect 137932 201218 138016 201454
rect 138252 201218 138336 201454
rect 138572 201218 138656 201454
rect 138892 201218 138976 201454
rect 139212 201218 139296 201454
rect 139532 201218 139616 201454
rect 139852 201218 139936 201454
rect 140172 201218 140256 201454
rect 140492 201218 140576 201454
rect 140812 201218 140896 201454
rect 141132 201218 141216 201454
rect 141452 201218 141536 201454
rect 141772 201218 141856 201454
rect 142092 201218 142176 201454
rect 142412 201218 142496 201454
rect 142732 201218 142816 201454
rect 143052 201218 143136 201454
rect 143372 201218 143456 201454
rect 143692 201218 143776 201454
rect 144012 201218 144096 201454
rect 144332 201218 144416 201454
rect 144652 201218 144736 201454
rect 144972 201218 145056 201454
rect 145292 201218 145376 201454
rect 145612 201218 145696 201454
rect 145932 201218 146016 201454
rect 146252 201218 146336 201454
rect 146572 201218 146656 201454
rect 146892 201218 146976 201454
rect 147212 201218 147296 201454
rect 147532 201218 147616 201454
rect 147852 201218 147936 201454
rect 148172 201218 148256 201454
rect 148492 201218 148576 201454
rect 148812 201218 148896 201454
rect 149132 201218 149216 201454
rect 149452 201218 149536 201454
rect 149772 201218 149856 201454
rect 150092 201218 150176 201454
rect 150412 201218 150496 201454
rect 150732 201218 150816 201454
rect 151052 201218 151136 201454
rect 151372 201218 151456 201454
rect 151692 201218 151776 201454
rect 152012 201218 152096 201454
rect 152332 201218 152416 201454
rect 152652 201218 152736 201454
rect 152972 201218 153056 201454
rect 153292 201218 153376 201454
rect 153612 201218 153696 201454
rect 153932 201218 154016 201454
rect 154252 201218 154336 201454
rect 154572 201218 154656 201454
rect 154892 201218 154976 201454
rect 155212 201218 155296 201454
rect 155532 201218 155616 201454
rect 155852 201218 155936 201454
rect 156172 201218 156256 201454
rect 156492 201218 156576 201454
rect 156812 201218 156896 201454
rect 157132 201218 157216 201454
rect 157452 201218 157536 201454
rect 157772 201218 157856 201454
rect 158092 201218 158176 201454
rect 158412 201218 158496 201454
rect 158732 201218 158816 201454
rect 159052 201218 159136 201454
rect 159372 201218 159456 201454
rect 159692 201218 159776 201454
rect 160012 201218 160096 201454
rect 160332 201218 160416 201454
rect 160652 201218 160736 201454
rect 160972 201218 161056 201454
rect 161292 201218 161376 201454
rect 161612 201218 161696 201454
rect 161932 201218 162016 201454
rect 162252 201218 162336 201454
rect 162572 201218 162656 201454
rect 162892 201218 162976 201454
rect 163212 201218 163296 201454
rect 163532 201218 163616 201454
rect 163852 201218 163936 201454
rect 164172 201218 164256 201454
rect 164492 201218 164576 201454
rect 164812 201218 164896 201454
rect 165132 201218 165216 201454
rect 165452 201218 165514 201454
rect 137314 201134 165514 201218
rect 137314 200898 137376 201134
rect 137612 200898 137696 201134
rect 137932 200898 138016 201134
rect 138252 200898 138336 201134
rect 138572 200898 138656 201134
rect 138892 200898 138976 201134
rect 139212 200898 139296 201134
rect 139532 200898 139616 201134
rect 139852 200898 139936 201134
rect 140172 200898 140256 201134
rect 140492 200898 140576 201134
rect 140812 200898 140896 201134
rect 141132 200898 141216 201134
rect 141452 200898 141536 201134
rect 141772 200898 141856 201134
rect 142092 200898 142176 201134
rect 142412 200898 142496 201134
rect 142732 200898 142816 201134
rect 143052 200898 143136 201134
rect 143372 200898 143456 201134
rect 143692 200898 143776 201134
rect 144012 200898 144096 201134
rect 144332 200898 144416 201134
rect 144652 200898 144736 201134
rect 144972 200898 145056 201134
rect 145292 200898 145376 201134
rect 145612 200898 145696 201134
rect 145932 200898 146016 201134
rect 146252 200898 146336 201134
rect 146572 200898 146656 201134
rect 146892 200898 146976 201134
rect 147212 200898 147296 201134
rect 147532 200898 147616 201134
rect 147852 200898 147936 201134
rect 148172 200898 148256 201134
rect 148492 200898 148576 201134
rect 148812 200898 148896 201134
rect 149132 200898 149216 201134
rect 149452 200898 149536 201134
rect 149772 200898 149856 201134
rect 150092 200898 150176 201134
rect 150412 200898 150496 201134
rect 150732 200898 150816 201134
rect 151052 200898 151136 201134
rect 151372 200898 151456 201134
rect 151692 200898 151776 201134
rect 152012 200898 152096 201134
rect 152332 200898 152416 201134
rect 152652 200898 152736 201134
rect 152972 200898 153056 201134
rect 153292 200898 153376 201134
rect 153612 200898 153696 201134
rect 153932 200898 154016 201134
rect 154252 200898 154336 201134
rect 154572 200898 154656 201134
rect 154892 200898 154976 201134
rect 155212 200898 155296 201134
rect 155532 200898 155616 201134
rect 155852 200898 155936 201134
rect 156172 200898 156256 201134
rect 156492 200898 156576 201134
rect 156812 200898 156896 201134
rect 157132 200898 157216 201134
rect 157452 200898 157536 201134
rect 157772 200898 157856 201134
rect 158092 200898 158176 201134
rect 158412 200898 158496 201134
rect 158732 200898 158816 201134
rect 159052 200898 159136 201134
rect 159372 200898 159456 201134
rect 159692 200898 159776 201134
rect 160012 200898 160096 201134
rect 160332 200898 160416 201134
rect 160652 200898 160736 201134
rect 160972 200898 161056 201134
rect 161292 200898 161376 201134
rect 161612 200898 161696 201134
rect 161932 200898 162016 201134
rect 162252 200898 162336 201134
rect 162572 200898 162656 201134
rect 162892 200898 162976 201134
rect 163212 200898 163296 201134
rect 163532 200898 163616 201134
rect 163852 200898 163936 201134
rect 164172 200898 164256 201134
rect 164492 200898 164576 201134
rect 164812 200898 164896 201134
rect 165132 200898 165216 201134
rect 165452 200898 165514 201134
rect 137314 200866 165514 200898
rect 144683 200700 144749 200701
rect 144683 200636 144684 200700
rect 144748 200636 144749 200700
rect 144683 200635 144749 200636
rect 144686 195669 144746 200635
rect 147627 199340 147693 199341
rect 147627 199276 147628 199340
rect 147692 199276 147693 199340
rect 147627 199275 147693 199276
rect 147630 196485 147690 199275
rect 147627 196484 147693 196485
rect 147627 196420 147628 196484
rect 147692 196420 147693 196484
rect 147627 196419 147693 196420
rect 151307 196076 151373 196077
rect 151307 196012 151308 196076
rect 151372 196012 151373 196076
rect 151307 196011 151373 196012
rect 144683 195668 144749 195669
rect 144683 195604 144684 195668
rect 144748 195604 144749 195668
rect 144683 195603 144749 195604
rect 149835 195668 149901 195669
rect 149835 195604 149836 195668
rect 149900 195604 149901 195668
rect 149835 195603 149901 195604
rect 143579 191808 143645 191809
rect 143579 191744 143580 191808
rect 143644 191744 143645 191808
rect 143579 191743 143645 191744
rect 141739 191316 141805 191317
rect 141739 191252 141740 191316
rect 141804 191252 141805 191316
rect 141739 191251 141805 191252
rect 140635 186964 140701 186965
rect 140635 186900 140636 186964
rect 140700 186900 140701 186964
rect 140635 186899 140701 186900
rect 140451 179212 140517 179213
rect 140451 179148 140452 179212
rect 140516 179148 140517 179212
rect 140451 179147 140517 179148
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 142000 132914 169398
rect 140454 143173 140514 179147
rect 140451 143172 140517 143173
rect 140451 143108 140452 143172
rect 140516 143108 140517 143172
rect 140451 143107 140517 143108
rect 140638 142765 140698 186899
rect 141742 166429 141802 191251
rect 141923 190636 141989 190637
rect 141923 190572 141924 190636
rect 141988 190572 141989 190636
rect 141923 190571 141989 190572
rect 141739 166428 141805 166429
rect 141739 166364 141740 166428
rect 141804 166364 141805 166428
rect 141739 166363 141805 166364
rect 141926 166293 141986 190571
rect 142659 178804 142725 178805
rect 142659 178740 142660 178804
rect 142724 178740 142725 178804
rect 142659 178739 142725 178740
rect 142662 176765 142722 178739
rect 142659 176764 142725 176765
rect 142659 176700 142660 176764
rect 142724 176700 142725 176764
rect 142659 176699 142725 176700
rect 142475 173908 142541 173909
rect 142475 173844 142476 173908
rect 142540 173844 142541 173908
rect 142475 173843 142541 173844
rect 142291 173772 142357 173773
rect 142291 173708 142292 173772
rect 142356 173708 142357 173772
rect 142291 173707 142357 173708
rect 142107 171324 142173 171325
rect 142107 171260 142108 171324
rect 142172 171260 142173 171324
rect 142107 171259 142173 171260
rect 142110 170917 142170 171259
rect 142107 170916 142173 170917
rect 142107 170852 142108 170916
rect 142172 170852 142173 170916
rect 142107 170851 142173 170852
rect 141923 166292 141989 166293
rect 141923 166228 141924 166292
rect 141988 166228 141989 166292
rect 141923 166227 141989 166228
rect 142107 161532 142173 161533
rect 142107 161530 142108 161532
rect 141926 161470 142108 161530
rect 140635 142764 140701 142765
rect 140635 142700 140636 142764
rect 140700 142700 140701 142764
rect 140635 142699 140701 142700
rect 141926 142490 141986 161470
rect 142107 161468 142108 161470
rect 142172 161468 142173 161532
rect 142107 161467 142173 161468
rect 142107 142492 142173 142493
rect 142107 142490 142108 142492
rect 141926 142430 142108 142490
rect 142107 142428 142108 142430
rect 142172 142428 142173 142492
rect 142107 142427 142173 142428
rect 142294 142221 142354 173707
rect 142478 143445 142538 173843
rect 142659 173636 142725 173637
rect 142659 173572 142660 173636
rect 142724 173572 142725 173636
rect 142659 173571 142725 173572
rect 142475 143444 142541 143445
rect 142475 143380 142476 143444
rect 142540 143380 142541 143444
rect 142475 143379 142541 143380
rect 142662 143309 142722 173571
rect 142659 143308 142725 143309
rect 142659 143244 142660 143308
rect 142724 143244 142725 143308
rect 142659 143243 142725 143244
rect 143582 142629 143642 191743
rect 149838 190637 149898 195603
rect 151310 191319 151370 196011
rect 151307 191318 151373 191319
rect 151307 191254 151308 191318
rect 151372 191254 151373 191318
rect 151307 191253 151373 191254
rect 149835 190636 149901 190637
rect 149835 190572 149836 190636
rect 149900 190572 149901 190636
rect 149835 190571 149901 190572
rect 146155 180708 146221 180709
rect 146155 180644 146156 180708
rect 146220 180644 146221 180708
rect 146155 180643 146221 180644
rect 144131 173772 144197 173773
rect 144131 173708 144132 173772
rect 144196 173708 144197 173772
rect 144131 173707 144197 173708
rect 144134 143037 144194 173707
rect 144131 143036 144197 143037
rect 144131 142972 144132 143036
rect 144196 142972 144197 143036
rect 144131 142971 144197 142972
rect 146158 142901 146218 180643
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 146155 142900 146221 142901
rect 146155 142836 146156 142900
rect 146220 142836 146221 142900
rect 146155 142835 146221 142836
rect 143579 142628 143645 142629
rect 143579 142564 143580 142628
rect 143644 142564 143645 142628
rect 143579 142563 143645 142564
rect 142291 142220 142357 142221
rect 142291 142156 142292 142220
rect 142356 142156 142357 142220
rect 142291 142155 142357 142156
rect 168294 142000 168914 169398
rect 172794 210454 173414 228484
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 142000 173414 173898
rect 177294 214954 177914 228484
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 142000 177914 142398
rect 181794 219454 182414 228484
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 142000 182414 146898
rect 186294 223954 186914 228484
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 139568 115954 139888 115986
rect 139568 115718 139610 115954
rect 139846 115718 139888 115954
rect 139568 115634 139888 115718
rect 139568 115398 139610 115634
rect 139846 115398 139888 115634
rect 139568 115366 139888 115398
rect 170288 115954 170608 115986
rect 170288 115718 170330 115954
rect 170566 115718 170608 115954
rect 170288 115634 170608 115718
rect 170288 115398 170330 115634
rect 170566 115398 170608 115634
rect 170288 115366 170608 115398
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 168051 80612 168117 80613
rect 168051 80548 168052 80612
rect 168116 80548 168117 80612
rect 168051 80547 168117 80548
rect 161979 80204 162045 80205
rect 161979 80140 161980 80204
rect 162044 80140 162045 80204
rect 161979 80139 162045 80140
rect 160139 80068 160205 80069
rect 160139 80004 160140 80068
rect 160204 80004 160205 80068
rect 160139 80003 160205 80004
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 125547 79932 125613 79933
rect 125547 79868 125548 79932
rect 125612 79868 125613 79932
rect 125547 79867 125613 79868
rect 128675 79932 128741 79933
rect 128675 79868 128676 79932
rect 128740 79930 128741 79932
rect 129043 79932 129109 79933
rect 128740 79870 128922 79930
rect 128740 79868 128741 79870
rect 128675 79867 128741 79868
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 78000
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 78000
rect 125550 64890 125610 79867
rect 127019 79796 127085 79797
rect 127019 79732 127020 79796
rect 127084 79732 127085 79796
rect 127019 79731 127085 79732
rect 128675 79796 128741 79797
rect 128675 79732 128676 79796
rect 128740 79732 128741 79796
rect 128675 79731 128741 79732
rect 125550 64830 125794 64890
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 125734 21317 125794 64830
rect 125731 21316 125797 21317
rect 125731 21252 125732 21316
rect 125796 21252 125797 21316
rect 125731 21251 125797 21252
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 127022 7581 127082 79731
rect 128491 78164 128557 78165
rect 128491 78100 128492 78164
rect 128556 78100 128557 78164
rect 128491 78099 128557 78100
rect 127203 75988 127269 75989
rect 127203 75924 127204 75988
rect 127268 75924 127269 75988
rect 127203 75923 127269 75924
rect 127206 35189 127266 75923
rect 127794 57454 128414 78000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127203 35188 127269 35189
rect 127203 35124 127204 35188
rect 127268 35124 127269 35188
rect 127203 35123 127269 35124
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127019 7580 127085 7581
rect 127019 7516 127020 7580
rect 127084 7516 127085 7580
rect 127019 7515 127085 7516
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 -4186 128414 20898
rect 128494 16590 128554 78099
rect 128678 71790 128738 79731
rect 128862 76394 128922 79870
rect 129043 79868 129044 79932
rect 129108 79868 129109 79932
rect 129043 79867 129109 79868
rect 129779 79932 129845 79933
rect 129779 79868 129780 79932
rect 129844 79868 129845 79932
rect 129779 79867 129845 79868
rect 130883 79932 130949 79933
rect 130883 79868 130884 79932
rect 130948 79868 130949 79932
rect 130883 79867 130949 79868
rect 133091 79932 133157 79933
rect 133091 79868 133092 79932
rect 133156 79868 133157 79932
rect 133091 79867 133157 79868
rect 133275 79932 133341 79933
rect 133275 79868 133276 79932
rect 133340 79868 133341 79932
rect 133275 79867 133341 79868
rect 133827 79932 133893 79933
rect 133827 79868 133828 79932
rect 133892 79868 133893 79932
rect 135483 79932 135549 79933
rect 135483 79930 135484 79932
rect 133827 79867 133893 79868
rect 135302 79870 135484 79930
rect 129046 77621 129106 79867
rect 129043 77620 129109 77621
rect 129043 77556 129044 77620
rect 129108 77556 129109 77620
rect 129043 77555 129109 77556
rect 128862 76334 129106 76394
rect 128678 71730 128922 71790
rect 128862 71093 128922 71730
rect 129046 71229 129106 76334
rect 129043 71228 129109 71229
rect 129043 71164 129044 71228
rect 129108 71164 129109 71228
rect 129043 71163 129109 71164
rect 128859 71092 128925 71093
rect 128859 71028 128860 71092
rect 128924 71028 128925 71092
rect 128859 71027 128925 71028
rect 128494 16530 128738 16590
rect 128678 8941 128738 16530
rect 129782 9077 129842 79867
rect 130886 78301 130946 79867
rect 131251 79796 131317 79797
rect 131251 79732 131252 79796
rect 131316 79732 131317 79796
rect 131251 79731 131317 79732
rect 130883 78300 130949 78301
rect 130883 78236 130884 78300
rect 130948 78236 130949 78300
rect 130883 78235 130949 78236
rect 130883 77620 130949 77621
rect 130883 77556 130884 77620
rect 130948 77556 130949 77620
rect 130883 77555 130949 77556
rect 129963 77348 130029 77349
rect 129963 77284 129964 77348
rect 130028 77284 130029 77348
rect 129963 77283 130029 77284
rect 129966 68237 130026 77283
rect 129963 68236 130029 68237
rect 129963 68172 129964 68236
rect 130028 68172 130029 68236
rect 129963 68171 130029 68172
rect 130886 14789 130946 77555
rect 131067 77212 131133 77213
rect 131067 77148 131068 77212
rect 131132 77148 131133 77212
rect 131067 77147 131133 77148
rect 130883 14788 130949 14789
rect 130883 14724 130884 14788
rect 130948 14724 130949 14788
rect 130883 14723 130949 14724
rect 131070 9213 131130 77147
rect 131254 69597 131314 79731
rect 133094 78301 133154 79867
rect 133278 78709 133338 79867
rect 133643 79660 133709 79661
rect 133643 79596 133644 79660
rect 133708 79596 133709 79660
rect 133643 79595 133709 79596
rect 133275 78708 133341 78709
rect 133275 78644 133276 78708
rect 133340 78644 133341 78708
rect 133275 78643 133341 78644
rect 133275 78436 133341 78437
rect 133275 78372 133276 78436
rect 133340 78372 133341 78436
rect 133275 78371 133341 78372
rect 133091 78300 133157 78301
rect 133091 78236 133092 78300
rect 133156 78236 133157 78300
rect 133091 78235 133157 78236
rect 133091 78164 133157 78165
rect 133091 78100 133092 78164
rect 133156 78100 133157 78164
rect 133091 78099 133157 78100
rect 131987 77892 132053 77893
rect 131987 77828 131988 77892
rect 132052 77828 132053 77892
rect 131987 77827 132053 77828
rect 131435 77348 131501 77349
rect 131435 77284 131436 77348
rect 131500 77284 131501 77348
rect 131435 77283 131501 77284
rect 131438 72453 131498 77283
rect 131435 72452 131501 72453
rect 131435 72388 131436 72452
rect 131500 72388 131501 72452
rect 131435 72387 131501 72388
rect 131251 69596 131317 69597
rect 131251 69532 131252 69596
rect 131316 69532 131317 69596
rect 131251 69531 131317 69532
rect 131067 9212 131133 9213
rect 131067 9148 131068 9212
rect 131132 9148 131133 9212
rect 131067 9147 131133 9148
rect 129779 9076 129845 9077
rect 129779 9012 129780 9076
rect 129844 9012 129845 9076
rect 129779 9011 129845 9012
rect 128675 8940 128741 8941
rect 128675 8876 128676 8940
rect 128740 8876 128741 8940
rect 128675 8875 128741 8876
rect 131990 3501 132050 77827
rect 132294 61954 132914 78000
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 131987 3500 132053 3501
rect 131987 3436 131988 3500
rect 132052 3436 132053 3500
rect 131987 3435 132053 3436
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 -5146 132914 25398
rect 133094 10301 133154 78099
rect 133278 68373 133338 78371
rect 133646 77213 133706 79595
rect 133643 77212 133709 77213
rect 133643 77148 133644 77212
rect 133708 77148 133709 77212
rect 133643 77147 133709 77148
rect 133275 68372 133341 68373
rect 133275 68308 133276 68372
rect 133340 68308 133341 68372
rect 133275 68307 133341 68308
rect 133091 10300 133157 10301
rect 133091 10236 133092 10300
rect 133156 10236 133157 10300
rect 133091 10235 133157 10236
rect 133830 7717 133890 79867
rect 134011 78708 134077 78709
rect 134011 78644 134012 78708
rect 134076 78644 134077 78708
rect 134011 78643 134077 78644
rect 134014 10437 134074 78643
rect 134931 78300 134997 78301
rect 134931 78236 134932 78300
rect 134996 78236 134997 78300
rect 134931 78235 134997 78236
rect 134011 10436 134077 10437
rect 134011 10372 134012 10436
rect 134076 10372 134077 10436
rect 134011 10371 134077 10372
rect 133827 7716 133893 7717
rect 133827 7652 133828 7716
rect 133892 7652 133893 7716
rect 133827 7651 133893 7652
rect 134934 3365 134994 78235
rect 135302 69597 135362 79870
rect 135483 79868 135484 79870
rect 135548 79868 135549 79932
rect 135483 79867 135549 79868
rect 136219 79932 136285 79933
rect 136219 79868 136220 79932
rect 136284 79868 136285 79932
rect 136219 79867 136285 79868
rect 137691 79932 137757 79933
rect 137691 79868 137692 79932
rect 137756 79868 137757 79932
rect 137691 79867 137757 79868
rect 138979 79932 139045 79933
rect 138979 79868 138980 79932
rect 139044 79868 139045 79932
rect 138979 79867 139045 79868
rect 139347 79932 139413 79933
rect 139347 79868 139348 79932
rect 139412 79868 139413 79932
rect 139347 79867 139413 79868
rect 142291 79932 142357 79933
rect 142291 79868 142292 79932
rect 142356 79868 142357 79932
rect 142291 79867 142357 79868
rect 144315 79932 144381 79933
rect 144315 79868 144316 79932
rect 144380 79868 144381 79932
rect 144315 79867 144381 79868
rect 145051 79932 145117 79933
rect 145051 79868 145052 79932
rect 145116 79868 145117 79932
rect 145051 79867 145117 79868
rect 145787 79932 145853 79933
rect 145787 79868 145788 79932
rect 145852 79868 145853 79932
rect 145787 79867 145853 79868
rect 146155 79932 146221 79933
rect 146155 79868 146156 79932
rect 146220 79868 146221 79932
rect 146155 79867 146221 79868
rect 147259 79932 147325 79933
rect 147259 79868 147260 79932
rect 147324 79868 147325 79932
rect 147259 79867 147325 79868
rect 149835 79932 149901 79933
rect 149835 79868 149836 79932
rect 149900 79868 149901 79932
rect 149835 79867 149901 79868
rect 150939 79932 151005 79933
rect 150939 79868 150940 79932
rect 151004 79868 151005 79932
rect 150939 79867 151005 79868
rect 152779 79932 152845 79933
rect 152779 79868 152780 79932
rect 152844 79868 152845 79932
rect 152779 79867 152845 79868
rect 153699 79932 153765 79933
rect 153699 79868 153700 79932
rect 153764 79868 153765 79932
rect 153699 79867 153765 79868
rect 154435 79932 154501 79933
rect 154435 79868 154436 79932
rect 154500 79868 154501 79932
rect 154435 79867 154501 79868
rect 154619 79932 154685 79933
rect 154619 79868 154620 79932
rect 154684 79868 154685 79932
rect 154619 79867 154685 79868
rect 155355 79932 155421 79933
rect 155355 79868 155356 79932
rect 155420 79868 155421 79932
rect 155355 79867 155421 79868
rect 157379 79932 157445 79933
rect 157379 79868 157380 79932
rect 157444 79868 157445 79932
rect 157379 79867 157445 79868
rect 158115 79932 158181 79933
rect 158115 79868 158116 79932
rect 158180 79868 158181 79932
rect 158115 79867 158181 79868
rect 158667 79932 158733 79933
rect 158667 79868 158668 79932
rect 158732 79868 158733 79932
rect 158667 79867 158733 79868
rect 159955 79932 160021 79933
rect 159955 79868 159956 79932
rect 160020 79868 160021 79932
rect 159955 79867 160021 79868
rect 135483 77348 135549 77349
rect 135483 77284 135484 77348
rect 135548 77284 135549 77348
rect 135483 77283 135549 77284
rect 135486 74493 135546 77283
rect 135483 74492 135549 74493
rect 135483 74428 135484 74492
rect 135548 74428 135549 74492
rect 135483 74427 135549 74428
rect 135299 69596 135365 69597
rect 135299 69532 135300 69596
rect 135364 69532 135365 69596
rect 135299 69531 135365 69532
rect 136222 10981 136282 79867
rect 136955 79796 137021 79797
rect 136955 79732 136956 79796
rect 137020 79732 137021 79796
rect 136955 79731 137021 79732
rect 136958 78709 137018 79731
rect 136955 78708 137021 78709
rect 136955 78644 136956 78708
rect 137020 78644 137021 78708
rect 136955 78643 137021 78644
rect 136403 78164 136469 78165
rect 136403 78100 136404 78164
rect 136468 78100 136469 78164
rect 136403 78099 136469 78100
rect 136219 10980 136285 10981
rect 136219 10916 136220 10980
rect 136284 10916 136285 10980
rect 136219 10915 136285 10916
rect 136406 3637 136466 78099
rect 136794 66454 137414 78000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 137694 44845 137754 79867
rect 137875 79796 137941 79797
rect 137875 79732 137876 79796
rect 137940 79732 137941 79796
rect 137875 79731 137941 79732
rect 138059 79796 138125 79797
rect 138059 79732 138060 79796
rect 138124 79732 138125 79796
rect 138059 79731 138125 79732
rect 138795 79796 138861 79797
rect 138795 79732 138796 79796
rect 138860 79732 138861 79796
rect 138795 79731 138861 79732
rect 137691 44844 137757 44845
rect 137691 44780 137692 44844
rect 137756 44780 137757 44844
rect 137691 44779 137757 44780
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136403 3636 136469 3637
rect 136403 3572 136404 3636
rect 136468 3572 136469 3636
rect 136403 3571 136469 3572
rect 134931 3364 134997 3365
rect 134931 3300 134932 3364
rect 134996 3300 134997 3364
rect 134931 3299 134997 3300
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 -6106 137414 29898
rect 137878 4861 137938 79731
rect 138062 78709 138122 79731
rect 138059 78708 138125 78709
rect 138059 78644 138060 78708
rect 138124 78644 138125 78708
rect 138059 78643 138125 78644
rect 138798 71093 138858 79731
rect 138795 71092 138861 71093
rect 138795 71028 138796 71092
rect 138860 71028 138861 71092
rect 138795 71027 138861 71028
rect 138982 67557 139042 79867
rect 139163 78300 139229 78301
rect 139163 78236 139164 78300
rect 139228 78236 139229 78300
rect 139163 78235 139229 78236
rect 138979 67556 139045 67557
rect 138979 67492 138980 67556
rect 139044 67492 139045 67556
rect 138979 67491 139045 67492
rect 139166 50285 139226 78235
rect 139350 75581 139410 79867
rect 141923 79796 141989 79797
rect 141923 79732 141924 79796
rect 141988 79732 141989 79796
rect 141923 79731 141989 79732
rect 140083 79660 140149 79661
rect 140083 79596 140084 79660
rect 140148 79596 140149 79660
rect 140083 79595 140149 79596
rect 139347 75580 139413 75581
rect 139347 75516 139348 75580
rect 139412 75516 139413 75580
rect 139347 75515 139413 75516
rect 140086 74357 140146 79595
rect 140451 78708 140517 78709
rect 140451 78644 140452 78708
rect 140516 78644 140517 78708
rect 140451 78643 140517 78644
rect 140267 77756 140333 77757
rect 140267 77692 140268 77756
rect 140332 77692 140333 77756
rect 140267 77691 140333 77692
rect 140083 74356 140149 74357
rect 140083 74292 140084 74356
rect 140148 74292 140149 74356
rect 140083 74291 140149 74292
rect 140270 65517 140330 77691
rect 140267 65516 140333 65517
rect 140267 65452 140268 65516
rect 140332 65452 140333 65516
rect 140267 65451 140333 65452
rect 139163 50284 139229 50285
rect 139163 50220 139164 50284
rect 139228 50220 139229 50284
rect 139163 50219 139229 50220
rect 140454 40901 140514 78643
rect 141926 78301 141986 79731
rect 141003 78300 141069 78301
rect 141003 78236 141004 78300
rect 141068 78236 141069 78300
rect 141003 78235 141069 78236
rect 141923 78300 141989 78301
rect 141923 78236 141924 78300
rect 141988 78236 141989 78300
rect 141923 78235 141989 78236
rect 140635 77484 140701 77485
rect 140635 77420 140636 77484
rect 140700 77420 140701 77484
rect 140635 77419 140701 77420
rect 140451 40900 140517 40901
rect 140451 40836 140452 40900
rect 140516 40836 140517 40900
rect 140451 40835 140517 40836
rect 140638 24445 140698 77419
rect 140635 24444 140701 24445
rect 140635 24380 140636 24444
rect 140700 24380 140701 24444
rect 140635 24379 140701 24380
rect 141006 17373 141066 78235
rect 141294 70954 141914 78000
rect 142294 77077 142354 79867
rect 143211 79796 143277 79797
rect 143211 79732 143212 79796
rect 143276 79732 143277 79796
rect 143211 79731 143277 79732
rect 143027 78300 143093 78301
rect 143027 78236 143028 78300
rect 143092 78236 143093 78300
rect 143027 78235 143093 78236
rect 142291 77076 142357 77077
rect 142291 77012 142292 77076
rect 142356 77012 142357 77076
rect 142291 77011 142357 77012
rect 142843 76804 142909 76805
rect 142843 76740 142844 76804
rect 142908 76740 142909 76804
rect 142843 76739 142909 76740
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141003 17372 141069 17373
rect 141003 17308 141004 17372
rect 141068 17308 141069 17372
rect 141003 17307 141069 17308
rect 137875 4860 137941 4861
rect 137875 4796 137876 4860
rect 137940 4796 137941 4860
rect 137875 4795 137941 4796
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 -7066 141914 34398
rect 142846 7853 142906 76739
rect 143030 58581 143090 78235
rect 143027 58580 143093 58581
rect 143027 58516 143028 58580
rect 143092 58516 143093 58580
rect 143027 58515 143093 58516
rect 143214 13701 143274 79731
rect 144318 78709 144378 79867
rect 144499 79796 144565 79797
rect 144499 79732 144500 79796
rect 144564 79732 144565 79796
rect 144499 79731 144565 79732
rect 143395 78708 143461 78709
rect 143395 78644 143396 78708
rect 143460 78644 143461 78708
rect 143395 78643 143461 78644
rect 144315 78708 144381 78709
rect 144315 78644 144316 78708
rect 144380 78644 144381 78708
rect 144315 78643 144381 78644
rect 143398 74221 143458 78643
rect 143395 74220 143461 74221
rect 143395 74156 143396 74220
rect 143460 74156 143461 74220
rect 143395 74155 143461 74156
rect 144315 73676 144381 73677
rect 144315 73612 144316 73676
rect 144380 73612 144381 73676
rect 144315 73611 144381 73612
rect 144318 19957 144378 73611
rect 144502 40765 144562 79731
rect 145054 76397 145114 79867
rect 145603 79660 145669 79661
rect 145603 79658 145604 79660
rect 145238 79598 145604 79658
rect 145051 76396 145117 76397
rect 145051 76332 145052 76396
rect 145116 76332 145117 76396
rect 145051 76331 145117 76332
rect 145238 57493 145298 79598
rect 145603 79596 145604 79598
rect 145668 79596 145669 79660
rect 145603 79595 145669 79596
rect 145790 78709 145850 79867
rect 146158 78709 146218 79867
rect 146523 79660 146589 79661
rect 146523 79596 146524 79660
rect 146588 79596 146589 79660
rect 146523 79595 146589 79596
rect 145787 78708 145853 78709
rect 145787 78644 145788 78708
rect 145852 78644 145853 78708
rect 145787 78643 145853 78644
rect 146155 78708 146221 78709
rect 146155 78644 146156 78708
rect 146220 78644 146221 78708
rect 146155 78643 146221 78644
rect 145603 78164 145669 78165
rect 145603 78100 145604 78164
rect 145668 78100 145669 78164
rect 145603 78099 145669 78100
rect 145419 76532 145485 76533
rect 145419 76468 145420 76532
rect 145484 76468 145485 76532
rect 145419 76467 145485 76468
rect 145235 57492 145301 57493
rect 145235 57428 145236 57492
rect 145300 57428 145301 57492
rect 145235 57427 145301 57428
rect 145422 42125 145482 76467
rect 145419 42124 145485 42125
rect 145419 42060 145420 42124
rect 145484 42060 145485 42124
rect 145419 42059 145485 42060
rect 144499 40764 144565 40765
rect 144499 40700 144500 40764
rect 144564 40700 144565 40764
rect 144499 40699 144565 40700
rect 144315 19956 144381 19957
rect 144315 19892 144316 19956
rect 144380 19892 144381 19956
rect 144315 19891 144381 19892
rect 143211 13700 143277 13701
rect 143211 13636 143212 13700
rect 143276 13636 143277 13700
rect 143211 13635 143277 13636
rect 145606 13565 145666 78099
rect 145794 75454 146414 78000
rect 146526 76669 146586 79595
rect 146523 76668 146589 76669
rect 146523 76604 146524 76668
rect 146588 76604 146589 76668
rect 146523 76603 146589 76604
rect 147075 76668 147141 76669
rect 147075 76604 147076 76668
rect 147140 76604 147141 76668
rect 147075 76603 147141 76604
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145603 13564 145669 13565
rect 145603 13500 145604 13564
rect 145668 13500 145669 13564
rect 145603 13499 145669 13500
rect 142843 7852 142909 7853
rect 142843 7788 142844 7852
rect 142908 7788 142909 7852
rect 142843 7787 142909 7788
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 3454 146414 38898
rect 147078 12341 147138 76603
rect 147075 12340 147141 12341
rect 147075 12276 147076 12340
rect 147140 12276 147141 12340
rect 147075 12275 147141 12276
rect 147262 9213 147322 79867
rect 148179 79796 148245 79797
rect 148179 79732 148180 79796
rect 148244 79732 148245 79796
rect 148179 79731 148245 79732
rect 148731 79796 148797 79797
rect 148731 79732 148732 79796
rect 148796 79732 148797 79796
rect 148731 79731 148797 79732
rect 149651 79796 149717 79797
rect 149651 79732 149652 79796
rect 149716 79732 149717 79796
rect 149651 79731 149717 79732
rect 148182 76533 148242 79731
rect 148547 78300 148613 78301
rect 148547 78236 148548 78300
rect 148612 78236 148613 78300
rect 148547 78235 148613 78236
rect 148363 77892 148429 77893
rect 148363 77828 148364 77892
rect 148428 77828 148429 77892
rect 148363 77827 148429 77828
rect 147443 76532 147509 76533
rect 147443 76468 147444 76532
rect 147508 76468 147509 76532
rect 147443 76467 147509 76468
rect 148179 76532 148245 76533
rect 148179 76468 148180 76532
rect 148244 76468 148245 76532
rect 148179 76467 148245 76468
rect 147259 9212 147325 9213
rect 147259 9148 147260 9212
rect 147324 9148 147325 9212
rect 147259 9147 147325 9148
rect 147446 6357 147506 76467
rect 148366 10709 148426 77827
rect 148550 55861 148610 78235
rect 148547 55860 148613 55861
rect 148547 55796 148548 55860
rect 148612 55796 148613 55860
rect 148547 55795 148613 55796
rect 148734 25669 148794 79731
rect 148731 25668 148797 25669
rect 148731 25604 148732 25668
rect 148796 25604 148797 25668
rect 148731 25603 148797 25604
rect 149654 17237 149714 79731
rect 149838 78165 149898 79867
rect 150942 78165 151002 79867
rect 151491 79796 151557 79797
rect 151491 79732 151492 79796
rect 151556 79732 151557 79796
rect 151491 79731 151557 79732
rect 152043 79796 152109 79797
rect 152043 79732 152044 79796
rect 152108 79732 152109 79796
rect 152043 79731 152109 79732
rect 152595 79796 152661 79797
rect 152595 79732 152596 79796
rect 152660 79732 152661 79796
rect 152595 79731 152661 79732
rect 151307 78708 151373 78709
rect 151307 78644 151308 78708
rect 151372 78644 151373 78708
rect 151307 78643 151373 78644
rect 149835 78164 149901 78165
rect 149835 78100 149836 78164
rect 149900 78100 149901 78164
rect 149835 78099 149901 78100
rect 150019 78164 150085 78165
rect 150019 78100 150020 78164
rect 150084 78100 150085 78164
rect 150019 78099 150085 78100
rect 150939 78164 151005 78165
rect 150939 78100 150940 78164
rect 151004 78100 151005 78164
rect 150939 78099 151005 78100
rect 149835 77892 149901 77893
rect 149835 77828 149836 77892
rect 149900 77828 149901 77892
rect 149835 77827 149901 77828
rect 149651 17236 149717 17237
rect 149651 17172 149652 17236
rect 149716 17172 149717 17236
rect 149651 17171 149717 17172
rect 149838 12205 149898 77827
rect 149835 12204 149901 12205
rect 149835 12140 149836 12204
rect 149900 12140 149901 12204
rect 149835 12139 149901 12140
rect 148363 10708 148429 10709
rect 148363 10644 148364 10708
rect 148428 10644 148429 10708
rect 148363 10643 148429 10644
rect 147443 6356 147509 6357
rect 147443 6292 147444 6356
rect 147508 6292 147509 6356
rect 147443 6291 147509 6292
rect 150022 6221 150082 78099
rect 150294 43954 150914 78000
rect 151310 62933 151370 78643
rect 151307 62932 151373 62933
rect 151307 62868 151308 62932
rect 151372 62868 151373 62932
rect 151307 62867 151373 62868
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 151494 12069 151554 79731
rect 151675 78436 151741 78437
rect 151675 78372 151676 78436
rect 151740 78372 151741 78436
rect 151675 78371 151741 78372
rect 151491 12068 151557 12069
rect 151491 12004 151492 12068
rect 151556 12004 151557 12068
rect 151491 12003 151557 12004
rect 151678 10573 151738 78371
rect 152046 77213 152106 79731
rect 152411 78436 152477 78437
rect 152411 78372 152412 78436
rect 152476 78372 152477 78436
rect 152411 78371 152477 78372
rect 152043 77212 152109 77213
rect 152043 77148 152044 77212
rect 152108 77148 152109 77212
rect 152043 77147 152109 77148
rect 152414 53413 152474 78371
rect 152411 53412 152477 53413
rect 152411 53348 152412 53412
rect 152476 53348 152477 53412
rect 152411 53347 152477 53348
rect 152598 21453 152658 79731
rect 152782 77485 152842 79867
rect 152963 78708 153029 78709
rect 152963 78644 152964 78708
rect 153028 78644 153029 78708
rect 152963 78643 153029 78644
rect 152779 77484 152845 77485
rect 152779 77420 152780 77484
rect 152844 77420 152845 77484
rect 152779 77419 152845 77420
rect 152779 77212 152845 77213
rect 152779 77148 152780 77212
rect 152844 77148 152845 77212
rect 152779 77147 152845 77148
rect 152595 21452 152661 21453
rect 152595 21388 152596 21452
rect 152660 21388 152661 21452
rect 152595 21387 152661 21388
rect 152782 21317 152842 77147
rect 152779 21316 152845 21317
rect 152779 21252 152780 21316
rect 152844 21252 152845 21316
rect 152779 21251 152845 21252
rect 152966 15877 153026 78643
rect 153702 77893 153762 79867
rect 154251 79796 154317 79797
rect 154251 79732 154252 79796
rect 154316 79732 154317 79796
rect 154251 79731 154317 79732
rect 154067 78164 154133 78165
rect 154067 78100 154068 78164
rect 154132 78100 154133 78164
rect 154067 78099 154133 78100
rect 153883 78028 153949 78029
rect 153883 77964 153884 78028
rect 153948 77964 153949 78028
rect 153883 77963 153949 77964
rect 153699 77892 153765 77893
rect 153699 77828 153700 77892
rect 153764 77828 153765 77892
rect 153699 77827 153765 77828
rect 153886 37909 153946 77963
rect 153883 37908 153949 37909
rect 153883 37844 153884 37908
rect 153948 37844 153949 37908
rect 153883 37843 153949 37844
rect 152963 15876 153029 15877
rect 152963 15812 152964 15876
rect 153028 15812 153029 15876
rect 152963 15811 153029 15812
rect 154070 14517 154130 78099
rect 154254 14653 154314 79731
rect 154251 14652 154317 14653
rect 154251 14588 154252 14652
rect 154316 14588 154317 14652
rect 154251 14587 154317 14588
rect 154067 14516 154133 14517
rect 154067 14452 154068 14516
rect 154132 14452 154133 14516
rect 154067 14451 154133 14452
rect 154438 13429 154498 79867
rect 154622 78029 154682 79867
rect 155358 78165 155418 79867
rect 156275 79796 156341 79797
rect 156275 79732 156276 79796
rect 156340 79732 156341 79796
rect 156275 79731 156341 79732
rect 155723 79660 155789 79661
rect 155723 79596 155724 79660
rect 155788 79596 155789 79660
rect 155723 79595 155789 79596
rect 155355 78164 155421 78165
rect 155355 78100 155356 78164
rect 155420 78100 155421 78164
rect 155355 78099 155421 78100
rect 154619 78028 154685 78029
rect 154619 77964 154620 78028
rect 154684 77964 154685 78028
rect 154619 77963 154685 77964
rect 154794 48454 155414 78000
rect 155539 77892 155605 77893
rect 155539 77828 155540 77892
rect 155604 77828 155605 77892
rect 155539 77827 155605 77828
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154435 13428 154501 13429
rect 154435 13364 154436 13428
rect 154500 13364 154501 13428
rect 154435 13363 154501 13364
rect 154794 12454 155414 47898
rect 155542 44845 155602 77827
rect 155539 44844 155605 44845
rect 155539 44780 155540 44844
rect 155604 44780 155605 44844
rect 155539 44779 155605 44780
rect 155726 26893 155786 79595
rect 156278 78709 156338 79731
rect 156827 79660 156893 79661
rect 156827 79596 156828 79660
rect 156892 79596 156893 79660
rect 156827 79595 156893 79596
rect 157195 79660 157261 79661
rect 157195 79596 157196 79660
rect 157260 79596 157261 79660
rect 157195 79595 157261 79596
rect 156275 78708 156341 78709
rect 156275 78644 156276 78708
rect 156340 78644 156341 78708
rect 156275 78643 156341 78644
rect 156643 78708 156709 78709
rect 156643 78644 156644 78708
rect 156708 78644 156709 78708
rect 156643 78643 156709 78644
rect 155723 26892 155789 26893
rect 155723 26828 155724 26892
rect 155788 26828 155789 26892
rect 155723 26827 155789 26828
rect 156646 24309 156706 78643
rect 156830 29613 156890 79595
rect 157198 70410 157258 79595
rect 157382 78437 157442 79867
rect 157931 79796 157997 79797
rect 157931 79732 157932 79796
rect 157996 79732 157997 79796
rect 157931 79731 157997 79732
rect 157379 78436 157445 78437
rect 157379 78372 157380 78436
rect 157444 78372 157445 78436
rect 157379 78371 157445 78372
rect 157934 77485 157994 79731
rect 157931 77484 157997 77485
rect 157931 77420 157932 77484
rect 157996 77420 157997 77484
rect 157931 77419 157997 77420
rect 157931 77212 157997 77213
rect 157931 77148 157932 77212
rect 157996 77148 157997 77212
rect 157931 77147 157997 77148
rect 157014 70350 157258 70410
rect 156827 29612 156893 29613
rect 156827 29548 156828 29612
rect 156892 29548 156893 29612
rect 156827 29547 156893 29548
rect 156643 24308 156709 24309
rect 156643 24244 156644 24308
rect 156708 24244 156709 24308
rect 156643 24243 156709 24244
rect 157014 24173 157074 70350
rect 157934 48925 157994 77147
rect 157931 48924 157997 48925
rect 157931 48860 157932 48924
rect 157996 48860 157997 48924
rect 157931 48859 157997 48860
rect 157011 24172 157077 24173
rect 157011 24108 157012 24172
rect 157076 24108 157077 24172
rect 157011 24107 157077 24108
rect 158118 22677 158178 79867
rect 158299 79796 158365 79797
rect 158299 79732 158300 79796
rect 158364 79732 158365 79796
rect 158299 79731 158365 79732
rect 158115 22676 158181 22677
rect 158115 22612 158116 22676
rect 158180 22612 158181 22676
rect 158115 22611 158181 22612
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 151675 10572 151741 10573
rect 151675 10508 151676 10572
rect 151740 10508 151741 10572
rect 151675 10507 151741 10508
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150019 6220 150085 6221
rect 150019 6156 150020 6220
rect 150084 6156 150085 6220
rect 150019 6155 150085 6156
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 -2266 155414 11898
rect 158302 7717 158362 79731
rect 158483 79660 158549 79661
rect 158483 79596 158484 79660
rect 158548 79596 158549 79660
rect 158483 79595 158549 79596
rect 158299 7716 158365 7717
rect 158299 7652 158300 7716
rect 158364 7652 158365 7716
rect 158299 7651 158365 7652
rect 158486 4997 158546 79595
rect 158670 77621 158730 79867
rect 159035 79660 159101 79661
rect 159035 79596 159036 79660
rect 159100 79596 159101 79660
rect 159035 79595 159101 79596
rect 158667 77620 158733 77621
rect 158667 77556 158668 77620
rect 158732 77556 158733 77620
rect 158667 77555 158733 77556
rect 159038 76533 159098 79595
rect 159958 78709 160018 79867
rect 159955 78708 160021 78709
rect 159955 78644 159956 78708
rect 160020 78644 160021 78708
rect 159955 78643 160021 78644
rect 159035 76532 159101 76533
rect 159035 76468 159036 76532
rect 159100 76468 159101 76532
rect 159035 76467 159101 76468
rect 159035 75308 159101 75309
rect 159035 75244 159036 75308
rect 159100 75244 159101 75308
rect 159035 75243 159101 75244
rect 158851 75172 158917 75173
rect 158851 75108 158852 75172
rect 158916 75108 158917 75172
rect 158851 75107 158917 75108
rect 158854 10437 158914 75107
rect 158851 10436 158917 10437
rect 158851 10372 158852 10436
rect 158916 10372 158917 10436
rect 158851 10371 158917 10372
rect 159038 10301 159098 75243
rect 159294 52954 159914 78000
rect 160142 75173 160202 80003
rect 160507 79932 160573 79933
rect 160507 79868 160508 79932
rect 160572 79868 160573 79932
rect 161059 79932 161125 79933
rect 161059 79930 161060 79932
rect 160507 79867 160573 79868
rect 160878 79870 161060 79930
rect 160510 78437 160570 79867
rect 160507 78436 160573 78437
rect 160507 78372 160508 78436
rect 160572 78372 160573 78436
rect 160507 78371 160573 78372
rect 160139 75172 160205 75173
rect 160139 75108 160140 75172
rect 160204 75108 160205 75172
rect 160139 75107 160205 75108
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159035 10300 159101 10301
rect 159035 10236 159036 10300
rect 159100 10236 159101 10300
rect 159035 10235 159101 10236
rect 158483 4996 158549 4997
rect 158483 4932 158484 4996
rect 158548 4932 158549 4996
rect 158483 4931 158549 4932
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 -3226 159914 16398
rect 160878 13293 160938 79870
rect 161059 79868 161060 79870
rect 161124 79868 161125 79932
rect 161059 79867 161125 79868
rect 161059 79796 161125 79797
rect 161059 79732 161060 79796
rect 161124 79732 161125 79796
rect 161059 79731 161125 79732
rect 161795 79796 161861 79797
rect 161795 79732 161796 79796
rect 161860 79732 161861 79796
rect 161795 79731 161861 79732
rect 161062 54501 161122 79731
rect 161798 77310 161858 79731
rect 161982 78981 162042 80139
rect 162715 79932 162781 79933
rect 162715 79868 162716 79932
rect 162780 79868 162781 79932
rect 162715 79867 162781 79868
rect 163451 79932 163517 79933
rect 163451 79868 163452 79932
rect 163516 79868 163517 79932
rect 163451 79867 163517 79868
rect 165107 79932 165173 79933
rect 165107 79868 165108 79932
rect 165172 79868 165173 79932
rect 165107 79867 165173 79868
rect 166395 79932 166461 79933
rect 166395 79868 166396 79932
rect 166460 79868 166461 79932
rect 166395 79867 166461 79868
rect 166763 79932 166829 79933
rect 166763 79868 166764 79932
rect 166828 79868 166829 79932
rect 167867 79932 167933 79933
rect 167867 79930 167868 79932
rect 166763 79867 166829 79868
rect 167502 79870 167868 79930
rect 162347 79796 162413 79797
rect 162347 79732 162348 79796
rect 162412 79732 162413 79796
rect 162347 79731 162413 79732
rect 161979 78980 162045 78981
rect 161979 78916 161980 78980
rect 162044 78916 162045 78980
rect 161979 78915 162045 78916
rect 161614 77250 161858 77310
rect 161614 75989 161674 77250
rect 161611 75988 161677 75989
rect 161611 75924 161612 75988
rect 161676 75924 161677 75988
rect 161611 75923 161677 75924
rect 162163 75036 162229 75037
rect 162163 74972 162164 75036
rect 162228 74972 162229 75036
rect 162163 74971 162229 74972
rect 161059 54500 161125 54501
rect 161059 54436 161060 54500
rect 161124 54436 161125 54500
rect 161059 54435 161125 54436
rect 160875 13292 160941 13293
rect 160875 13228 160876 13292
rect 160940 13228 160941 13292
rect 160875 13227 160941 13228
rect 162166 9077 162226 74971
rect 162350 11797 162410 79731
rect 162531 79116 162597 79117
rect 162531 79052 162532 79116
rect 162596 79052 162597 79116
rect 162531 79051 162597 79052
rect 162534 11933 162594 79051
rect 162718 78709 162778 79867
rect 162715 78708 162781 78709
rect 162715 78644 162716 78708
rect 162780 78644 162781 78708
rect 162715 78643 162781 78644
rect 163454 57221 163514 79867
rect 163635 79796 163701 79797
rect 163635 79732 163636 79796
rect 163700 79732 163701 79796
rect 163635 79731 163701 79732
rect 163451 57220 163517 57221
rect 163451 57156 163452 57220
rect 163516 57156 163517 57220
rect 163451 57155 163517 57156
rect 162531 11932 162597 11933
rect 162531 11868 162532 11932
rect 162596 11868 162597 11932
rect 162531 11867 162597 11868
rect 162347 11796 162413 11797
rect 162347 11732 162348 11796
rect 162412 11732 162413 11796
rect 162347 11731 162413 11732
rect 162163 9076 162229 9077
rect 162163 9012 162164 9076
rect 162228 9012 162229 9076
rect 162163 9011 162229 9012
rect 163638 4861 163698 79731
rect 164739 79660 164805 79661
rect 164739 79596 164740 79660
rect 164804 79596 164805 79660
rect 164739 79595 164805 79596
rect 164923 79660 164989 79661
rect 164923 79596 164924 79660
rect 164988 79596 164989 79660
rect 164923 79595 164989 79596
rect 163794 57454 164414 78000
rect 164742 75173 164802 79595
rect 164739 75172 164805 75173
rect 164739 75108 164740 75172
rect 164804 75108 164805 75172
rect 164739 75107 164805 75108
rect 164926 64157 164986 79595
rect 164923 64156 164989 64157
rect 164923 64092 164924 64156
rect 164988 64092 164989 64156
rect 164923 64091 164989 64092
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 165110 53277 165170 79867
rect 165475 79796 165541 79797
rect 165475 79732 165476 79796
rect 165540 79732 165541 79796
rect 165475 79731 165541 79732
rect 165291 75988 165357 75989
rect 165291 75924 165292 75988
rect 165356 75924 165357 75988
rect 165291 75923 165357 75924
rect 165107 53276 165173 53277
rect 165107 53212 165108 53276
rect 165172 53212 165173 53276
rect 165107 53211 165173 53212
rect 165294 40629 165354 75923
rect 165291 40628 165357 40629
rect 165291 40564 165292 40628
rect 165356 40564 165357 40628
rect 165291 40563 165357 40564
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163635 4860 163701 4861
rect 163635 4796 163636 4860
rect 163700 4796 163701 4860
rect 163635 4795 163701 4796
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 -4186 164414 20898
rect 165478 13157 165538 79731
rect 166398 79389 166458 79867
rect 166395 79388 166461 79389
rect 166395 79324 166396 79388
rect 166460 79324 166461 79388
rect 166395 79323 166461 79324
rect 166211 77892 166277 77893
rect 166211 77828 166212 77892
rect 166276 77828 166277 77892
rect 166211 77827 166277 77828
rect 166214 69597 166274 77827
rect 166395 77484 166461 77485
rect 166395 77420 166396 77484
rect 166460 77420 166461 77484
rect 166395 77419 166461 77420
rect 166211 69596 166277 69597
rect 166211 69532 166212 69596
rect 166276 69532 166277 69596
rect 166211 69531 166277 69532
rect 166398 51781 166458 77419
rect 166579 77348 166645 77349
rect 166579 77284 166580 77348
rect 166644 77284 166645 77348
rect 166579 77283 166645 77284
rect 166395 51780 166461 51781
rect 166395 51716 166396 51780
rect 166460 51716 166461 51780
rect 166395 51715 166461 51716
rect 166582 39269 166642 77283
rect 166579 39268 166645 39269
rect 166579 39204 166580 39268
rect 166644 39204 166645 39268
rect 166579 39203 166645 39204
rect 166766 25533 166826 79867
rect 167315 79388 167381 79389
rect 167315 79324 167316 79388
rect 167380 79324 167381 79388
rect 167315 79323 167381 79324
rect 167318 75989 167378 79323
rect 167315 75988 167381 75989
rect 167315 75924 167316 75988
rect 167380 75924 167381 75988
rect 167315 75923 167381 75924
rect 167502 62797 167562 79870
rect 167867 79868 167868 79870
rect 167932 79868 167933 79932
rect 167867 79867 167933 79868
rect 167683 79660 167749 79661
rect 167683 79596 167684 79660
rect 167748 79596 167749 79660
rect 167683 79595 167749 79596
rect 167499 62796 167565 62797
rect 167499 62732 167500 62796
rect 167564 62732 167565 62796
rect 167499 62731 167565 62732
rect 167686 46205 167746 79595
rect 167867 79388 167933 79389
rect 167867 79324 167868 79388
rect 167932 79324 167933 79388
rect 167867 79323 167933 79324
rect 167683 46204 167749 46205
rect 167683 46140 167684 46204
rect 167748 46140 167749 46204
rect 167683 46139 167749 46140
rect 166763 25532 166829 25533
rect 166763 25468 166764 25532
rect 166828 25468 166829 25532
rect 166763 25467 166829 25468
rect 167870 18597 167930 79323
rect 168054 78709 168114 80547
rect 172283 80340 172349 80341
rect 172283 80276 172284 80340
rect 172348 80276 172349 80340
rect 172283 80275 172349 80276
rect 168419 79932 168485 79933
rect 168419 79868 168420 79932
rect 168484 79868 168485 79932
rect 168419 79867 168485 79868
rect 168971 79932 169037 79933
rect 168971 79868 168972 79932
rect 169036 79868 169037 79932
rect 168971 79867 169037 79868
rect 169523 79932 169589 79933
rect 169523 79868 169524 79932
rect 169588 79868 169589 79932
rect 169523 79867 169589 79868
rect 169891 79932 169957 79933
rect 169891 79868 169892 79932
rect 169956 79868 169957 79932
rect 169891 79867 169957 79868
rect 170443 79932 170509 79933
rect 170443 79868 170444 79932
rect 170508 79868 170509 79932
rect 170443 79867 170509 79868
rect 170811 79932 170877 79933
rect 170811 79868 170812 79932
rect 170876 79868 170877 79932
rect 170811 79867 170877 79868
rect 171179 79932 171245 79933
rect 171179 79868 171180 79932
rect 171244 79868 171245 79932
rect 171179 79867 171245 79868
rect 171731 79932 171797 79933
rect 171731 79868 171732 79932
rect 171796 79868 171797 79932
rect 171731 79867 171797 79868
rect 171915 79932 171981 79933
rect 171915 79868 171916 79932
rect 171980 79868 171981 79932
rect 172145 79932 172211 79933
rect 172145 79930 172146 79932
rect 171915 79867 171981 79868
rect 172102 79868 172146 79930
rect 172210 79868 172211 79932
rect 172102 79867 172211 79868
rect 168051 78708 168117 78709
rect 168051 78644 168052 78708
rect 168116 78644 168117 78708
rect 168051 78643 168117 78644
rect 168422 78165 168482 79867
rect 168974 79389 169034 79867
rect 168787 79388 168853 79389
rect 168787 79324 168788 79388
rect 168852 79324 168853 79388
rect 168787 79323 168853 79324
rect 168971 79388 169037 79389
rect 168971 79324 168972 79388
rect 169036 79324 169037 79388
rect 168971 79323 169037 79324
rect 168790 78301 168850 79323
rect 169526 78690 169586 79867
rect 169894 79389 169954 79867
rect 169891 79388 169957 79389
rect 169891 79324 169892 79388
rect 169956 79324 169957 79388
rect 169891 79323 169957 79324
rect 170259 79388 170325 79389
rect 170259 79324 170260 79388
rect 170324 79324 170325 79388
rect 170259 79323 170325 79324
rect 169342 78630 169586 78690
rect 168787 78300 168853 78301
rect 168787 78236 168788 78300
rect 168852 78236 168853 78300
rect 168787 78235 168853 78236
rect 168419 78164 168485 78165
rect 168419 78100 168420 78164
rect 168484 78100 168485 78164
rect 168419 78099 168485 78100
rect 168051 75988 168117 75989
rect 168051 75924 168052 75988
rect 168116 75924 168117 75988
rect 168051 75923 168117 75924
rect 167867 18596 167933 18597
rect 167867 18532 167868 18596
rect 167932 18532 167933 18596
rect 167867 18531 167933 18532
rect 165475 13156 165541 13157
rect 165475 13092 165476 13156
rect 165540 13092 165541 13156
rect 165475 13091 165541 13092
rect 168054 7581 168114 75923
rect 168294 61954 168914 78000
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168051 7580 168117 7581
rect 168051 7516 168052 7580
rect 168116 7516 168117 7580
rect 168051 7515 168117 7516
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 -5146 168914 25398
rect 169342 13021 169402 78630
rect 170262 78301 170322 79323
rect 170259 78300 170325 78301
rect 170259 78236 170260 78300
rect 170324 78236 170325 78300
rect 170259 78235 170325 78236
rect 169339 13020 169405 13021
rect 169339 12956 169340 13020
rect 169404 12956 169405 13020
rect 169339 12955 169405 12956
rect 170446 8941 170506 79867
rect 170627 77484 170693 77485
rect 170627 77420 170628 77484
rect 170692 77420 170693 77484
rect 170627 77419 170693 77420
rect 170630 53141 170690 77419
rect 170627 53140 170693 53141
rect 170627 53076 170628 53140
rect 170692 53076 170693 53140
rect 170627 53075 170693 53076
rect 170814 11661 170874 79867
rect 171182 79389 171242 79867
rect 171179 79388 171245 79389
rect 171179 79324 171180 79388
rect 171244 79324 171245 79388
rect 171179 79323 171245 79324
rect 170995 78708 171061 78709
rect 170995 78644 170996 78708
rect 171060 78644 171061 78708
rect 170995 78643 171061 78644
rect 170998 73813 171058 78643
rect 171547 78436 171613 78437
rect 171547 78372 171548 78436
rect 171612 78372 171613 78436
rect 171547 78371 171613 78372
rect 170995 73812 171061 73813
rect 170995 73748 170996 73812
rect 171060 73748 171061 73812
rect 170995 73747 171061 73748
rect 171550 59941 171610 78371
rect 171734 77757 171794 79867
rect 171918 78573 171978 79867
rect 171915 78572 171981 78573
rect 171915 78508 171916 78572
rect 171980 78508 171981 78572
rect 171915 78507 171981 78508
rect 172102 78165 172162 79867
rect 172286 78709 172346 80275
rect 186294 79954 186914 115398
rect 172467 79932 172533 79933
rect 172467 79868 172468 79932
rect 172532 79868 172533 79932
rect 172467 79867 172533 79868
rect 173755 79932 173821 79933
rect 173755 79868 173756 79932
rect 173820 79868 173821 79932
rect 173755 79867 173821 79868
rect 172470 78709 172530 79867
rect 172835 79660 172901 79661
rect 172835 79596 172836 79660
rect 172900 79596 172901 79660
rect 172835 79595 172901 79596
rect 172838 79386 172898 79595
rect 173203 79388 173269 79389
rect 173203 79386 173204 79388
rect 172838 79326 173204 79386
rect 173203 79324 173204 79326
rect 173268 79324 173269 79388
rect 173203 79323 173269 79324
rect 173758 79253 173818 79867
rect 173939 79796 174005 79797
rect 173939 79732 173940 79796
rect 174004 79732 174005 79796
rect 173939 79731 174005 79732
rect 173942 79525 174002 79731
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 173939 79524 174005 79525
rect 173939 79460 173940 79524
rect 174004 79460 174005 79524
rect 173939 79459 174005 79460
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 173755 79252 173821 79253
rect 173755 79188 173756 79252
rect 173820 79188 173821 79252
rect 173755 79187 173821 79188
rect 172283 78708 172349 78709
rect 172283 78644 172284 78708
rect 172348 78644 172349 78708
rect 172283 78643 172349 78644
rect 172467 78708 172533 78709
rect 172467 78644 172468 78708
rect 172532 78644 172533 78708
rect 172467 78643 172533 78644
rect 172099 78164 172165 78165
rect 172099 78100 172100 78164
rect 172164 78100 172165 78164
rect 172099 78099 172165 78100
rect 171731 77756 171797 77757
rect 171731 77692 171732 77756
rect 171796 77692 171797 77756
rect 171731 77691 171797 77692
rect 172283 77620 172349 77621
rect 172283 77556 172284 77620
rect 172348 77556 172349 77620
rect 172283 77555 172349 77556
rect 171731 75988 171797 75989
rect 171731 75924 171732 75988
rect 171796 75924 171797 75988
rect 171731 75923 171797 75924
rect 171547 59940 171613 59941
rect 171547 59876 171548 59940
rect 171612 59876 171613 59940
rect 171547 59875 171613 59876
rect 171734 31789 171794 75923
rect 172286 57357 172346 77555
rect 172794 66454 173414 78000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172283 57356 172349 57357
rect 172283 57292 172284 57356
rect 172348 57292 172349 57356
rect 172283 57291 172349 57292
rect 171731 31788 171797 31789
rect 171731 31724 171732 31788
rect 171796 31724 171797 31788
rect 171731 31723 171797 31724
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 170811 11660 170877 11661
rect 170811 11596 170812 11660
rect 170876 11596 170877 11660
rect 170811 11595 170877 11596
rect 170443 8940 170509 8941
rect 170443 8876 170444 8940
rect 170508 8876 170509 8940
rect 170443 8875 170509 8876
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 70954 177914 78000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 75454 182414 78000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 228453 191414 228484
rect 190794 228217 190826 228453
rect 191062 228217 191146 228453
rect 191382 228217 191414 228453
rect 190794 228133 191414 228217
rect 190794 227897 190826 228133
rect 191062 227897 191146 228133
rect 191382 227897 191414 228133
rect 190794 192454 191414 227897
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 196954 195914 228484
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 201454 200414 228484
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 205954 204914 228484
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 210454 209414 228484
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 214954 213914 228484
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 219454 218414 228484
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 223954 222914 228484
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 228453 227414 228484
rect 226794 228217 226826 228453
rect 227062 228217 227146 228453
rect 227382 228217 227414 228453
rect 226794 228133 227414 228217
rect 226794 227897 226826 228133
rect 227062 227897 227146 228133
rect 227382 227897 227414 228133
rect 226794 192454 227414 227897
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 196954 231914 228484
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 201454 236414 228484
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 205954 240914 228484
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 210454 245414 228484
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 214954 249914 228484
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 219454 254414 228484
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 223954 258914 228484
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 228453 263414 228484
rect 262794 228217 262826 228453
rect 263062 228217 263146 228453
rect 263382 228217 263414 228453
rect 262794 228133 263414 228217
rect 262794 227897 262826 228133
rect 263062 227897 263146 228133
rect 263382 227897 263414 228133
rect 262794 192454 263414 227897
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 196954 267914 228484
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 201454 272414 228484
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 205954 276914 228484
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 210454 281414 228484
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 214954 285914 228484
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 219454 290414 228484
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 223954 294914 228484
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 228453 299414 228484
rect 298794 228217 298826 228453
rect 299062 228217 299146 228453
rect 299382 228217 299414 228453
rect 298794 228133 299414 228217
rect 298794 227897 298826 228133
rect 299062 227897 299146 228133
rect 299382 227897 299414 228133
rect 298794 192454 299414 227897
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 196954 303914 228484
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 201454 308414 228484
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 205954 312914 228484
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 210454 317414 228484
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 214954 321914 228484
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 219454 326414 228484
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 223954 330914 228484
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 228453 335414 228484
rect 334794 228217 334826 228453
rect 335062 228217 335146 228453
rect 335382 228217 335414 228453
rect 334794 228133 335414 228217
rect 334794 227897 334826 228133
rect 335062 227897 335146 228133
rect 335382 227897 335414 228133
rect 334794 192454 335414 227897
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 196954 339914 228484
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 201454 344414 228484
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 205954 348914 228484
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 210454 353414 228484
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 214954 357914 228484
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 219454 362414 228484
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 223954 366914 228484
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 228453 371414 228484
rect 370794 228217 370826 228453
rect 371062 228217 371146 228453
rect 371382 228217 371414 228453
rect 370794 228133 371414 228217
rect 370794 227897 370826 228133
rect 371062 227897 371146 228133
rect 371382 227897 371414 228133
rect 370794 192454 371414 227897
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 196954 375914 228484
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 201454 380414 228484
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 205954 384914 228484
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 210454 389414 228484
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 214954 393914 228484
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 396582 78165 396642 696899
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 248684 398414 254898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 397794 219454 398414 228484
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 396579 78164 396645 78165
rect 396579 78100 396580 78164
rect 396644 78100 396645 78164
rect 396579 78099 396645 78100
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 65342 246067 65578 246303
rect 65662 246067 65898 246303
rect 65982 246067 66218 246303
rect 66302 246067 66538 246303
rect 66622 246067 66858 246303
rect 66942 246067 67178 246303
rect 67262 246067 67498 246303
rect 67582 246067 67818 246303
rect 67902 246067 68138 246303
rect 68222 246067 68458 246303
rect 68542 246067 68778 246303
rect 68862 246067 69098 246303
rect 69182 246067 69418 246303
rect 69502 246067 69738 246303
rect 69822 246067 70058 246303
rect 65462 241717 65698 241953
rect 65782 241717 66018 241953
rect 66102 241717 66338 241953
rect 66422 241717 66658 241953
rect 66742 241717 66978 241953
rect 67062 241717 67298 241953
rect 67382 241717 67618 241953
rect 67702 241717 67938 241953
rect 68022 241717 68258 241953
rect 68342 241717 68578 241953
rect 68662 241717 68898 241953
rect 68982 241717 69218 241953
rect 69302 241717 69538 241953
rect 69622 241717 69858 241953
rect 69942 241717 70178 241953
rect 70262 241717 70498 241953
rect 70582 241717 70818 241953
rect 70902 241717 71138 241953
rect 65462 241397 65698 241633
rect 65782 241397 66018 241633
rect 66102 241397 66338 241633
rect 66422 241397 66658 241633
rect 66742 241397 66978 241633
rect 67062 241397 67298 241633
rect 67382 241397 67618 241633
rect 67702 241397 67938 241633
rect 68022 241397 68258 241633
rect 68342 241397 68578 241633
rect 68662 241397 68898 241633
rect 68982 241397 69218 241633
rect 69302 241397 69538 241633
rect 69622 241397 69858 241633
rect 69942 241397 70178 241633
rect 70262 241397 70498 241633
rect 70582 241397 70818 241633
rect 70902 241397 71138 241633
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 228217 47062 228453
rect 47146 228217 47382 228453
rect 46826 227897 47062 228133
rect 47146 227897 47382 228133
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 228217 83062 228453
rect 83146 228217 83382 228453
rect 82826 227897 83062 228133
rect 83146 227897 83382 228133
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 118826 228217 119062 228453
rect 119146 228217 119382 228453
rect 118826 227897 119062 228133
rect 119146 227897 119382 228133
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 136036 205718 136272 205954
rect 136356 205718 136592 205954
rect 136676 205718 136912 205954
rect 136996 205718 137232 205954
rect 137316 205718 137552 205954
rect 137636 205718 137872 205954
rect 137956 205718 138192 205954
rect 138276 205718 138512 205954
rect 138596 205718 138832 205954
rect 138916 205718 139152 205954
rect 139236 205718 139472 205954
rect 139556 205718 139792 205954
rect 139876 205718 140112 205954
rect 140196 205718 140432 205954
rect 140516 205718 140752 205954
rect 140836 205718 141072 205954
rect 141156 205718 141392 205954
rect 141476 205718 141712 205954
rect 141796 205718 142032 205954
rect 142116 205718 142352 205954
rect 142436 205718 142672 205954
rect 142756 205718 142992 205954
rect 143076 205718 143312 205954
rect 143396 205718 143632 205954
rect 143716 205718 143952 205954
rect 144036 205718 144272 205954
rect 144356 205718 144592 205954
rect 144676 205718 144912 205954
rect 144996 205718 145232 205954
rect 145316 205718 145552 205954
rect 145636 205718 145872 205954
rect 145956 205718 146192 205954
rect 146276 205718 146512 205954
rect 146596 205718 146832 205954
rect 146916 205718 147152 205954
rect 147236 205718 147472 205954
rect 147556 205718 147792 205954
rect 147876 205718 148112 205954
rect 148196 205718 148432 205954
rect 148516 205718 148752 205954
rect 148836 205718 149072 205954
rect 149156 205718 149392 205954
rect 149476 205718 149712 205954
rect 149796 205718 150032 205954
rect 150116 205718 150352 205954
rect 150436 205718 150672 205954
rect 150756 205718 150992 205954
rect 151076 205718 151312 205954
rect 151396 205718 151632 205954
rect 151716 205718 151952 205954
rect 152036 205718 152272 205954
rect 152356 205718 152592 205954
rect 152676 205718 152912 205954
rect 152996 205718 153232 205954
rect 153316 205718 153552 205954
rect 153636 205718 153872 205954
rect 153956 205718 154192 205954
rect 154276 205718 154512 205954
rect 154596 205718 154832 205954
rect 154916 205718 155152 205954
rect 155236 205718 155472 205954
rect 155556 205718 155792 205954
rect 155876 205718 156112 205954
rect 156196 205718 156432 205954
rect 156516 205718 156752 205954
rect 156836 205718 157072 205954
rect 157156 205718 157392 205954
rect 157476 205718 157712 205954
rect 157796 205718 158032 205954
rect 158116 205718 158352 205954
rect 158436 205718 158672 205954
rect 158756 205718 158992 205954
rect 159076 205718 159312 205954
rect 159396 205718 159632 205954
rect 159716 205718 159952 205954
rect 160036 205718 160272 205954
rect 160356 205718 160592 205954
rect 160676 205718 160912 205954
rect 160996 205718 161232 205954
rect 161316 205718 161552 205954
rect 161636 205718 161872 205954
rect 161956 205718 162192 205954
rect 162276 205718 162512 205954
rect 162596 205718 162832 205954
rect 162916 205718 163152 205954
rect 163236 205718 163472 205954
rect 163556 205718 163792 205954
rect 163876 205718 164112 205954
rect 164196 205718 164432 205954
rect 164516 205718 164752 205954
rect 164836 205718 165072 205954
rect 165156 205718 165392 205954
rect 136036 205398 136272 205634
rect 136356 205398 136592 205634
rect 136676 205398 136912 205634
rect 136996 205398 137232 205634
rect 137316 205398 137552 205634
rect 137636 205398 137872 205634
rect 137956 205398 138192 205634
rect 138276 205398 138512 205634
rect 138596 205398 138832 205634
rect 138916 205398 139152 205634
rect 139236 205398 139472 205634
rect 139556 205398 139792 205634
rect 139876 205398 140112 205634
rect 140196 205398 140432 205634
rect 140516 205398 140752 205634
rect 140836 205398 141072 205634
rect 141156 205398 141392 205634
rect 141476 205398 141712 205634
rect 141796 205398 142032 205634
rect 142116 205398 142352 205634
rect 142436 205398 142672 205634
rect 142756 205398 142992 205634
rect 143076 205398 143312 205634
rect 143396 205398 143632 205634
rect 143716 205398 143952 205634
rect 144036 205398 144272 205634
rect 144356 205398 144592 205634
rect 144676 205398 144912 205634
rect 144996 205398 145232 205634
rect 145316 205398 145552 205634
rect 145636 205398 145872 205634
rect 145956 205398 146192 205634
rect 146276 205398 146512 205634
rect 146596 205398 146832 205634
rect 146916 205398 147152 205634
rect 147236 205398 147472 205634
rect 147556 205398 147792 205634
rect 147876 205398 148112 205634
rect 148196 205398 148432 205634
rect 148516 205398 148752 205634
rect 148836 205398 149072 205634
rect 149156 205398 149392 205634
rect 149476 205398 149712 205634
rect 149796 205398 150032 205634
rect 150116 205398 150352 205634
rect 150436 205398 150672 205634
rect 150756 205398 150992 205634
rect 151076 205398 151312 205634
rect 151396 205398 151632 205634
rect 151716 205398 151952 205634
rect 152036 205398 152272 205634
rect 152356 205398 152592 205634
rect 152676 205398 152912 205634
rect 152996 205398 153232 205634
rect 153316 205398 153552 205634
rect 153636 205398 153872 205634
rect 153956 205398 154192 205634
rect 154276 205398 154512 205634
rect 154596 205398 154832 205634
rect 154916 205398 155152 205634
rect 155236 205398 155472 205634
rect 155556 205398 155792 205634
rect 155876 205398 156112 205634
rect 156196 205398 156432 205634
rect 156516 205398 156752 205634
rect 156836 205398 157072 205634
rect 157156 205398 157392 205634
rect 157476 205398 157712 205634
rect 157796 205398 158032 205634
rect 158116 205398 158352 205634
rect 158436 205398 158672 205634
rect 158756 205398 158992 205634
rect 159076 205398 159312 205634
rect 159396 205398 159632 205634
rect 159716 205398 159952 205634
rect 160036 205398 160272 205634
rect 160356 205398 160592 205634
rect 160676 205398 160912 205634
rect 160996 205398 161232 205634
rect 161316 205398 161552 205634
rect 161636 205398 161872 205634
rect 161956 205398 162192 205634
rect 162276 205398 162512 205634
rect 162596 205398 162832 205634
rect 162916 205398 163152 205634
rect 163236 205398 163472 205634
rect 163556 205398 163792 205634
rect 163876 205398 164112 205634
rect 164196 205398 164432 205634
rect 164516 205398 164752 205634
rect 164836 205398 165072 205634
rect 165156 205398 165392 205634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 137376 201218 137612 201454
rect 137696 201218 137932 201454
rect 138016 201218 138252 201454
rect 138336 201218 138572 201454
rect 138656 201218 138892 201454
rect 138976 201218 139212 201454
rect 139296 201218 139532 201454
rect 139616 201218 139852 201454
rect 139936 201218 140172 201454
rect 140256 201218 140492 201454
rect 140576 201218 140812 201454
rect 140896 201218 141132 201454
rect 141216 201218 141452 201454
rect 141536 201218 141772 201454
rect 141856 201218 142092 201454
rect 142176 201218 142412 201454
rect 142496 201218 142732 201454
rect 142816 201218 143052 201454
rect 143136 201218 143372 201454
rect 143456 201218 143692 201454
rect 143776 201218 144012 201454
rect 144096 201218 144332 201454
rect 144416 201218 144652 201454
rect 144736 201218 144972 201454
rect 145056 201218 145292 201454
rect 145376 201218 145612 201454
rect 145696 201218 145932 201454
rect 146016 201218 146252 201454
rect 146336 201218 146572 201454
rect 146656 201218 146892 201454
rect 146976 201218 147212 201454
rect 147296 201218 147532 201454
rect 147616 201218 147852 201454
rect 147936 201218 148172 201454
rect 148256 201218 148492 201454
rect 148576 201218 148812 201454
rect 148896 201218 149132 201454
rect 149216 201218 149452 201454
rect 149536 201218 149772 201454
rect 149856 201218 150092 201454
rect 150176 201218 150412 201454
rect 150496 201218 150732 201454
rect 150816 201218 151052 201454
rect 151136 201218 151372 201454
rect 151456 201218 151692 201454
rect 151776 201218 152012 201454
rect 152096 201218 152332 201454
rect 152416 201218 152652 201454
rect 152736 201218 152972 201454
rect 153056 201218 153292 201454
rect 153376 201218 153612 201454
rect 153696 201218 153932 201454
rect 154016 201218 154252 201454
rect 154336 201218 154572 201454
rect 154656 201218 154892 201454
rect 154976 201218 155212 201454
rect 155296 201218 155532 201454
rect 155616 201218 155852 201454
rect 155936 201218 156172 201454
rect 156256 201218 156492 201454
rect 156576 201218 156812 201454
rect 156896 201218 157132 201454
rect 157216 201218 157452 201454
rect 157536 201218 157772 201454
rect 157856 201218 158092 201454
rect 158176 201218 158412 201454
rect 158496 201218 158732 201454
rect 158816 201218 159052 201454
rect 159136 201218 159372 201454
rect 159456 201218 159692 201454
rect 159776 201218 160012 201454
rect 160096 201218 160332 201454
rect 160416 201218 160652 201454
rect 160736 201218 160972 201454
rect 161056 201218 161292 201454
rect 161376 201218 161612 201454
rect 161696 201218 161932 201454
rect 162016 201218 162252 201454
rect 162336 201218 162572 201454
rect 162656 201218 162892 201454
rect 162976 201218 163212 201454
rect 163296 201218 163532 201454
rect 163616 201218 163852 201454
rect 163936 201218 164172 201454
rect 164256 201218 164492 201454
rect 164576 201218 164812 201454
rect 164896 201218 165132 201454
rect 165216 201218 165452 201454
rect 137376 200898 137612 201134
rect 137696 200898 137932 201134
rect 138016 200898 138252 201134
rect 138336 200898 138572 201134
rect 138656 200898 138892 201134
rect 138976 200898 139212 201134
rect 139296 200898 139532 201134
rect 139616 200898 139852 201134
rect 139936 200898 140172 201134
rect 140256 200898 140492 201134
rect 140576 200898 140812 201134
rect 140896 200898 141132 201134
rect 141216 200898 141452 201134
rect 141536 200898 141772 201134
rect 141856 200898 142092 201134
rect 142176 200898 142412 201134
rect 142496 200898 142732 201134
rect 142816 200898 143052 201134
rect 143136 200898 143372 201134
rect 143456 200898 143692 201134
rect 143776 200898 144012 201134
rect 144096 200898 144332 201134
rect 144416 200898 144652 201134
rect 144736 200898 144972 201134
rect 145056 200898 145292 201134
rect 145376 200898 145612 201134
rect 145696 200898 145932 201134
rect 146016 200898 146252 201134
rect 146336 200898 146572 201134
rect 146656 200898 146892 201134
rect 146976 200898 147212 201134
rect 147296 200898 147532 201134
rect 147616 200898 147852 201134
rect 147936 200898 148172 201134
rect 148256 200898 148492 201134
rect 148576 200898 148812 201134
rect 148896 200898 149132 201134
rect 149216 200898 149452 201134
rect 149536 200898 149772 201134
rect 149856 200898 150092 201134
rect 150176 200898 150412 201134
rect 150496 200898 150732 201134
rect 150816 200898 151052 201134
rect 151136 200898 151372 201134
rect 151456 200898 151692 201134
rect 151776 200898 152012 201134
rect 152096 200898 152332 201134
rect 152416 200898 152652 201134
rect 152736 200898 152972 201134
rect 153056 200898 153292 201134
rect 153376 200898 153612 201134
rect 153696 200898 153932 201134
rect 154016 200898 154252 201134
rect 154336 200898 154572 201134
rect 154656 200898 154892 201134
rect 154976 200898 155212 201134
rect 155296 200898 155532 201134
rect 155616 200898 155852 201134
rect 155936 200898 156172 201134
rect 156256 200898 156492 201134
rect 156576 200898 156812 201134
rect 156896 200898 157132 201134
rect 157216 200898 157452 201134
rect 157536 200898 157772 201134
rect 157856 200898 158092 201134
rect 158176 200898 158412 201134
rect 158496 200898 158732 201134
rect 158816 200898 159052 201134
rect 159136 200898 159372 201134
rect 159456 200898 159692 201134
rect 159776 200898 160012 201134
rect 160096 200898 160332 201134
rect 160416 200898 160652 201134
rect 160736 200898 160972 201134
rect 161056 200898 161292 201134
rect 161376 200898 161612 201134
rect 161696 200898 161932 201134
rect 162016 200898 162252 201134
rect 162336 200898 162572 201134
rect 162656 200898 162892 201134
rect 162976 200898 163212 201134
rect 163296 200898 163532 201134
rect 163616 200898 163852 201134
rect 163936 200898 164172 201134
rect 164256 200898 164492 201134
rect 164576 200898 164812 201134
rect 164896 200898 165132 201134
rect 165216 200898 165452 201134
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 139610 115718 139846 115954
rect 139610 115398 139846 115634
rect 170330 115718 170566 115954
rect 170330 115398 170566 115634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 228217 191062 228453
rect 191146 228217 191382 228453
rect 190826 227897 191062 228133
rect 191146 227897 191382 228133
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 228217 227062 228453
rect 227146 228217 227382 228453
rect 226826 227897 227062 228133
rect 227146 227897 227382 228133
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 228217 263062 228453
rect 263146 228217 263382 228453
rect 262826 227897 263062 228133
rect 263146 227897 263382 228133
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 228217 299062 228453
rect 299146 228217 299382 228453
rect 298826 227897 299062 228133
rect 299146 227897 299382 228133
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 228217 335062 228453
rect 335146 228217 335382 228453
rect 334826 227897 335062 228133
rect 335146 227897 335382 228133
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 228217 371062 228453
rect 371146 228217 371382 228453
rect 370826 227897 371062 228133
rect 371146 227897 371382 228133
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246303 424826 246454
rect 29382 246218 65342 246303
rect -8726 246134 65342 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 246067 65342 246134
rect 65578 246067 65662 246303
rect 65898 246067 65982 246303
rect 66218 246067 66302 246303
rect 66538 246067 66622 246303
rect 66858 246067 66942 246303
rect 67178 246067 67262 246303
rect 67498 246067 67582 246303
rect 67818 246067 67902 246303
rect 68138 246067 68222 246303
rect 68458 246067 68542 246303
rect 68778 246067 68862 246303
rect 69098 246067 69182 246303
rect 69418 246067 69502 246303
rect 69738 246067 69822 246303
rect 70058 246218 424826 246303
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect 70058 246134 592650 246218
rect 70058 246067 424826 246134
rect 29382 245898 424826 246067
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241953 420326 241954
rect 24882 241718 65462 241953
rect -8726 241717 65462 241718
rect 65698 241717 65782 241953
rect 66018 241717 66102 241953
rect 66338 241717 66422 241953
rect 66658 241717 66742 241953
rect 66978 241717 67062 241953
rect 67298 241717 67382 241953
rect 67618 241717 67702 241953
rect 67938 241717 68022 241953
rect 68258 241717 68342 241953
rect 68578 241717 68662 241953
rect 68898 241717 68982 241953
rect 69218 241717 69302 241953
rect 69538 241717 69622 241953
rect 69858 241717 69942 241953
rect 70178 241717 70262 241953
rect 70498 241717 70582 241953
rect 70818 241717 70902 241953
rect 71138 241718 420326 241953
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect 71138 241717 592650 241718
rect -8726 241634 592650 241717
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241633 420326 241634
rect 24882 241398 65462 241633
rect -8726 241397 65462 241398
rect 65698 241397 65782 241633
rect 66018 241397 66102 241633
rect 66338 241397 66422 241633
rect 66658 241397 66742 241633
rect 66978 241397 67062 241633
rect 67298 241397 67382 241633
rect 67618 241397 67702 241633
rect 67938 241397 68022 241633
rect 68258 241397 68342 241633
rect 68578 241397 68662 241633
rect 68898 241397 68982 241633
rect 69218 241397 69302 241633
rect 69538 241397 69622 241633
rect 69858 241397 69942 241633
rect 70178 241397 70262 241633
rect 70498 241397 70582 241633
rect 70818 241397 70902 241633
rect 71138 241398 420326 241633
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect 71138 241397 592650 241398
rect -8726 241366 592650 241397
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228453 406826 228454
rect 11382 228218 46826 228453
rect -8726 228217 46826 228218
rect 47062 228217 47146 228453
rect 47382 228217 82826 228453
rect 83062 228217 83146 228453
rect 83382 228217 118826 228453
rect 119062 228217 119146 228453
rect 119382 228217 190826 228453
rect 191062 228217 191146 228453
rect 191382 228217 226826 228453
rect 227062 228217 227146 228453
rect 227382 228217 262826 228453
rect 263062 228217 263146 228453
rect 263382 228217 298826 228453
rect 299062 228217 299146 228453
rect 299382 228217 334826 228453
rect 335062 228217 335146 228453
rect 335382 228217 370826 228453
rect 371062 228217 371146 228453
rect 371382 228218 406826 228453
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect 371382 228217 592650 228218
rect -8726 228134 592650 228217
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 228133 406826 228134
rect 11382 227898 46826 228133
rect -8726 227897 46826 227898
rect 47062 227897 47146 228133
rect 47382 227897 82826 228133
rect 83062 227897 83146 228133
rect 83382 227897 118826 228133
rect 119062 227897 119146 228133
rect 119382 227897 190826 228133
rect 191062 227897 191146 228133
rect 191382 227897 226826 228133
rect 227062 227897 227146 228133
rect 227382 227897 262826 228133
rect 263062 227897 263146 228133
rect 263382 227897 298826 228133
rect 299062 227897 299146 228133
rect 299382 227897 334826 228133
rect 335062 227897 335146 228133
rect 335382 227897 370826 228133
rect 371062 227897 371146 228133
rect 371382 227898 406826 228133
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect 371382 227897 592650 227898
rect -8726 227866 592650 227897
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 136036 205954
rect 136272 205718 136356 205954
rect 136592 205718 136676 205954
rect 136912 205718 136996 205954
rect 137232 205718 137316 205954
rect 137552 205718 137636 205954
rect 137872 205718 137956 205954
rect 138192 205718 138276 205954
rect 138512 205718 138596 205954
rect 138832 205718 138916 205954
rect 139152 205718 139236 205954
rect 139472 205718 139556 205954
rect 139792 205718 139876 205954
rect 140112 205718 140196 205954
rect 140432 205718 140516 205954
rect 140752 205718 140836 205954
rect 141072 205718 141156 205954
rect 141392 205718 141476 205954
rect 141712 205718 141796 205954
rect 142032 205718 142116 205954
rect 142352 205718 142436 205954
rect 142672 205718 142756 205954
rect 142992 205718 143076 205954
rect 143312 205718 143396 205954
rect 143632 205718 143716 205954
rect 143952 205718 144036 205954
rect 144272 205718 144356 205954
rect 144592 205718 144676 205954
rect 144912 205718 144996 205954
rect 145232 205718 145316 205954
rect 145552 205718 145636 205954
rect 145872 205718 145956 205954
rect 146192 205718 146276 205954
rect 146512 205718 146596 205954
rect 146832 205718 146916 205954
rect 147152 205718 147236 205954
rect 147472 205718 147556 205954
rect 147792 205718 147876 205954
rect 148112 205718 148196 205954
rect 148432 205718 148516 205954
rect 148752 205718 148836 205954
rect 149072 205718 149156 205954
rect 149392 205718 149476 205954
rect 149712 205718 149796 205954
rect 150032 205718 150116 205954
rect 150352 205718 150436 205954
rect 150672 205718 150756 205954
rect 150992 205718 151076 205954
rect 151312 205718 151396 205954
rect 151632 205718 151716 205954
rect 151952 205718 152036 205954
rect 152272 205718 152356 205954
rect 152592 205718 152676 205954
rect 152912 205718 152996 205954
rect 153232 205718 153316 205954
rect 153552 205718 153636 205954
rect 153872 205718 153956 205954
rect 154192 205718 154276 205954
rect 154512 205718 154596 205954
rect 154832 205718 154916 205954
rect 155152 205718 155236 205954
rect 155472 205718 155556 205954
rect 155792 205718 155876 205954
rect 156112 205718 156196 205954
rect 156432 205718 156516 205954
rect 156752 205718 156836 205954
rect 157072 205718 157156 205954
rect 157392 205718 157476 205954
rect 157712 205718 157796 205954
rect 158032 205718 158116 205954
rect 158352 205718 158436 205954
rect 158672 205718 158756 205954
rect 158992 205718 159076 205954
rect 159312 205718 159396 205954
rect 159632 205718 159716 205954
rect 159952 205718 160036 205954
rect 160272 205718 160356 205954
rect 160592 205718 160676 205954
rect 160912 205718 160996 205954
rect 161232 205718 161316 205954
rect 161552 205718 161636 205954
rect 161872 205718 161956 205954
rect 162192 205718 162276 205954
rect 162512 205718 162596 205954
rect 162832 205718 162916 205954
rect 163152 205718 163236 205954
rect 163472 205718 163556 205954
rect 163792 205718 163876 205954
rect 164112 205718 164196 205954
rect 164432 205718 164516 205954
rect 164752 205718 164836 205954
rect 165072 205718 165156 205954
rect 165392 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 136036 205634
rect 136272 205398 136356 205634
rect 136592 205398 136676 205634
rect 136912 205398 136996 205634
rect 137232 205398 137316 205634
rect 137552 205398 137636 205634
rect 137872 205398 137956 205634
rect 138192 205398 138276 205634
rect 138512 205398 138596 205634
rect 138832 205398 138916 205634
rect 139152 205398 139236 205634
rect 139472 205398 139556 205634
rect 139792 205398 139876 205634
rect 140112 205398 140196 205634
rect 140432 205398 140516 205634
rect 140752 205398 140836 205634
rect 141072 205398 141156 205634
rect 141392 205398 141476 205634
rect 141712 205398 141796 205634
rect 142032 205398 142116 205634
rect 142352 205398 142436 205634
rect 142672 205398 142756 205634
rect 142992 205398 143076 205634
rect 143312 205398 143396 205634
rect 143632 205398 143716 205634
rect 143952 205398 144036 205634
rect 144272 205398 144356 205634
rect 144592 205398 144676 205634
rect 144912 205398 144996 205634
rect 145232 205398 145316 205634
rect 145552 205398 145636 205634
rect 145872 205398 145956 205634
rect 146192 205398 146276 205634
rect 146512 205398 146596 205634
rect 146832 205398 146916 205634
rect 147152 205398 147236 205634
rect 147472 205398 147556 205634
rect 147792 205398 147876 205634
rect 148112 205398 148196 205634
rect 148432 205398 148516 205634
rect 148752 205398 148836 205634
rect 149072 205398 149156 205634
rect 149392 205398 149476 205634
rect 149712 205398 149796 205634
rect 150032 205398 150116 205634
rect 150352 205398 150436 205634
rect 150672 205398 150756 205634
rect 150992 205398 151076 205634
rect 151312 205398 151396 205634
rect 151632 205398 151716 205634
rect 151952 205398 152036 205634
rect 152272 205398 152356 205634
rect 152592 205398 152676 205634
rect 152912 205398 152996 205634
rect 153232 205398 153316 205634
rect 153552 205398 153636 205634
rect 153872 205398 153956 205634
rect 154192 205398 154276 205634
rect 154512 205398 154596 205634
rect 154832 205398 154916 205634
rect 155152 205398 155236 205634
rect 155472 205398 155556 205634
rect 155792 205398 155876 205634
rect 156112 205398 156196 205634
rect 156432 205398 156516 205634
rect 156752 205398 156836 205634
rect 157072 205398 157156 205634
rect 157392 205398 157476 205634
rect 157712 205398 157796 205634
rect 158032 205398 158116 205634
rect 158352 205398 158436 205634
rect 158672 205398 158756 205634
rect 158992 205398 159076 205634
rect 159312 205398 159396 205634
rect 159632 205398 159716 205634
rect 159952 205398 160036 205634
rect 160272 205398 160356 205634
rect 160592 205398 160676 205634
rect 160912 205398 160996 205634
rect 161232 205398 161316 205634
rect 161552 205398 161636 205634
rect 161872 205398 161956 205634
rect 162192 205398 162276 205634
rect 162512 205398 162596 205634
rect 162832 205398 162916 205634
rect 163152 205398 163236 205634
rect 163472 205398 163556 205634
rect 163792 205398 163876 205634
rect 164112 205398 164196 205634
rect 164432 205398 164516 205634
rect 164752 205398 164836 205634
rect 165072 205398 165156 205634
rect 165392 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 137376 201454
rect 137612 201218 137696 201454
rect 137932 201218 138016 201454
rect 138252 201218 138336 201454
rect 138572 201218 138656 201454
rect 138892 201218 138976 201454
rect 139212 201218 139296 201454
rect 139532 201218 139616 201454
rect 139852 201218 139936 201454
rect 140172 201218 140256 201454
rect 140492 201218 140576 201454
rect 140812 201218 140896 201454
rect 141132 201218 141216 201454
rect 141452 201218 141536 201454
rect 141772 201218 141856 201454
rect 142092 201218 142176 201454
rect 142412 201218 142496 201454
rect 142732 201218 142816 201454
rect 143052 201218 143136 201454
rect 143372 201218 143456 201454
rect 143692 201218 143776 201454
rect 144012 201218 144096 201454
rect 144332 201218 144416 201454
rect 144652 201218 144736 201454
rect 144972 201218 145056 201454
rect 145292 201218 145376 201454
rect 145612 201218 145696 201454
rect 145932 201218 146016 201454
rect 146252 201218 146336 201454
rect 146572 201218 146656 201454
rect 146892 201218 146976 201454
rect 147212 201218 147296 201454
rect 147532 201218 147616 201454
rect 147852 201218 147936 201454
rect 148172 201218 148256 201454
rect 148492 201218 148576 201454
rect 148812 201218 148896 201454
rect 149132 201218 149216 201454
rect 149452 201218 149536 201454
rect 149772 201218 149856 201454
rect 150092 201218 150176 201454
rect 150412 201218 150496 201454
rect 150732 201218 150816 201454
rect 151052 201218 151136 201454
rect 151372 201218 151456 201454
rect 151692 201218 151776 201454
rect 152012 201218 152096 201454
rect 152332 201218 152416 201454
rect 152652 201218 152736 201454
rect 152972 201218 153056 201454
rect 153292 201218 153376 201454
rect 153612 201218 153696 201454
rect 153932 201218 154016 201454
rect 154252 201218 154336 201454
rect 154572 201218 154656 201454
rect 154892 201218 154976 201454
rect 155212 201218 155296 201454
rect 155532 201218 155616 201454
rect 155852 201218 155936 201454
rect 156172 201218 156256 201454
rect 156492 201218 156576 201454
rect 156812 201218 156896 201454
rect 157132 201218 157216 201454
rect 157452 201218 157536 201454
rect 157772 201218 157856 201454
rect 158092 201218 158176 201454
rect 158412 201218 158496 201454
rect 158732 201218 158816 201454
rect 159052 201218 159136 201454
rect 159372 201218 159456 201454
rect 159692 201218 159776 201454
rect 160012 201218 160096 201454
rect 160332 201218 160416 201454
rect 160652 201218 160736 201454
rect 160972 201218 161056 201454
rect 161292 201218 161376 201454
rect 161612 201218 161696 201454
rect 161932 201218 162016 201454
rect 162252 201218 162336 201454
rect 162572 201218 162656 201454
rect 162892 201218 162976 201454
rect 163212 201218 163296 201454
rect 163532 201218 163616 201454
rect 163852 201218 163936 201454
rect 164172 201218 164256 201454
rect 164492 201218 164576 201454
rect 164812 201218 164896 201454
rect 165132 201218 165216 201454
rect 165452 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 137376 201134
rect 137612 200898 137696 201134
rect 137932 200898 138016 201134
rect 138252 200898 138336 201134
rect 138572 200898 138656 201134
rect 138892 200898 138976 201134
rect 139212 200898 139296 201134
rect 139532 200898 139616 201134
rect 139852 200898 139936 201134
rect 140172 200898 140256 201134
rect 140492 200898 140576 201134
rect 140812 200898 140896 201134
rect 141132 200898 141216 201134
rect 141452 200898 141536 201134
rect 141772 200898 141856 201134
rect 142092 200898 142176 201134
rect 142412 200898 142496 201134
rect 142732 200898 142816 201134
rect 143052 200898 143136 201134
rect 143372 200898 143456 201134
rect 143692 200898 143776 201134
rect 144012 200898 144096 201134
rect 144332 200898 144416 201134
rect 144652 200898 144736 201134
rect 144972 200898 145056 201134
rect 145292 200898 145376 201134
rect 145612 200898 145696 201134
rect 145932 200898 146016 201134
rect 146252 200898 146336 201134
rect 146572 200898 146656 201134
rect 146892 200898 146976 201134
rect 147212 200898 147296 201134
rect 147532 200898 147616 201134
rect 147852 200898 147936 201134
rect 148172 200898 148256 201134
rect 148492 200898 148576 201134
rect 148812 200898 148896 201134
rect 149132 200898 149216 201134
rect 149452 200898 149536 201134
rect 149772 200898 149856 201134
rect 150092 200898 150176 201134
rect 150412 200898 150496 201134
rect 150732 200898 150816 201134
rect 151052 200898 151136 201134
rect 151372 200898 151456 201134
rect 151692 200898 151776 201134
rect 152012 200898 152096 201134
rect 152332 200898 152416 201134
rect 152652 200898 152736 201134
rect 152972 200898 153056 201134
rect 153292 200898 153376 201134
rect 153612 200898 153696 201134
rect 153932 200898 154016 201134
rect 154252 200898 154336 201134
rect 154572 200898 154656 201134
rect 154892 200898 154976 201134
rect 155212 200898 155296 201134
rect 155532 200898 155616 201134
rect 155852 200898 155936 201134
rect 156172 200898 156256 201134
rect 156492 200898 156576 201134
rect 156812 200898 156896 201134
rect 157132 200898 157216 201134
rect 157452 200898 157536 201134
rect 157772 200898 157856 201134
rect 158092 200898 158176 201134
rect 158412 200898 158496 201134
rect 158732 200898 158816 201134
rect 159052 200898 159136 201134
rect 159372 200898 159456 201134
rect 159692 200898 159776 201134
rect 160012 200898 160096 201134
rect 160332 200898 160416 201134
rect 160652 200898 160736 201134
rect 160972 200898 161056 201134
rect 161292 200898 161376 201134
rect 161612 200898 161696 201134
rect 161932 200898 162016 201134
rect 162252 200898 162336 201134
rect 162572 200898 162656 201134
rect 162892 200898 162976 201134
rect 163212 200898 163296 201134
rect 163532 200898 163616 201134
rect 163852 200898 163936 201134
rect 164172 200898 164256 201134
rect 164492 200898 164576 201134
rect 164812 200898 164896 201134
rect 165132 200898 165216 201134
rect 165452 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 139610 115954
rect 139846 115718 170330 115954
rect 170566 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 139610 115634
rect 139846 115398 170330 115634
rect 170566 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 154970 111454
rect 155206 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 154970 111134
rect 155206 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use PD_M1_M2  PD_M1_M2_macro0
timestamp 0
transform 1 0 16000 0 1 232484
box 30000 -2000 380500 14200
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 120000 0 1 80000
box 0 0 60000 60000
use SystemLevel  sl_macro0
timestamp 0
transform 1 0 148914 0 1 188066
box -13000 -14480 17120 18000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 248684 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 248684 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 248684 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 142000 182414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 248684 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 248684 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 248684 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 248684 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 248684 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 248684 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 248684 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 248684 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 248684 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 142000 119414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 248684 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 248684 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 248684 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 248684 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 248684 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 248684 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 248684 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 248684 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 248684 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 248684 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 142000 128414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 248684 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 248684 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 248684 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 248684 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 248684 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 248684 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 248684 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 248684 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 248684 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 248684 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 248684 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 142000 173414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 248684 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 248684 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 248684 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 248684 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 248684 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 248684 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 248684 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 248684 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 248684 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 142000 132914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 248684 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 142000 168914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 248684 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 248684 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 248684 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 248684 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 248684 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 248684 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 248684 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 248684 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 248684 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 248684 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 142000 177914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 248684 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 248684 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 248684 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 248684 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 248684 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 248684 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 248684 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 248684 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 248684 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 248684 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 248684 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 248684 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 248684 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 248684 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 248684 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 248684 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 248684 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 248684 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 142000 123914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 248684 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 248684 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 248684 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 248684 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 248684 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 248684 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 248684 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 248684 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
