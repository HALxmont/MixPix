* NGSPICE file created from pixel_macro.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_2 abstract view
.subckt sky130_fd_sc_hd__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

.subckt pixel_macro io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2]
+ io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103]
+ la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108]
+ la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113]
+ la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118]
+ la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123]
+ la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35]
+ la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40]
+ la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
+ la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51]
+ la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57]
+ la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62]
+ la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68]
+ la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73]
+ la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79]
+ la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84]
+ la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8]
+ la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95]
+ la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0]
+ la_data_out[100] la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104]
+ la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109]
+ la_data_out[10] la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113]
+ la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118]
+ la_data_out[119] la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61]
+ la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66]
+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71]
+ la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
+ la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100]
+ la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107]
+ la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113]
+ la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11]
+ la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126]
+ la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
+ la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
+ la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2]
+ la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36]
+ la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42]
+ la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49]
+ la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55]
+ la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61]
+ la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68]
+ la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74]
+ la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80]
+ la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87]
+ la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93]
+ la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9]
+ vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0422__B _0820_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0613__A _1141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output56_A _0829_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater71 _0442_/X vssd1 vssd1 vccd1 vccd1 repeater71/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater82 repeater83/X vssd1 vssd1 vccd1 vccd1 repeater82/X sky130_fd_sc_hd__clkbuf_2
X_0419_ _0823_/Q _0433_/B vssd1 vssd1 vccd1 vccd1 _0503_/B sky130_fd_sc_hd__nand2b_2
XFILLER_27_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0417__B _0438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xpixel_macro_283 vssd1 vssd1 vccd1 vccd1 pixel_macro_283/HI wbs_dat_o[19] sky130_fd_sc_hd__conb_1
Xpixel_macro_272 vssd1 vssd1 vccd1 vccd1 pixel_macro_272/HI la_data_out[121] sky130_fd_sc_hd__conb_1
Xpixel_macro_250 vssd1 vssd1 vccd1 vccd1 pixel_macro_250/HI la_data_out[99] sky130_fd_sc_hd__conb_1
Xpixel_macro_261 vssd1 vssd1 vccd1 vccd1 pixel_macro_261/HI la_data_out[110] sky130_fd_sc_hd__conb_1
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xpixel_macro_294 vssd1 vssd1 vccd1 vccd1 pixel_macro_294/HI wbs_dat_o[30] sky130_fd_sc_hd__conb_1
XFILLER_7_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0770_ _0794_/B vssd1 vssd1 vccd1 vccd1 _0780_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0899_ _0899_/D _0436_/Y vssd1 vssd1 vccd1 vccd1 _0899_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_23_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0822_ _0921_/CLK _0822_/D _0751_/Y vssd1 vssd1 vccd1 vccd1 _0822_/Q sky130_fd_sc_hd__dfrtp_1
X_0753_ input1/X _0754_/B vssd1 vssd1 vccd1 vccd1 _0824_/D sky130_fd_sc_hd__nor2_1
X_0684_ _0684_/A _0684_/B vssd1 vssd1 vccd1 vccd1 _0686_/C sky130_fd_sc_hd__and2_1
XFILLER_6_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_515 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0832__CLK _0838_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0805_ _0829_/CLK _0805_/D vssd1 vssd1 vccd1 vccd1 _0805_/Q sky130_fd_sc_hd__dfxtp_1
X_0667_ _0667_/A vssd1 vssd1 vccd1 vccd1 _0917_/D sky130_fd_sc_hd__clkbuf_1
X_0598_ _0598_/A vssd1 vssd1 vccd1 vccd1 _0881_/D sky130_fd_sc_hd__clkbuf_1
X_0736_ _0736_/A vssd1 vssd1 vccd1 vccd1 _0736_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0706__A _0706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0762__A1 _0756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0616__A _0622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input18_A wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0452_ _0452_/A vssd1 vssd1 vccd1 vccd1 _0452_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0521_ _0666_/B vssd1 vssd1 vccd1 vccd1 _0627_/B sky130_fd_sc_hd__clkbuf_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0719_ _0754_/A input6/X _0719_/C vssd1 vssd1 vccd1 vccd1 _0737_/A sky130_fd_sc_hd__nor3_2
XFILLER_15_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput42 _0433_/B vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
Xoutput31 _1140_/A vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
Xoutput53 _0826_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
XFILLER_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0504_ _0659_/B vssd1 vssd1 vccd1 vccd1 _0649_/B sky130_fd_sc_hd__clkbuf_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0435_ _0560_/B _0756_/C vssd1 vssd1 vccd1 vccd1 _0435_/Y sky130_fd_sc_hd__nor2_1
XTAP_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0414__B1 _0918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0717__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0708__A1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater83 _0477_/X vssd1 vssd1 vccd1 vccd1 repeater83/X sky130_fd_sc_hd__clkbuf_1
Xrepeater72 _0436_/Y vssd1 vssd1 vccd1 vccd1 _0444_/A sky130_fd_sc_hd__clkbuf_1
X_0418_ _0438_/A vssd1 vssd1 vccd1 vccd1 _0451_/A sky130_fd_sc_hd__inv_2
XFILLER_27_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_284 vssd1 vssd1 vccd1 vccd1 pixel_macro_284/HI wbs_dat_o[20] sky130_fd_sc_hd__conb_1
Xpixel_macro_273 vssd1 vssd1 vccd1 vccd1 pixel_macro_273/HI la_data_out[122] sky130_fd_sc_hd__conb_1
Xpixel_macro_262 vssd1 vssd1 vccd1 vccd1 pixel_macro_262/HI la_data_out[111] sky130_fd_sc_hd__conb_1
Xpixel_macro_240 vssd1 vssd1 vccd1 vccd1 pixel_macro_240/HI la_data_out[89] sky130_fd_sc_hd__conb_1
Xpixel_macro_251 vssd1 vssd1 vccd1 vccd1 pixel_macro_251/HI la_data_out[100] sky130_fd_sc_hd__conb_1
Xpixel_macro_295 vssd1 vssd1 vccd1 vccd1 pixel_macro_295/HI wbs_dat_o[31] sky130_fd_sc_hd__conb_1
XANTENNA__0714__A _0731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0433__B _0433_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0534__A _0538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0898_ _0898_/D _0442_/X vssd1 vssd1 vccd1 vccd1 _0910_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA__0428__B _0655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0752_ _0797_/A vssd1 vssd1 vccd1 vccd1 _0752_/Y sky130_fd_sc_hd__inv_2
X_0821_ _0921_/CLK _0821_/D _0750_/Y vssd1 vssd1 vccd1 vccd1 _0821_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_9_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0683_ input9/X _0754_/C vssd1 vssd1 vccd1 vccd1 _0705_/A sky130_fd_sc_hd__nor2_2
XFILLER_6_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0529__A _0551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_232 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output31_A _1140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0735_ _0735_/A vssd1 vssd1 vccd1 vccd1 _0735_/X sky130_fd_sc_hd__clkbuf_2
X_0804_ _0829_/CLK _0804_/D vssd1 vssd1 vccd1 vccd1 _0804_/Q sky130_fd_sc_hd__dfxtp_1
X_0597_ _0605_/A _0649_/B vssd1 vssd1 vccd1 vccd1 _0598_/A sky130_fd_sc_hd__and2_1
X_0666_ _0756_/B _0666_/B vssd1 vssd1 vccd1 vccd1 _0667_/A sky130_fd_sc_hd__and2_1
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_335 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0632__A _0640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0520_ _0520_/A vssd1 vssd1 vccd1 vccd1 _0850_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0451_ _0451_/A _0666_/B vssd1 vssd1 vccd1 vccd1 _0452_/A sky130_fd_sc_hd__or2_1
XANTENNA__0729__C1 _0714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0718_ input9/X vssd1 vssd1 vccd1 vccd1 _0754_/A sky130_fd_sc_hd__inv_2
X_0649_ _0649_/A _0649_/B vssd1 vssd1 vccd1 vccd1 _0650_/A sky130_fd_sc_hd__and2_1
XFILLER_15_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0822__CLK _0921_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput43 _0823_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
Xoutput32 _1141_/A vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput54 _0827_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
XANTENNA__0627__A _0649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0434_ _0434_/A _0510_/B vssd1 vssd1 vccd1 vccd1 _0756_/C sky130_fd_sc_hd__nor2_2
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0503_ _0510_/A _0503_/B vssd1 vssd1 vccd1 vccd1 _0659_/B sky130_fd_sc_hd__nor2_1
XANTENNA__0414__A1 _0756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_190 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater62 _0450_/X vssd1 vssd1 vccd1 vccd1 repeater62/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater73 _0931_/Q vssd1 vssd1 vccd1 vccd1 _0551_/A sky130_fd_sc_hd__clkbuf_2
Xrepeater84 _0477_/X vssd1 vssd1 vccd1 vccd1 repeater84/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0417_ _0756_/A _0438_/A vssd1 vssd1 vccd1 vccd1 _0417_/Y sky130_fd_sc_hd__nor2_1
Xpixel_macro_285 vssd1 vssd1 vccd1 vccd1 pixel_macro_285/HI wbs_dat_o[21] sky130_fd_sc_hd__conb_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xpixel_macro_252 vssd1 vssd1 vccd1 vccd1 pixel_macro_252/HI la_data_out[101] sky130_fd_sc_hd__conb_1
Xpixel_macro_230 vssd1 vssd1 vccd1 vccd1 pixel_macro_230/HI la_data_out[79] sky130_fd_sc_hd__conb_1
Xpixel_macro_263 vssd1 vssd1 vccd1 vccd1 pixel_macro_263/HI la_data_out[112] sky130_fd_sc_hd__conb_1
Xpixel_macro_241 vssd1 vssd1 vccd1 vccd1 pixel_macro_241/HI la_data_out[90] sky130_fd_sc_hd__conb_1
Xpixel_macro_274 vssd1 vssd1 vccd1 vccd1 pixel_macro_274/HI la_data_out[123] sky130_fd_sc_hd__conb_1
XFILLER_10_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0640__A _0640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0897_ _0897_/D _0435_/Y vssd1 vssd1 vccd1 vccd1 _0897_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_4_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0820_ _0921_/CLK _0820_/D _0680_/X vssd1 vssd1 vccd1 vccd1 _0820_/Q sky130_fd_sc_hd__dfstp_1
X_0751_ _0797_/A vssd1 vssd1 vccd1 vccd1 _0751_/Y sky130_fd_sc_hd__inv_2
X_0682_ input3/X input2/X input6/X vssd1 vssd1 vccd1 vccd1 _0754_/C sky130_fd_sc_hd__or3b_1
XFILLER_25_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0545__A _0549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0665_ _0665_/A vssd1 vssd1 vccd1 vccd1 _0903_/D sky130_fd_sc_hd__clkbuf_1
X_0734_ input19/X _0721_/X _0733_/X _0731_/X vssd1 vssd1 vccd1 vccd1 _0814_/D sky130_fd_sc_hd__o211a_1
X_0803_ _0829_/CLK _0803_/D vssd1 vssd1 vccd1 vccd1 _0803_/Q sky130_fd_sc_hd__dfxtp_1
X_0596_ _0609_/A vssd1 vssd1 vccd1 vccd1 _0605_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_347 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0450_ _0450_/A vssd1 vssd1 vccd1 vccd1 _0450_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0648_ _0648_/A vssd1 vssd1 vccd1 vccd1 _0912_/D sky130_fd_sc_hd__clkbuf_1
X_0717_ input24/X _0704_/X _0716_/X _0714_/X vssd1 vssd1 vccd1 vccd1 _0809_/D sky130_fd_sc_hd__o211a_1
XFILLER_26_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0579_ _0579_/A _0627_/B vssd1 vssd1 vccd1 vccd1 _0580_/A sky130_fd_sc_hd__and2_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput44 _1138_/X vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
Xoutput33 _0609_/A vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
Xoutput55 _0828_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XANTENNA_input23_A wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0643__A _0661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0408__C1 _0918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0502_ _0525_/A vssd1 vssd1 vccd1 vccd1 _0519_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0433_ _0433_/A _0433_/B vssd1 vssd1 vccd1 vccd1 _0510_/B sky130_fd_sc_hd__or2_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0414__A2 _0925_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0638__A _0640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_431 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater63 _0448_/X vssd1 vssd1 vccd1 vccd1 repeater63/X sky130_fd_sc_hd__clkbuf_1
Xrepeater85 _0439_/B vssd1 vssd1 vccd1 vccd1 repeater85/X sky130_fd_sc_hd__clkbuf_1
Xrepeater74 _0930_/Q vssd1 vssd1 vccd1 vccd1 _0525_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_242 vssd1 vssd1 vccd1 vccd1 pixel_macro_242/HI la_data_out[91] sky130_fd_sc_hd__conb_1
Xpixel_macro_231 vssd1 vssd1 vccd1 vccd1 pixel_macro_231/HI la_data_out[80] sky130_fd_sc_hd__conb_1
Xpixel_macro_220 vssd1 vssd1 vccd1 vccd1 pixel_macro_220/HI la_data_out[69] sky130_fd_sc_hd__conb_1
X_0416_ _0823_/Q _0822_/Q _0821_/Q vssd1 vssd1 vccd1 vccd1 _0438_/A sky130_fd_sc_hd__or3b_2
XANTENNA__0812__CLK _0838_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xpixel_macro_264 vssd1 vssd1 vccd1 vccd1 pixel_macro_264/HI la_data_out[113] sky130_fd_sc_hd__conb_1
Xpixel_macro_253 vssd1 vssd1 vccd1 vccd1 pixel_macro_253/HI la_data_out[102] sky130_fd_sc_hd__conb_1
Xpixel_macro_275 vssd1 vssd1 vccd1 vccd1 pixel_macro_275/HI la_data_out[124] sky130_fd_sc_hd__conb_1
Xpixel_macro_286 vssd1 vssd1 vccd1 vccd1 pixel_macro_286/HI wbs_dat_o[22] sky130_fd_sc_hd__conb_1
XFILLER_12_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0835__CLK _0838_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0896_ _0896_/D _0429_/X vssd1 vssd1 vccd1 vccd1 _0908_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_11_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0681_ _0799_/Q _0677_/Y _0678_/X _0680_/X vssd1 vssd1 vccd1 vccd1 _0799_/D sky130_fd_sc_hd__o211a_1
X_0750_ _0797_/A vssd1 vssd1 vccd1 vccd1 _0750_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0774__A1 _0913_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0879_ _0879_/D _0762_/A2 vssd1 vssd1 vccd1 vccd1 _0916_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_18_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0802_ _0829_/CLK _0802_/D vssd1 vssd1 vccd1 vccd1 _0802_/Q sky130_fd_sc_hd__dfxtp_1
X_0733_ _0722_/X _0723_/X _0814_/Q vssd1 vssd1 vccd1 vccd1 _0733_/X sky130_fd_sc_hd__a21o_1
X_0664_ _0756_/B _0664_/B vssd1 vssd1 vccd1 vccd1 _0665_/A sky130_fd_sc_hd__and2_1
X_0595_ _0595_/A vssd1 vssd1 vccd1 vccd1 _0887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0729__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0647_ _0649_/A _0647_/B vssd1 vssd1 vccd1 vccd1 _0648_/A sky130_fd_sc_hd__and2_1
X_0716_ _0705_/X _0706_/X _0809_/Q vssd1 vssd1 vccd1 vccd1 _0716_/X sky130_fd_sc_hd__a21o_1
XFILLER_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0578_ _0578_/A vssd1 vssd1 vccd1 vccd1 _0876_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0919__CLK _0921_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput34 _0579_/A vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
Xoutput45 _1139_/X vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
Xoutput56 _0829_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
XANTENNA_input16_A wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0501_ _0501_/A vssd1 vssd1 vccd1 vccd1 _0848_/D sky130_fd_sc_hd__clkbuf_1
X_0432_ _0668_/B vssd1 vssd1 vccd1 vccd1 _0918_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input8_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater64 _0429_/X vssd1 vssd1 vccd1 vccd1 repeater64/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater75 _0655_/A vssd1 vssd1 vccd1 vccd1 _1141_/A sky130_fd_sc_hd__clkbuf_1
Xrepeater86 _0441_/A vssd1 vssd1 vccd1 vccd1 _0439_/B sky130_fd_sc_hd__clkbuf_1
X_0415_ _0756_/A _0406_/C _0414_/Y vssd1 vssd1 vccd1 vccd1 _0820_/D sky130_fd_sc_hd__o21a_1
XFILLER_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xpixel_macro_243 vssd1 vssd1 vccd1 vccd1 pixel_macro_243/HI la_data_out[92] sky130_fd_sc_hd__conb_1
Xpixel_macro_232 vssd1 vssd1 vccd1 vccd1 pixel_macro_232/HI la_data_out[81] sky130_fd_sc_hd__conb_1
Xpixel_macro_221 vssd1 vssd1 vccd1 vccd1 pixel_macro_221/HI la_data_out[70] sky130_fd_sc_hd__conb_1
Xpixel_macro_210 vssd1 vssd1 vccd1 vccd1 pixel_macro_210/HI la_data_out[59] sky130_fd_sc_hd__conb_1
Xpixel_macro_265 vssd1 vssd1 vccd1 vccd1 pixel_macro_265/HI la_data_out[114] sky130_fd_sc_hd__conb_1
Xpixel_macro_254 vssd1 vssd1 vccd1 vccd1 pixel_macro_254/HI la_data_out[103] sky130_fd_sc_hd__conb_1
XANTENNA__0564__A _0566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xpixel_macro_287 vssd1 vssd1 vccd1 vccd1 pixel_macro_287/HI wbs_dat_o[23] sky130_fd_sc_hd__conb_1
XFILLER_11_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xpixel_macro_276 vssd1 vssd1 vccd1 vccd1 pixel_macro_276/HI la_data_out[125] sky130_fd_sc_hd__conb_1
XFILLER_10_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0795__C1 _0731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0649__A _0649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0895_ _0895_/D repeater62/X vssd1 vssd1 vccd1 vccd1 _0907_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA__0710__C1 _0700_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0701__C1 _0700_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0680_ _0781_/A vssd1 vssd1 vccd1 vccd1 _0680_/X sky130_fd_sc_hd__buf_2
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0802__CLK _0829_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0878_ _0878_/D repeater63/X vssd1 vssd1 vccd1 vccd1 _0915_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_18_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0825__CLK _0838_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0801_ _0838_/CLK _0801_/D vssd1 vssd1 vccd1 vccd1 _0801_/Q sky130_fd_sc_hd__dfxtp_1
X_0594_ _0594_/A _0647_/B vssd1 vssd1 vccd1 vccd1 _0595_/A sky130_fd_sc_hd__and2_1
X_0732_ input18/X _0721_/X _0730_/X _0731_/X vssd1 vssd1 vccd1 vccd1 _0813_/D sky130_fd_sc_hd__o211a_1
XFILLER_6_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0663_ _0927_/Q vssd1 vssd1 vccd1 vccd1 _0756_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_25_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0657__A _0661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0715_ input23/X _0704_/X _0713_/X _0714_/X vssd1 vssd1 vccd1 vccd1 _0808_/D sky130_fd_sc_hd__o211a_1
X_0577_ _0577_/A _0625_/B vssd1 vssd1 vccd1 vccd1 _0578_/A sky130_fd_sc_hd__and2_1
X_0646_ _0646_/A vssd1 vssd1 vccd1 vccd1 _0902_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput35 _0525_/A vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput46 _0824_/Q vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
XFILLER_5_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput57 _0830_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XFILLER_16_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0500_ _0500_/A _0647_/B vssd1 vssd1 vccd1 vccd1 _0501_/A sky130_fd_sc_hd__and2_1
X_0431_ _0486_/B _0495_/B vssd1 vssd1 vccd1 vccd1 _0668_/B sky130_fd_sc_hd__nor2_2
XTAP_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0629_ _0649_/A _0668_/B vssd1 vssd1 vccd1 vccd1 _0630_/A sky130_fd_sc_hd__and2_1
XFILLER_26_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater65 _0445_/X vssd1 vssd1 vccd1 vccd1 repeater65/X sky130_fd_sc_hd__clkbuf_1
Xrepeater87 repeater88/X vssd1 vssd1 vccd1 vccd1 repeater87/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater76 _0929_/Q vssd1 vssd1 vccd1 vccd1 _0655_/A sky130_fd_sc_hd__clkbuf_1
X_0414_ _0756_/A _0925_/Q _0918_/Q vssd1 vssd1 vccd1 vccd1 _0414_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xpixel_macro_288 vssd1 vssd1 vccd1 vccd1 pixel_macro_288/HI wbs_dat_o[24] sky130_fd_sc_hd__conb_1
Xpixel_macro_266 vssd1 vssd1 vccd1 vccd1 pixel_macro_266/HI la_data_out[115] sky130_fd_sc_hd__conb_1
Xpixel_macro_255 vssd1 vssd1 vccd1 vccd1 pixel_macro_255/HI la_data_out[104] sky130_fd_sc_hd__conb_1
Xpixel_macro_244 vssd1 vssd1 vccd1 vccd1 pixel_macro_244/HI la_data_out[93] sky130_fd_sc_hd__conb_1
Xpixel_macro_233 vssd1 vssd1 vccd1 vccd1 pixel_macro_233/HI la_data_out[82] sky130_fd_sc_hd__conb_1
Xpixel_macro_222 vssd1 vssd1 vccd1 vccd1 pixel_macro_222/HI la_data_out[71] sky130_fd_sc_hd__conb_1
Xpixel_macro_211 vssd1 vssd1 vccd1 vccd1 pixel_macro_211/HI la_data_out[60] sky130_fd_sc_hd__conb_1
Xpixel_macro_200 vssd1 vssd1 vccd1 vccd1 pixel_macro_200/HI la_data_out[49] sky130_fd_sc_hd__conb_1
Xpixel_macro_277 vssd1 vssd1 vccd1 vccd1 pixel_macro_277/HI la_data_out[126] sky130_fd_sc_hd__conb_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0490__A _0500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0894_ _0894_/D repeater65/X vssd1 vssd1 vccd1 vccd1 _0904_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_9_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0575__A _0577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0485__A _0525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0877_ _0877_/D repeater65/X vssd1 vssd1 vccd1 vccd1 _0904_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_0_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0695__C1 _0680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_520 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0731_ _0731_/A vssd1 vssd1 vccd1 vccd1 _0731_/X sky130_fd_sc_hd__clkbuf_2
X_0800_ _0838_/CLK _0800_/D vssd1 vssd1 vccd1 vccd1 _0800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0593_ _0593_/A vssd1 vssd1 vccd1 vccd1 _0880_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0662_ _0662_/A vssd1 vssd1 vccd1 vccd1 _0898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0929_ _0929_/D repeater82/X vssd1 vssd1 vccd1 vccd1 _0929_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_0_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0714_ _0731_/A vssd1 vssd1 vccd1 vccd1 _0714_/X sky130_fd_sc_hd__clkbuf_2
X_0645_ _0661_/A _0645_/B vssd1 vssd1 vccd1 vccd1 _0646_/A sky130_fd_sc_hd__and2_1
X_0576_ _0576_/A vssd1 vssd1 vccd1 vccd1 _0871_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0815__CLK _0829_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput36 _0551_/A vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
Xoutput58 _0831_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
Xoutput47 _0825_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0493__A _0500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0408__A2 _0560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0668__A _0756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0430_ _0433_/B _0433_/A vssd1 vssd1 vccd1 vccd1 _0495_/B sky130_fd_sc_hd__nand2b_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0838__CLK _0838_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0628_ _0628_/A vssd1 vssd1 vccd1 vccd1 _0909_/D sky130_fd_sc_hd__clkbuf_1
X_0559_ _0559_/A vssd1 vssd1 vccd1 vccd1 _0877_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0488__A _0500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input21_A wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater66 _0449_/B vssd1 vssd1 vccd1 vccd1 repeater66/X sky130_fd_sc_hd__clkbuf_1
Xrepeater77 _0928_/Q vssd1 vssd1 vccd1 vccd1 _0609_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater88 _0451_/A vssd1 vssd1 vccd1 vccd1 repeater88/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0398__A _0823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0413_ _0918_/Q _0413_/B _0413_/C vssd1 vssd1 vccd1 vccd1 _0821_/D sky130_fd_sc_hd__nor3_1
Xpixel_macro_289 vssd1 vssd1 vccd1 vccd1 pixel_macro_289/HI wbs_dat_o[25] sky130_fd_sc_hd__conb_1
Xpixel_macro_278 vssd1 vssd1 vccd1 vccd1 pixel_macro_278/HI la_data_out[127] sky130_fd_sc_hd__conb_1
Xpixel_macro_267 vssd1 vssd1 vccd1 vccd1 pixel_macro_267/HI la_data_out[116] sky130_fd_sc_hd__conb_1
Xpixel_macro_256 vssd1 vssd1 vccd1 vccd1 pixel_macro_256/HI la_data_out[105] sky130_fd_sc_hd__conb_1
Xpixel_macro_223 vssd1 vssd1 vccd1 vccd1 pixel_macro_223/HI la_data_out[72] sky130_fd_sc_hd__conb_1
Xpixel_macro_201 vssd1 vssd1 vccd1 vccd1 pixel_macro_201/HI la_data_out[50] sky130_fd_sc_hd__conb_1
Xpixel_macro_212 vssd1 vssd1 vccd1 vccd1 pixel_macro_212/HI la_data_out[61] sky130_fd_sc_hd__conb_1
Xpixel_macro_245 vssd1 vssd1 vccd1 vccd1 pixel_macro_245/HI la_data_out[94] sky130_fd_sc_hd__conb_1
Xpixel_macro_234 vssd1 vssd1 vccd1 vccd1 pixel_macro_234/HI la_data_out[83] sky130_fd_sc_hd__conb_1
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_220 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0490__B _0560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0771__A _0829_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0893_ _0893_/D _0436_/Y vssd1 vssd1 vccd1 vccd1 _0899_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_9_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0575__B _0653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0710__A1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0701__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0876_ _0876_/D repeater85/X vssd1 vssd1 vccd1 vccd1 _0914_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_18_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_532 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0730_ _0722_/X _0723_/X _0813_/Q vssd1 vssd1 vccd1 vccd1 _0730_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0661_ _0661_/A _0661_/B vssd1 vssd1 vccd1 vccd1 _0662_/A sky130_fd_sc_hd__and2_1
XFILLER_27_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0592_ _0594_/A _0620_/B vssd1 vssd1 vccd1 vccd1 _0593_/A sky130_fd_sc_hd__and2_1
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0859_ _0859_/D _0444_/A vssd1 vssd1 vccd1 vccd1 _0899_/Q sky130_fd_sc_hd__dlxtn_1
X_0928_ _0928_/D repeater84/X vssd1 vssd1 vccd1 vccd1 _0928_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0713_ _0705_/X _0706_/X _0808_/Q vssd1 vssd1 vccd1 vccd1 _0713_/X sky130_fd_sc_hd__a21o_1
X_0644_ _0644_/A vssd1 vssd1 vccd1 vccd1 _0916_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0575_ _0577_/A _0653_/B vssd1 vssd1 vccd1 vccd1 _0576_/A sky130_fd_sc_hd__and2_1
XFILLER_25_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0758__B _0758_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput37 _0406_/C vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
Xoutput59 _0832_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
Xoutput48 _0835_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
XFILLER_16_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0668__B _0668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0558_ _0566_/A _0614_/B vssd1 vssd1 vccd1 vccd1 _0559_/A sky130_fd_sc_hd__and2_1
XFILLER_7_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0627_ _0649_/A _0627_/B vssd1 vssd1 vccd1 vccd1 _0628_/A sky130_fd_sc_hd__and2_1
XFILLER_26_424 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0489_ _0489_/A vssd1 vssd1 vccd1 vccd1 _0851_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input14_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater67 _0447_/A vssd1 vssd1 vccd1 vccd1 _0449_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_8_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater78 _0927_/Q vssd1 vssd1 vccd1 vccd1 _1140_/A sky130_fd_sc_hd__clkbuf_2
Xrepeater89 _0822_/Q vssd1 vssd1 vccd1 vccd1 _0433_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__0679__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0805__CLK _0829_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0412_ _0756_/A _0925_/Q _0434_/A vssd1 vssd1 vccd1 vccd1 _0413_/C sky130_fd_sc_hd__a21oi_1
Xpixel_macro_224 vssd1 vssd1 vccd1 vccd1 pixel_macro_224/HI la_data_out[73] sky130_fd_sc_hd__conb_1
Xpixel_macro_213 vssd1 vssd1 vccd1 vccd1 pixel_macro_213/HI la_data_out[62] sky130_fd_sc_hd__conb_1
Xpixel_macro_202 vssd1 vssd1 vccd1 vccd1 pixel_macro_202/HI la_data_out[51] sky130_fd_sc_hd__conb_1
XFILLER_23_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xpixel_macro_279 vssd1 vssd1 vccd1 vccd1 pixel_macro_279/HI wbs_dat_o[15] sky130_fd_sc_hd__conb_1
Xpixel_macro_268 vssd1 vssd1 vccd1 vccd1 pixel_macro_268/HI la_data_out[117] sky130_fd_sc_hd__conb_1
Xpixel_macro_235 vssd1 vssd1 vccd1 vccd1 pixel_macro_235/HI la_data_out[84] sky130_fd_sc_hd__conb_1
Xpixel_macro_257 vssd1 vssd1 vccd1 vccd1 pixel_macro_257/HI la_data_out[106] sky130_fd_sc_hd__conb_1
Xpixel_macro_246 vssd1 vssd1 vccd1 vccd1 pixel_macro_246/HI la_data_out[95] sky130_fd_sc_hd__conb_1
XANTENNA_input6_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_232 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0828__CLK _0839_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0892_ _0892_/D repeater68/X vssd1 vssd1 vccd1 vccd1 _0897_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0875_ _0875_/D repeater69/X vssd1 vssd1 vccd1 vccd1 _0913_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA__0695__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_544 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0660_ _0660_/A vssd1 vssd1 vccd1 vccd1 _0896_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0591_ _0591_/A vssd1 vssd1 vccd1 vccd1 _0885_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__0687__A _0706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0927_ _0927_/D repeater82/X vssd1 vssd1 vccd1 vccd1 _0927_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA__0597__A _0605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0789_ _0910_/Q _0777_/X _0788_/X _0781_/X vssd1 vssd1 vccd1 vccd1 _0836_/D sky130_fd_sc_hd__o211a_1
X_0858_ _0858_/D repeater71/X vssd1 vssd1 vccd1 vccd1 _0910_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0712_ input22/X _0704_/X _0711_/X _0700_/X vssd1 vssd1 vccd1 vccd1 _0807_/D sky130_fd_sc_hd__o211a_1
X_0574_ _0574_/A vssd1 vssd1 vccd1 vccd1 _0866_/D sky130_fd_sc_hd__clkbuf_1
X_0643_ _0661_/A _0643_/B vssd1 vssd1 vccd1 vccd1 _0644_/A sky130_fd_sc_hd__and2_1
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0929__GATE_N repeater82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput38 _0474_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
Xoutput49 _0836_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0626_ _0626_/A vssd1 vssd1 vccd1 vccd1 _0914_/D sky130_fd_sc_hd__clkbuf_1
X_0557_ _0579_/A vssd1 vssd1 vccd1 vccd1 _0566_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_436 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0488_ _0500_/A _0614_/B vssd1 vssd1 vccd1 vccd1 _0489_/A sky130_fd_sc_hd__and2_1
XFILLER_21_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater79 _0926_/Q vssd1 vssd1 vccd1 vccd1 _0579_/A sky130_fd_sc_hd__clkbuf_2
Xrepeater68 _0435_/Y vssd1 vssd1 vccd1 vccd1 repeater68/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0411_ _0426_/A vssd1 vssd1 vccd1 vccd1 _0756_/A sky130_fd_sc_hd__clkbuf_2
Xpixel_macro_247 vssd1 vssd1 vccd1 vccd1 pixel_macro_247/HI la_data_out[96] sky130_fd_sc_hd__conb_1
Xpixel_macro_214 vssd1 vssd1 vccd1 vccd1 pixel_macro_214/HI la_data_out[63] sky130_fd_sc_hd__conb_1
Xpixel_macro_203 vssd1 vssd1 vccd1 vccd1 pixel_macro_203/HI la_data_out[52] sky130_fd_sc_hd__conb_1
Xpixel_macro_225 vssd1 vssd1 vccd1 vccd1 pixel_macro_225/HI la_data_out[74] sky130_fd_sc_hd__conb_1
Xpixel_macro_236 vssd1 vssd1 vccd1 vccd1 pixel_macro_236/HI la_data_out[85] sky130_fd_sc_hd__conb_1
XFILLER_23_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_491 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xpixel_macro_258 vssd1 vssd1 vccd1 vccd1 pixel_macro_258/HI la_data_out[107] sky130_fd_sc_hd__conb_1
Xpixel_macro_269 vssd1 vssd1 vccd1 vccd1 pixel_macro_269/HI la_data_out[118] sky130_fd_sc_hd__conb_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0609_ _0609_/A _0645_/B vssd1 vssd1 vccd1 vccd1 _0610_/A sky130_fd_sc_hd__and2_1
XFILLER_26_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0891_ _0891_/D repeater63/X vssd1 vssd1 vccd1 vccd1 _0915_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_9_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output38_A _0474_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0874_ _0874_/D repeater66/X vssd1 vssd1 vccd1 vccd1 _0912_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_9_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0818__CLK _0829_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0590_ _0594_/A _0618_/B vssd1 vssd1 vccd1 vccd1 _0591_/A sky130_fd_sc_hd__and2_1
XFILLER_10_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0926_ _0926_/D repeater82/X vssd1 vssd1 vccd1 vccd1 _0926_/Q sky130_fd_sc_hd__dlxtn_1
X_0857_ _0857_/D repeater68/X vssd1 vssd1 vccd1 vccd1 _0897_/Q sky130_fd_sc_hd__dlxtn_1
X_0788_ _0836_/Q _0792_/B vssd1 vssd1 vccd1 vccd1 _0788_/X sky130_fd_sc_hd__or2_1
XFILLER_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0711_ _0705_/X _0706_/X _0807_/Q vssd1 vssd1 vccd1 vccd1 _0711_/X sky130_fd_sc_hd__a21o_1
X_0573_ _0577_/A _0643_/B vssd1 vssd1 vccd1 vccd1 _0574_/A sky130_fd_sc_hd__and2_1
X_0642_ _0927_/Q vssd1 vssd1 vccd1 vccd1 _0661_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput28 _0820_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
Xoutput39 _0821_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
X_0909_ _0909_/D repeater88/X vssd1 vssd1 vccd1 vccd1 _0917_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA__0401__A _0821_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0625_ _0649_/A _0625_/B vssd1 vssd1 vccd1 vccd1 _0626_/A sky130_fd_sc_hd__and2_1
XFILLER_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0556_ _0556_/A vssd1 vssd1 vccd1 vccd1 _0865_/D sky130_fd_sc_hd__clkbuf_1
X_0487_ _0632_/B vssd1 vssd1 vccd1 vccd1 _0614_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_26_448 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater69 _0428_/A vssd1 vssd1 vccd1 vccd1 repeater69/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_603 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0410_ _0400_/B _0413_/B _0409_/Y vssd1 vssd1 vccd1 vccd1 _0822_/D sky130_fd_sc_hd__o21a_1
XFILLER_23_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xpixel_macro_237 vssd1 vssd1 vccd1 vccd1 pixel_macro_237/HI la_data_out[86] sky130_fd_sc_hd__conb_1
Xpixel_macro_226 vssd1 vssd1 vccd1 vccd1 pixel_macro_226/HI la_data_out[75] sky130_fd_sc_hd__conb_1
Xpixel_macro_215 vssd1 vssd1 vccd1 vccd1 pixel_macro_215/HI la_data_out[64] sky130_fd_sc_hd__conb_1
Xpixel_macro_204 vssd1 vssd1 vccd1 vccd1 pixel_macro_204/HI la_data_out[53] sky130_fd_sc_hd__conb_1
Xpixel_macro_248 vssd1 vssd1 vccd1 vccd1 pixel_macro_248/HI la_data_out[97] sky130_fd_sc_hd__conb_1
Xpixel_macro_259 vssd1 vssd1 vccd1 vccd1 pixel_macro_259/HI la_data_out[108] sky130_fd_sc_hd__conb_1
XANTENNA__0789__A1 _0910_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0608_ _0608_/A vssd1 vssd1 vccd1 vccd1 _0882_/D sky130_fd_sc_hd__clkbuf_1
X_0539_ _0539_/A vssd1 vssd1 vccd1 vccd1 _0861_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_256 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0890_ _0890_/D _0445_/X vssd1 vssd1 vccd1 vccd1 _0904_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_4_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0873_ _0873_/D repeater70/X vssd1 vssd1 vccd1 vccd1 _0911_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_24_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0404__A _0514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1141_ _1141_/A vssd1 vssd1 vccd1 vccd1 _1141_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0925_ _0925_/D repeater83/X vssd1 vssd1 vccd1 vccd1 _0925_/Q sky130_fd_sc_hd__dlxtn_1
X_0787_ _0907_/Q _0777_/X _0786_/X _0781_/X vssd1 vssd1 vccd1 vccd1 _0835_/D sky130_fd_sc_hd__o211a_1
X_0856_ _0856_/D repeater87/X vssd1 vssd1 vccd1 vccd1 _0917_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_24_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0761__C1 _0745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0710_ input21/X _0704_/X _0709_/X _0700_/X vssd1 vssd1 vccd1 vccd1 _0806_/D sky130_fd_sc_hd__o211a_1
X_0641_ _0641_/A vssd1 vssd1 vccd1 vccd1 _0900_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0808__CLK _0921_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0572_ _0572_/A vssd1 vssd1 vccd1 vccd1 _0873_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0908_ _0908_/D repeater64/X vssd1 vssd1 vccd1 vccd1 _0908_/Q sky130_fd_sc_hd__dlxtn_1
Xoutput29 _1140_/X vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
X_0839_ _0839_/CLK _0839_/D vssd1 vssd1 vccd1 vccd1 _0839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0743__C1 _0731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0734__C1 _0731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0502__A _0525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0624_ _0655_/A vssd1 vssd1 vccd1 vccd1 _0649_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__0725__C1 _0714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0555_ _0931_/Q _0918_/D vssd1 vssd1 vccd1 vccd1 _0556_/A sky130_fd_sc_hd__and2_1
X_0486_ _0514_/A _0486_/B vssd1 vssd1 vccd1 vccd1 _0632_/B sky130_fd_sc_hd__nor2_1
XFILLER_26_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_238 vssd1 vssd1 vccd1 vccd1 pixel_macro_238/HI la_data_out[87] sky130_fd_sc_hd__conb_1
Xpixel_macro_227 vssd1 vssd1 vccd1 vccd1 pixel_macro_227/HI la_data_out[76] sky130_fd_sc_hd__conb_1
Xpixel_macro_216 vssd1 vssd1 vccd1 vccd1 pixel_macro_216/HI la_data_out[65] sky130_fd_sc_hd__conb_1
Xpixel_macro_205 vssd1 vssd1 vccd1 vccd1 pixel_macro_205/HI la_data_out[54] sky130_fd_sc_hd__conb_1
Xpixel_macro_249 vssd1 vssd1 vccd1 vccd1 pixel_macro_249/HI la_data_out[98] sky130_fd_sc_hd__conb_1
XANTENNA__0410__A1 _0400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0538_ _0538_/A _0647_/B vssd1 vssd1 vccd1 vccd1 _0539_/A sky130_fd_sc_hd__and2_1
X_0607_ _0928_/Q _0627_/B vssd1 vssd1 vccd1 vccd1 _0608_/A sky130_fd_sc_hd__and2_1
X_0469_ _0817_/Q _0816_/Q _0815_/Q _0814_/Q vssd1 vssd1 vccd1 vccd1 _0470_/D sky130_fd_sc_hd__or4_1
XFILLER_26_268 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_603 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input12_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0872_ _0872_/D _0444_/A vssd1 vssd1 vccd1 vccd1 _0899_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0510__A _0510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0404__B _0510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0420__A _0821_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output43_A _0823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1140_ _1140_/A vssd1 vssd1 vccd1 vccd1 _1140_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0505__A _0519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0924_ _0924_/D repeater84/X vssd1 vssd1 vccd1 vccd1 _0924_/Q sky130_fd_sc_hd__dlxtn_1
X_0855_ _0855_/D repeater64/X vssd1 vssd1 vccd1 vccd1 _0908_/Q sky130_fd_sc_hd__dlxtn_1
X_0786_ _0835_/Q _0792_/B vssd1 vssd1 vccd1 vccd1 _0786_/X sky130_fd_sc_hd__or2_1
XFILLER_24_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_322 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0571_ _0577_/A _0622_/B vssd1 vssd1 vccd1 vccd1 _0572_/A sky130_fd_sc_hd__and2_1
X_0640_ _0640_/A _0640_/B vssd1 vssd1 vccd1 vccd1 _0641_/A sky130_fd_sc_hd__and2_1
X_0907_ _0907_/D _0450_/X vssd1 vssd1 vccd1 vccd1 _0907_/Q sky130_fd_sc_hd__dlxtn_1
X_0838_ _0838_/CLK _0838_/D vssd1 vssd1 vccd1 vccd1 _0838_/Q sky130_fd_sc_hd__dfxtp_1
X_0769_ _0917_/Q _0764_/X _0767_/X _0768_/X vssd1 vssd1 vccd1 vccd1 _0828_/D sky130_fd_sc_hd__o211a_1
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0623_ _0623_/A vssd1 vssd1 vccd1 vccd1 _0911_/D sky130_fd_sc_hd__clkbuf_1
X_0554_ _0554_/A vssd1 vssd1 vccd1 vccd1 _0862_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0485_ _0525_/A vssd1 vssd1 vccd1 vccd1 _0500_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0603__A _0605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_239 vssd1 vssd1 vccd1 vccd1 pixel_macro_239/HI la_data_out[88] sky130_fd_sc_hd__conb_1
Xpixel_macro_217 vssd1 vssd1 vccd1 vccd1 pixel_macro_217/HI la_data_out[66] sky130_fd_sc_hd__conb_1
Xpixel_macro_206 vssd1 vssd1 vccd1 vccd1 pixel_macro_206/HI la_data_out[55] sky130_fd_sc_hd__conb_1
Xpixel_macro_228 vssd1 vssd1 vccd1 vccd1 pixel_macro_228/HI la_data_out[77] sky130_fd_sc_hd__conb_1
X_0537_ _0537_/A vssd1 vssd1 vccd1 vccd1 _0854_/D sky130_fd_sc_hd__clkbuf_1
X_0606_ _0606_/A vssd1 vssd1 vccd1 vccd1 _0889_/D sky130_fd_sc_hd__clkbuf_1
X_0468_ _0813_/Q _0812_/Q _0811_/Q _0810_/Q vssd1 vssd1 vccd1 vccd1 _0470_/C sky130_fd_sc_hd__or4_2
X_0399_ _0822_/Q vssd1 vssd1 vccd1 vccd1 _0400_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0508__A _0519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0418__A _0438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0871_ _0871_/D repeater71/X vssd1 vssd1 vccd1 vccd1 _0910_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_27_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output36_A _0551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0854_ _0854_/D repeater62/X vssd1 vssd1 vccd1 vccd1 _0907_/Q sky130_fd_sc_hd__dlxtn_1
X_0923_ _0923_/D repeater82/X vssd1 vssd1 vccd1 vccd1 _0923_/Q sky130_fd_sc_hd__dlxtn_1
X_0785_ _0915_/Q _0777_/X _0784_/X _0781_/X vssd1 vssd1 vccd1 vccd1 _0834_/D sky130_fd_sc_hd__o211a_1
XFILLER_24_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0831__CLK _0921_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0431__A _0486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_584 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0570_ _0570_/A vssd1 vssd1 vccd1 vccd1 _0868_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0516__A _0519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0837_ _0838_/CLK _0837_/D vssd1 vssd1 vccd1 vccd1 _0837_/Q sky130_fd_sc_hd__dfxtp_1
X_0906_ _0906_/D _0417_/Y vssd1 vssd1 vccd1 vccd1 _0916_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA__0743__A1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0699_ _0781_/A vssd1 vssd1 vccd1 vccd1 _0731_/A sky130_fd_sc_hd__clkbuf_2
X_0768_ _0781_/A vssd1 vssd1 vccd1 vccd1 _0768_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0734__A1 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0725__A1 _0678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0622_ _0622_/A _0622_/B vssd1 vssd1 vccd1 vccd1 _0623_/A sky130_fd_sc_hd__and2_1
X_0484_ _0484_/A vssd1 vssd1 vccd1 vccd1 _0924_/D sky130_fd_sc_hd__clkbuf_1
X_0553_ _0931_/Q _0645_/B vssd1 vssd1 vccd1 vccd1 _0554_/A sky130_fd_sc_hd__and2_1
XFILLER_22_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_178 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0603__B _0653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_229 vssd1 vssd1 vccd1 vccd1 pixel_macro_229/HI la_data_out[78] sky130_fd_sc_hd__conb_1
Xpixel_macro_207 vssd1 vssd1 vccd1 vccd1 pixel_macro_207/HI la_data_out[56] sky130_fd_sc_hd__conb_1
Xpixel_macro_218 vssd1 vssd1 vccd1 vccd1 pixel_macro_218/HI la_data_out[67] sky130_fd_sc_hd__conb_1
XFILLER_7_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0536_ _0538_/A _0620_/B vssd1 vssd1 vccd1 vccd1 _0537_/A sky130_fd_sc_hd__and2_1
X_0605_ _0605_/A _0625_/B vssd1 vssd1 vccd1 vccd1 _0606_/A sky130_fd_sc_hd__and2_1
X_0467_ _0467_/A vssd1 vssd1 vccd1 vccd1 _0925_/D sky130_fd_sc_hd__clkbuf_1
X_0398_ _0823_/Q vssd1 vssd1 vccd1 vccd1 _0433_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0614__A _0622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0524__A _0655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0519_ _0519_/A _0625_/B vssd1 vssd1 vccd1 vccd1 _0520_/A sky130_fd_sc_hd__and2_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0609__A _0609_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0870_ _0870_/D repeater68/X vssd1 vssd1 vccd1 vccd1 _0897_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_9_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0519__A _0519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0922_ _0922_/D repeater83/X vssd1 vssd1 vccd1 vccd1 _0922_/Q sky130_fd_sc_hd__dlxtn_1
X_0853_ _0853_/D _0762_/A2 vssd1 vssd1 vccd1 vccd1 _0916_/Q sky130_fd_sc_hd__dlxtn_1
X_0784_ _0834_/Q _0792_/B vssd1 vssd1 vccd1 vccd1 _0784_/X sky130_fd_sc_hd__or2_1
Xinput1 wb_rst_i vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_2
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_90 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0746__C1 _0745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0622__A _0622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_596 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0516__B _0653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0532__A _0538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0905_ _0905_/D _0448_/X vssd1 vssd1 vccd1 vccd1 _0915_/Q sky130_fd_sc_hd__dlxtn_2
X_0836_ _0838_/CLK _0836_/D vssd1 vssd1 vccd1 vccd1 _0836_/Q sky130_fd_sc_hd__dfxtp_1
X_0767_ _0828_/Q _0767_/B vssd1 vssd1 vccd1 vccd1 _0767_/X sky130_fd_sc_hd__or2_1
X_0698_ _0690_/X _0691_/X _0803_/Q vssd1 vssd1 vccd1 vccd1 _0698_/X sky130_fd_sc_hd__a21o_1
XFILLER_24_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0621_ _0621_/A vssd1 vssd1 vccd1 vccd1 _0907_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0821__CLK _0921_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0552_ _0552_/A vssd1 vssd1 vccd1 vccd1 _0856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0483_ _0483_/A _0483_/B _0483_/C vssd1 vssd1 vccd1 vccd1 _0484_/A sky130_fd_sc_hd__and3_1
XFILLER_21_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0819_ _0829_/CLK _0819_/D vssd1 vssd1 vccd1 vccd1 _0819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_419 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_219 vssd1 vssd1 vccd1 vccd1 pixel_macro_219/HI la_data_out[68] sky130_fd_sc_hd__conb_1
Xpixel_macro_208 vssd1 vssd1 vccd1 vccd1 pixel_macro_208/HI la_data_out[57] sky130_fd_sc_hd__conb_1
XFILLER_7_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0604_ _0604_/A vssd1 vssd1 vccd1 vccd1 _0884_/D sky130_fd_sc_hd__clkbuf_1
X_0466_ _0466_/A _0466_/B _0476_/B vssd1 vssd1 vccd1 vccd1 _0467_/A sky130_fd_sc_hd__and3_1
X_0535_ _0535_/A vssd1 vssd1 vccd1 vccd1 _0859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0899__GATE_N _0436_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0540__A _0551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0518_ _0664_/B vssd1 vssd1 vccd1 vccd1 _0625_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0449_ _0668_/B _0449_/B _0657_/B vssd1 vssd1 vccd1 vccd1 _0450_/A sky130_fd_sc_hd__or3_1
XFILLER_2_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input10_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0625__A _0649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input2_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0921_ _0921_/CLK _0924_/Q _0798_/Y vssd1 vssd1 vccd1 vccd1 _0921_/Q sky130_fd_sc_hd__dfrtp_1
X_0852_ _0852_/D repeater63/X vssd1 vssd1 vccd1 vccd1 _0915_/Q sky130_fd_sc_hd__dlxtn_2
X_0783_ _0794_/B vssd1 vssd1 vccd1 vccd1 _0792_/B sky130_fd_sc_hd__clkbuf_1
Xinput2 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_91 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output41_A _0918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0904_ _0904_/D _0445_/X vssd1 vssd1 vccd1 vccd1 _0904_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA__0532__B _0560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0697_ input17/X _0689_/X _0696_/X _0680_/X vssd1 vssd1 vccd1 vccd1 _0802_/D sky130_fd_sc_hd__o211a_1
X_0835_ _0838_/CLK _0835_/D vssd1 vssd1 vccd1 vccd1 _0835_/Q sky130_fd_sc_hd__dfxtp_1
X_0766_ _0916_/Q _0764_/X _0765_/X _0745_/X vssd1 vssd1 vccd1 vccd1 _0827_/D sky130_fd_sc_hd__o211a_1
XFILLER_24_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0723__A _0737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0620_ _0622_/A _0620_/B vssd1 vssd1 vccd1 vccd1 _0621_/A sky130_fd_sc_hd__and2_1
XFILLER_7_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0551_ _0551_/A _0627_/B vssd1 vssd1 vccd1 vccd1 _0552_/A sky130_fd_sc_hd__and2_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0482_ _0927_/D _0474_/Y _0479_/Y vssd1 vssd1 vccd1 vccd1 _0923_/D sky130_fd_sc_hd__a21o_1
XFILLER_3_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0543__A _0549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0818_ _0829_/CLK _0818_/D vssd1 vssd1 vccd1 vccd1 _0818_/Q sky130_fd_sc_hd__dfxtp_1
X_0749_ input1/X vssd1 vssd1 vccd1 vccd1 _0797_/A sky130_fd_sc_hd__buf_2
XFILLER_16_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xpixel_macro_209 vssd1 vssd1 vccd1 vccd1 pixel_macro_209/HI la_data_out[58] sky130_fd_sc_hd__conb_1
X_0534_ _0538_/A _0618_/B vssd1 vssd1 vccd1 vccd1 _0535_/A sky130_fd_sc_hd__and2_1
XFILLER_7_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0603_ _0605_/A _0653_/B vssd1 vssd1 vccd1 vccd1 _0604_/A sky130_fd_sc_hd__and2_1
XANTENNA__0538__A _0538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0465_ _0931_/D vssd1 vssd1 vccd1 vccd1 _0930_/D sky130_fd_sc_hd__inv_2
XFILLER_22_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0720__B _0737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0448__A _0448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0811__CLK _0839_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0517_ _0517_/A vssd1 vssd1 vccd1 vccd1 _0845_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0448_ _0448_/A vssd1 vssd1 vccd1 vccd1 _0448_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0834__CLK _0838_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0731__A _0731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0551__A _0551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0636__A _0640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0920_ _0921_/CLK _0923_/Q _0797_/Y vssd1 vssd1 vccd1 vccd1 _0920_/Q sky130_fd_sc_hd__dfrtp_1
X_0851_ _0851_/D repeater65/X vssd1 vssd1 vccd1 vccd1 _0904_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0782_ _0912_/Q _0777_/X _0780_/X _0781_/X vssd1 vssd1 vccd1 vccd1 _0833_/D sky130_fd_sc_hd__o211a_1
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput3 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XTAP_92 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0746__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output34_A _0579_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0903_ _0903_/D _0439_/B vssd1 vssd1 vccd1 vccd1 _0914_/Q sky130_fd_sc_hd__dlxtn_1
X_0834_ _0838_/CLK _0834_/D vssd1 vssd1 vccd1 vccd1 _0834_/Q sky130_fd_sc_hd__dfxtp_1
X_0765_ _0827_/Q _0767_/B vssd1 vssd1 vccd1 vccd1 _0765_/X sky130_fd_sc_hd__or2_1
X_0696_ _0690_/X _0691_/X _0802_/Q vssd1 vssd1 vccd1 vccd1 _0696_/X sky130_fd_sc_hd__a21o_1
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0918__CLK _0921_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0550_ _0550_/A vssd1 vssd1 vccd1 vccd1 _0863_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0481_ _0475_/Y _0478_/X _0479_/Y _0480_/X vssd1 vssd1 vccd1 vccd1 _0922_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_19_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0817_ _0829_/CLK _0817_/D vssd1 vssd1 vccd1 vccd1 _0817_/Q sky130_fd_sc_hd__dfxtp_1
X_0679_ input1/X vssd1 vssd1 vccd1 vccd1 _0781_/A sky130_fd_sc_hd__inv_2
X_0748_ input24/X _0735_/X _0747_/X _0745_/X vssd1 vssd1 vccd1 vccd1 _0819_/D sky130_fd_sc_hd__o211a_1
XFILLER_16_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0602_ _0602_/A vssd1 vssd1 vccd1 vccd1 _0879_/D sky130_fd_sc_hd__clkbuf_1
X_0533_ _0533_/A vssd1 vssd1 vccd1 vccd1 _0857_/D sky130_fd_sc_hd__clkbuf_1
X_0464_ _0466_/B _0476_/B vssd1 vssd1 vccd1 vccd1 _0931_/D sky130_fd_sc_hd__nor2_1
XFILLER_19_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0549__A _0549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0447_ _0447_/A _0657_/B vssd1 vssd1 vccd1 vccd1 _0448_/A sky130_fd_sc_hd__or2_1
X_0516_ _0519_/A _0653_/B vssd1 vssd1 vccd1 vccd1 _0517_/A sky130_fd_sc_hd__and2_1
XFILLER_22_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0459__A _0929_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0801__CLK _0838_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0850_ _0850_/D repeater85/X vssd1 vssd1 vccd1 vccd1 _0914_/Q sky130_fd_sc_hd__dlxtn_1
X_0781_ _0781_/A vssd1 vssd1 vccd1 vccd1 _0781_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0824__CLK _0839_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput4 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XTAP_93 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_60 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0562__A _0566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0737__A _0737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_190 vssd1 vssd1 vccd1 vccd1 pixel_macro_190/HI la_data_out[39] sky130_fd_sc_hd__conb_1
XFILLER_7_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0647__A _0649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0833_ _0838_/CLK _0833_/D vssd1 vssd1 vccd1 vccd1 _0833_/Q sky130_fd_sc_hd__dfxtp_1
X_0902_ _0902_/D repeater69/X vssd1 vssd1 vccd1 vccd1 _0913_/Q sky130_fd_sc_hd__dlxtn_1
X_0764_ _0764_/A vssd1 vssd1 vccd1 vccd1 _0764_/X sky130_fd_sc_hd__clkbuf_2
X_0695_ input16/X _0689_/X _0694_/X _0680_/X vssd1 vssd1 vccd1 vccd1 _0801_/D sky130_fd_sc_hd__o211a_1
XANTENNA__0557__A _0579_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0407__A1 _0400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0480_ _0466_/A _0483_/A _0474_/A _0478_/X vssd1 vssd1 vccd1 vccd1 _0480_/X sky130_fd_sc_hd__a31o_1
XFILLER_7_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0747_ _0736_/X _0737_/X _0819_/Q vssd1 vssd1 vccd1 vccd1 _0747_/X sky130_fd_sc_hd__a21o_1
X_0816_ _0829_/CLK _0816_/D vssd1 vssd1 vccd1 vccd1 _0816_/Q sky130_fd_sc_hd__dfxtp_1
X_0678_ _0678_/A _0754_/B _0678_/C _0678_/D vssd1 vssd1 vccd1 vccd1 _0678_/X sky130_fd_sc_hd__or4_1
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input26_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0601_ _0605_/A _0643_/B vssd1 vssd1 vccd1 vccd1 _0602_/A sky130_fd_sc_hd__and2_1
XFILLER_21_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0463_ _0928_/D vssd1 vssd1 vccd1 vccd1 _0927_/D sky130_fd_sc_hd__inv_2
X_0532_ _0538_/A _0560_/B vssd1 vssd1 vccd1 vccd1 _0533_/A sky130_fd_sc_hd__and2_1
XFILLER_19_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0446_ _0446_/A _0495_/B vssd1 vssd1 vccd1 vccd1 _0657_/B sky130_fd_sc_hd__nor2_1
X_0515_ _0661_/B vssd1 vssd1 vccd1 vccd1 _0653_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0475__A _0799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output57_A _0830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0429_ _0429_/A vssd1 vssd1 vccd1 vccd1 _0429_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0780_ _0833_/Q _0780_/B vssd1 vssd1 vccd1 vccd1 _0780_/X sky130_fd_sc_hd__or2_1
Xinput5 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_72 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_94 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0799__CLK _0838_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0753__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_191 vssd1 vssd1 vccd1 vccd1 pixel_macro_191/HI la_data_out[40] sky130_fd_sc_hd__conb_1
Xpixel_macro_180 vssd1 vssd1 vccd1 vccd1 pixel_macro_180/HI la_data_out[29] sky130_fd_sc_hd__conb_1
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0901_ _0901_/D _0447_/A vssd1 vssd1 vccd1 vccd1 _0912_/Q sky130_fd_sc_hd__dlxtn_1
X_0763_ _0826_/Q _0767_/B _0762_/X _0745_/X vssd1 vssd1 vccd1 vccd1 _0826_/D sky130_fd_sc_hd__o211a_1
X_0832_ _0838_/CLK _0832_/D vssd1 vssd1 vccd1 vccd1 _0832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0694_ _0690_/X _0691_/X _0801_/Q vssd1 vssd1 vccd1 vccd1 _0694_/X sky130_fd_sc_hd__a21o_1
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0573__A _0577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0814__CLK _0839_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0671__A_N input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0815_ _0829_/CLK _0815_/D vssd1 vssd1 vccd1 vccd1 _0815_/Q sky130_fd_sc_hd__dfxtp_1
X_0746_ input23/X _0735_/X _0744_/X _0745_/X vssd1 vssd1 vccd1 vccd1 _0818_/D sky130_fd_sc_hd__o211a_1
XANTENNA__0568__A _0579_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0677_ _0754_/B _0678_/C _0678_/D vssd1 vssd1 vccd1 vccd1 _0677_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__0837__CLK _0838_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input19_A wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0531_ _0531_/A vssd1 vssd1 vccd1 vccd1 _0864_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0600_ _0600_/A vssd1 vssd1 vccd1 vccd1 _0886_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0462_ _0462_/A vssd1 vssd1 vccd1 vccd1 _0928_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_250 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0729_ input17/X _0721_/X _0728_/X _0714_/X vssd1 vssd1 vccd1 vccd1 _0812_/D sky130_fd_sc_hd__o211a_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _0921_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0655__B _0655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0785__A1 _0915_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0514_ _0514_/A _0514_/B vssd1 vssd1 vccd1 vccd1 _0661_/B sky130_fd_sc_hd__nor2_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0445_ _0445_/A vssd1 vssd1 vccd1 vccd1 _0445_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0776__A1 _0908_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0756__A _0756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0666__A _0756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater72_A _0436_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0428_ _0428_/A _0655_/B vssd1 vssd1 vccd1 vccd1 _0429_/A sky130_fd_sc_hd__or2_1
XFILLER_10_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0486__A _0514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput6 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_73 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_95 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_170 vssd1 vssd1 vccd1 vccd1 pixel_macro_170/HI la_data_out[5] sky130_fd_sc_hd__conb_1
Xpixel_macro_192 vssd1 vssd1 vccd1 vccd1 pixel_macro_192/HI la_data_out[41] sky130_fd_sc_hd__conb_1
Xpixel_macro_181 vssd1 vssd1 vccd1 vccd1 pixel_macro_181/HI la_data_out[30] sky130_fd_sc_hd__conb_1
XFILLER_23_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0900_ _0900_/D repeater70/X vssd1 vssd1 vccd1 vccd1 _0911_/Q sky130_fd_sc_hd__dlxtn_1
X_0693_ _0678_/A _0689_/X _0692_/X _0680_/X vssd1 vssd1 vccd1 vccd1 _0800_/D sky130_fd_sc_hd__o211a_1
X_0762_ _0756_/B _0762_/A2 _0767_/B vssd1 vssd1 vccd1 vccd1 _0762_/X sky130_fd_sc_hd__a21bo_1
X_0831_ _0921_/CLK _0831_/D vssd1 vssd1 vccd1 vccd1 _0831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_26 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output32_A _1141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0814_ _0839_/CLK _0814_/D vssd1 vssd1 vccd1 vccd1 _0814_/Q sky130_fd_sc_hd__dfxtp_1
Xinput20 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_2
X_0676_ input9/X _0676_/B _0719_/C _0676_/D vssd1 vssd1 vccd1 vccd1 _0678_/D sky130_fd_sc_hd__or4_1
X_0745_ _0781_/A vssd1 vssd1 vccd1 vccd1 _0745_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_2__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _0829_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_479 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0530_ _0538_/A _0614_/B vssd1 vssd1 vccd1 vccd1 _0531_/A sky130_fd_sc_hd__and2_1
X_0461_ _0920_/Q _0466_/B _0921_/Q vssd1 vssd1 vccd1 vccd1 _0462_/A sky130_fd_sc_hd__or3_1
XFILLER_19_262 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0579__A _0579_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0659_ _0661_/A _0659_/B vssd1 vssd1 vccd1 vccd1 _0660_/A sky130_fd_sc_hd__and2_1
XANTENNA__0804__CLK _0829_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0728_ _0722_/X _0723_/X _0812_/Q vssd1 vssd1 vccd1 vccd1 _0728_/X sky130_fd_sc_hd__a21o_1
XANTENNA__0712__C1 _0700_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0703__C1 _0700_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0827__CLK _0839_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0444_ _0444_/A _0636_/B vssd1 vssd1 vccd1 vccd1 _0445_/A sky130_fd_sc_hd__or2_1
X_0513_ _0513_/A vssd1 vssd1 vccd1 vccd1 _0840_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0756__B _0756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0427_ _0486_/B _0503_/B vssd1 vssd1 vccd1 vccd1 _0655_/B sky130_fd_sc_hd__nor2_2
XFILLER_24_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0486__B _0486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
XTAP_74 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_96 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_160 vssd1 vssd1 vccd1 vccd1 pixel_macro_160/HI io_out[32] sky130_fd_sc_hd__conb_1
XFILLER_27_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_193 vssd1 vssd1 vccd1 vccd1 pixel_macro_193/HI la_data_out[42] sky130_fd_sc_hd__conb_1
Xpixel_macro_171 vssd1 vssd1 vccd1 vccd1 pixel_macro_171/HI la_data_out[6] sky130_fd_sc_hd__conb_1
Xpixel_macro_182 vssd1 vssd1 vccd1 vccd1 pixel_macro_182/HI la_data_out[31] sky130_fd_sc_hd__conb_1
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0497__A _0500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0830_ _0838_/CLK _0830_/D vssd1 vssd1 vccd1 vccd1 _0830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_591 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0692_ _0690_/X _0691_/X _0800_/Q vssd1 vssd1 vccd1 vccd1 _0692_/X sky130_fd_sc_hd__a21o_1
X_0761_ _0764_/A _0756_/X _0760_/X _0745_/X vssd1 vssd1 vccd1 vccd1 _0825_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_2_1__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _0838_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_38 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0483__C _0483_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput10 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 _0676_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__0690__A _0705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0813_ _0839_/CLK _0813_/D vssd1 vssd1 vccd1 vccd1 _0813_/Q sky130_fd_sc_hd__dfxtp_1
Xinput21 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_2
X_0744_ _0736_/X _0737_/X _0818_/Q vssd1 vssd1 vccd1 vccd1 _0744_/X sky130_fd_sc_hd__a21o_1
X_0675_ input6/X _0685_/A _0685_/B _0685_/C vssd1 vssd1 vccd1 vccd1 _0676_/D sky130_fd_sc_hd__or4_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0775__A _0831_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0460_ _0919_/Q vssd1 vssd1 vccd1 vccd1 _0466_/B sky130_fd_sc_hd__inv_2
XFILLER_19_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0727_ input16/X _0721_/X _0726_/X _0714_/X vssd1 vssd1 vccd1 vccd1 _0811_/D sky130_fd_sc_hd__o211a_1
XFILLER_8_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0658_ _0658_/A vssd1 vssd1 vccd1 vccd1 _0901_/D sky130_fd_sc_hd__clkbuf_1
X_0589_ _0589_/A vssd1 vssd1 vccd1 vccd1 _0883_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input24_A wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0482__A2 _0474_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0512_ _0519_/A _0643_/B vssd1 vssd1 vccd1 vccd1 _0513_/A sky130_fd_sc_hd__and2_1
X_0443_ _0514_/A _0446_/A vssd1 vssd1 vccd1 vccd1 _0636_/B sky130_fd_sc_hd__nor2_1
XANTENNA__0921__CLK _0921_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0697__C1 _0680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0426_ _0426_/A _0434_/A vssd1 vssd1 vccd1 vccd1 _0486_/B sky130_fd_sc_hd__or2b_2
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0817__CLK _0829_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0820__SET_B _0680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_0__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _0839_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_75 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_97 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0409_ _0400_/B _0413_/B _0918_/Q vssd1 vssd1 vccd1 vccd1 _0409_/Y sky130_fd_sc_hd__a21oi_1
Xpixel_macro_161 vssd1 vssd1 vccd1 vccd1 pixel_macro_161/HI io_out[33] sky130_fd_sc_hd__conb_1
Xpixel_macro_150 vssd1 vssd1 vccd1 vccd1 pixel_macro_150/HI io_out[22] sky130_fd_sc_hd__conb_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_183 vssd1 vssd1 vccd1 vccd1 pixel_macro_183/HI la_data_out[32] sky130_fd_sc_hd__conb_1
Xpixel_macro_194 vssd1 vssd1 vccd1 vccd1 pixel_macro_194/HI la_data_out[43] sky130_fd_sc_hd__conb_1
Xpixel_macro_172 vssd1 vssd1 vccd1 vccd1 pixel_macro_172/HI la_data_out[7] sky130_fd_sc_hd__conb_1
XFILLER_2_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0760_ _0825_/Q _0767_/B vssd1 vssd1 vccd1 vccd1 _0760_/X sky130_fd_sc_hd__or2_1
XANTENNA__0688__A _0705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0691_ _0736_/A vssd1 vssd1 vccd1 vccd1 _0691_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0889_ _0889_/D repeater85/X vssd1 vssd1 vccd1 vccd1 _0914_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput11 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 _0685_/A sky130_fd_sc_hd__clkbuf_1
Xinput22 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_2
X_0743_ input22/X _0735_/X _0742_/X _0731_/X vssd1 vssd1 vccd1 vccd1 _0817_/D sky130_fd_sc_hd__o211a_1
X_0812_ _0838_/CLK _0812_/D vssd1 vssd1 vccd1 vccd1 _0812_/Q sky130_fd_sc_hd__dfxtp_1
X_0674_ input3/X input2/X vssd1 vssd1 vccd1 vccd1 _0719_/C sky130_fd_sc_hd__or2_1
XFILLER_16_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0726_ _0722_/X _0723_/X _0811_/Q vssd1 vssd1 vccd1 vccd1 _0726_/X sky130_fd_sc_hd__a21o_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0657_ _0661_/A _0657_/B vssd1 vssd1 vccd1 vccd1 _0658_/A sky130_fd_sc_hd__and2_1
XANTENNA__0712__A1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0588_ _0594_/A _0634_/B vssd1 vssd1 vccd1 vccd1 _0589_/A sky130_fd_sc_hd__and2_1
XFILLER_27_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input17_A wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0703__A1 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0511_ _0651_/B vssd1 vssd1 vccd1 vccd1 _0643_/B sky130_fd_sc_hd__clkbuf_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0442_ _0442_/A vssd1 vssd1 vccd1 vccd1 _0442_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0430__A_N _0433_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0709_ _0705_/X _0706_/X _0806_/Q vssd1 vssd1 vccd1 vccd1 _0709_/X sky130_fd_sc_hd__a21o_1
XANTENNA_input9_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xpixel_macro_90 vssd1 vssd1 vccd1 vccd1 pixel_macro_90/HI io_oeb[0] sky130_fd_sc_hd__conb_1
XANTENNA__1140__A _1140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0425_ _0425_/A vssd1 vssd1 vccd1 vccd1 _0428_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_76 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_98 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_140 vssd1 vssd1 vccd1 vccd1 pixel_macro_140/HI io_out[12] sky130_fd_sc_hd__conb_1
X_0408_ _0406_/C _0560_/B _0407_/Y _0918_/Q vssd1 vssd1 vccd1 vccd1 _0823_/D sky130_fd_sc_hd__a211oi_1
Xpixel_macro_162 vssd1 vssd1 vccd1 vccd1 pixel_macro_162/HI io_out[34] sky130_fd_sc_hd__conb_1
Xpixel_macro_151 vssd1 vssd1 vccd1 vccd1 pixel_macro_151/HI io_out[23] sky130_fd_sc_hd__conb_1
XFILLER_11_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_173 vssd1 vssd1 vccd1 vccd1 pixel_macro_173/HI la_data_out[22] sky130_fd_sc_hd__conb_1
Xpixel_macro_195 vssd1 vssd1 vccd1 vccd1 pixel_macro_195/HI la_data_out[44] sky130_fd_sc_hd__conb_1
Xpixel_macro_184 vssd1 vssd1 vccd1 vccd1 pixel_macro_184/HI la_data_out[33] sky130_fd_sc_hd__conb_1
XFILLER_18_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0690_ _0705_/A vssd1 vssd1 vccd1 vccd1 _0690_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0888_ _0888_/D _0428_/A vssd1 vssd1 vccd1 vccd1 _0913_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0807__CLK _0921_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput12 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 _0685_/C sky130_fd_sc_hd__clkbuf_1
X_0673_ _0684_/A _0684_/B vssd1 vssd1 vccd1 vccd1 _0678_/C sky130_fd_sc_hd__nand2_1
X_0811_ _0839_/CLK _0811_/D vssd1 vssd1 vccd1 vccd1 _0811_/Q sky130_fd_sc_hd__dfxtp_1
X_0742_ _0736_/X _0737_/X _0817_/Q vssd1 vssd1 vccd1 vccd1 _0742_/X sky130_fd_sc_hd__a21o_1
Xinput23 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0402__A _0820_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0715__C1 _0714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0725_ _0678_/A _0721_/X _0724_/X _0714_/X vssd1 vssd1 vccd1 vccd1 _0810_/D sky130_fd_sc_hd__o211a_1
XFILLER_6_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0656_ _0656_/A vssd1 vssd1 vccd1 vccd1 _0913_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0587_ _0587_/A vssd1 vssd1 vccd1 vccd1 _0890_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1139_ _1141_/A vssd1 vssd1 vccd1 vccd1 _1139_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1138__A _1140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0510_ _0510_/A _0510_/B vssd1 vssd1 vccd1 vccd1 _0651_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0441_ _0441_/A _0495_/B vssd1 vssd1 vccd1 vccd1 _0442_/A sky130_fd_sc_hd__or2b_1
XFILLER_3_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0708_ input20/X _0704_/X _0707_/X _0700_/X vssd1 vssd1 vccd1 vccd1 _0805_/D sky130_fd_sc_hd__o211a_1
X_0639_ _0639_/A vssd1 vssd1 vccd1 vccd1 _0895_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0697__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xpixel_macro_91 vssd1 vssd1 vccd1 vccd1 pixel_macro_91/HI io_oeb[1] sky130_fd_sc_hd__conb_1
XFILLER_8_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0500__A _0500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0424_ _0451_/A _0640_/B _0666_/B vssd1 vssd1 vccd1 vccd1 _0425_/A sky130_fd_sc_hd__or3_1
XFILLER_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_77 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_99 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0407_ _0400_/B _0413_/B _0433_/A vssd1 vssd1 vccd1 vccd1 _0407_/Y sky130_fd_sc_hd__a21oi_1
Xpixel_macro_163 vssd1 vssd1 vccd1 vccd1 pixel_macro_163/HI io_out[35] sky130_fd_sc_hd__conb_1
Xpixel_macro_152 vssd1 vssd1 vccd1 vccd1 pixel_macro_152/HI io_out[24] sky130_fd_sc_hd__conb_1
Xpixel_macro_141 vssd1 vssd1 vccd1 vccd1 pixel_macro_141/HI io_out[13] sky130_fd_sc_hd__conb_1
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xpixel_macro_130 vssd1 vssd1 vccd1 vccd1 pixel_macro_130/HI io_out[2] sky130_fd_sc_hd__conb_1
Xpixel_macro_174 vssd1 vssd1 vccd1 vccd1 pixel_macro_174/HI la_data_out[23] sky130_fd_sc_hd__conb_1
Xpixel_macro_196 vssd1 vssd1 vccd1 vccd1 pixel_macro_196/HI la_data_out[45] sky130_fd_sc_hd__conb_1
Xpixel_macro_185 vssd1 vssd1 vccd1 vccd1 pixel_macro_185/HI la_data_out[34] sky130_fd_sc_hd__conb_1
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0887_ _0887_/D repeater66/X vssd1 vssd1 vccd1 vccd1 _0912_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput13 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 _0685_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_14_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0810_ _0839_/CLK _0810_/D vssd1 vssd1 vccd1 vccd1 _0810_/Q sky130_fd_sc_hd__dfxtp_1
X_0672_ _0758_/A _0758_/B vssd1 vssd1 vccd1 vccd1 _0754_/B sky130_fd_sc_hd__nand2_1
Xinput24 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0741_ input21/X _0735_/X _0740_/X _0731_/X vssd1 vssd1 vccd1 vccd1 _0816_/D sky130_fd_sc_hd__o211a_1
XFILLER_25_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0586_ _0594_/A _0614_/B vssd1 vssd1 vccd1 vccd1 _0587_/A sky130_fd_sc_hd__and2_1
XANTENNA__0503__A _0510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0655_ _0655_/A _0655_/B vssd1 vssd1 vccd1 vccd1 _0656_/A sky130_fd_sc_hd__and2_1
X_0724_ _0722_/X _0723_/X _0810_/Q vssd1 vssd1 vccd1 vccd1 _0724_/X sky130_fd_sc_hd__a21o_1
XFILLER_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1138_ _1140_/A vssd1 vssd1 vccd1 vccd1 _1138_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0413__A _0918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0440_ _0440_/A vssd1 vssd1 vccd1 vccd1 _0447_/A sky130_fd_sc_hd__clkbuf_1
X_0707_ _0705_/X _0706_/X _0805_/Q vssd1 vssd1 vccd1 vccd1 _0707_/X sky130_fd_sc_hd__a21o_1
X_0569_ _0577_/A _0649_/B vssd1 vssd1 vccd1 vccd1 _0570_/A sky130_fd_sc_hd__and2_1
X_0638_ _0640_/A _0638_/B vssd1 vssd1 vccd1 vccd1 _0639_/A sky130_fd_sc_hd__and2_1
XFILLER_26_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input22_A wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_92 vssd1 vssd1 vccd1 vccd1 pixel_macro_92/HI io_oeb[2] sky130_fd_sc_hd__conb_1
XFILLER_12_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0423_ _0514_/B _0503_/B vssd1 vssd1 vccd1 vccd1 _0666_/B sky130_fd_sc_hd__nor2_1
XFILLER_27_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_397 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0601__A _0605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_67 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_89 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0406_ _0434_/A _0426_/A _0406_/C vssd1 vssd1 vccd1 vccd1 _0413_/B sky130_fd_sc_hd__and3_1
Xpixel_macro_164 vssd1 vssd1 vccd1 vccd1 pixel_macro_164/HI io_out[36] sky130_fd_sc_hd__conb_1
Xpixel_macro_120 vssd1 vssd1 vccd1 vccd1 pixel_macro_120/HI io_oeb[30] sky130_fd_sc_hd__conb_1
Xpixel_macro_153 vssd1 vssd1 vccd1 vccd1 pixel_macro_153/HI io_out[25] sky130_fd_sc_hd__conb_1
Xpixel_macro_142 vssd1 vssd1 vccd1 vccd1 pixel_macro_142/HI io_out[14] sky130_fd_sc_hd__conb_1
XFILLER_27_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_131 vssd1 vssd1 vccd1 vccd1 pixel_macro_131/HI io_out[3] sky130_fd_sc_hd__conb_1
Xpixel_macro_197 vssd1 vssd1 vccd1 vccd1 pixel_macro_197/HI la_data_out[46] sky130_fd_sc_hd__conb_1
Xpixel_macro_186 vssd1 vssd1 vccd1 vccd1 pixel_macro_186/HI la_data_out[35] sky130_fd_sc_hd__conb_1
Xpixel_macro_175 vssd1 vssd1 vccd1 vccd1 pixel_macro_175/HI la_data_out[24] sky130_fd_sc_hd__conb_1
XFILLER_11_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0830__CLK _0838_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0886_ _0886_/D _0452_/X vssd1 vssd1 vccd1 vccd1 _0911_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_9_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0416__A _0823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 _0670_/B sky130_fd_sc_hd__clkbuf_1
Xinput25 wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 _0684_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0740_ _0736_/X _0737_/X _0816_/Q vssd1 vssd1 vccd1 vccd1 _0740_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0671_ input8/X input7/X input5/X input4/X vssd1 vssd1 vccd1 vccd1 _0758_/B sky130_fd_sc_hd__and4bb_1
XFILLER_25_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0869_ _0869_/D repeater87/X vssd1 vssd1 vccd1 vccd1 _0917_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_9_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0715__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0723_ _0737_/A vssd1 vssd1 vccd1 vccd1 _0723_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0654_ _0654_/A vssd1 vssd1 vccd1 vccd1 _0910_/D sky130_fd_sc_hd__clkbuf_1
X_0585_ _0609_/A vssd1 vssd1 vccd1 vccd1 _0594_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0514__A _0514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0706_ _0706_/A vssd1 vssd1 vccd1 vccd1 _0706_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0499_ _0657_/B vssd1 vssd1 vccd1 vccd1 _0647_/B sky130_fd_sc_hd__clkbuf_1
X_0568_ _0579_/A vssd1 vssd1 vccd1 vccd1 _0577_/A sky130_fd_sc_hd__clkbuf_2
X_0637_ _0637_/A vssd1 vssd1 vccd1 vccd1 _0899_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input15_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xpixel_macro_93 vssd1 vssd1 vccd1 vccd1 pixel_macro_93/HI io_oeb[3] sky130_fd_sc_hd__conb_1
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0422_ _0821_/Q _0820_/Q vssd1 vssd1 vccd1 vccd1 _0514_/B sky130_fd_sc_hd__or2_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input7_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0763__C1 _0745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_68 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0405_ _0634_/B vssd1 vssd1 vccd1 vccd1 _0560_/B sky130_fd_sc_hd__clkbuf_2
Xpixel_macro_165 vssd1 vssd1 vccd1 vccd1 pixel_macro_165/HI io_out[37] sky130_fd_sc_hd__conb_1
Xpixel_macro_121 vssd1 vssd1 vccd1 vccd1 pixel_macro_121/HI io_oeb[31] sky130_fd_sc_hd__conb_1
Xpixel_macro_154 vssd1 vssd1 vccd1 vccd1 pixel_macro_154/HI io_out[26] sky130_fd_sc_hd__conb_1
Xpixel_macro_110 vssd1 vssd1 vccd1 vccd1 pixel_macro_110/HI io_oeb[20] sky130_fd_sc_hd__conb_1
Xpixel_macro_143 vssd1 vssd1 vccd1 vccd1 pixel_macro_143/HI io_out[15] sky130_fd_sc_hd__conb_1
Xpixel_macro_132 vssd1 vssd1 vccd1 vccd1 pixel_macro_132/HI io_out[4] sky130_fd_sc_hd__conb_1
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xpixel_macro_198 vssd1 vssd1 vccd1 vccd1 pixel_macro_198/HI la_data_out[47] sky130_fd_sc_hd__conb_1
Xpixel_macro_176 vssd1 vssd1 vccd1 vccd1 pixel_macro_176/HI la_data_out[25] sky130_fd_sc_hd__conb_1
Xpixel_macro_187 vssd1 vssd1 vccd1 vccd1 pixel_macro_187/HI la_data_out[36] sky130_fd_sc_hd__conb_1
XANTENNA__0421__B _0446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0885_ _0885_/D _0436_/Y vssd1 vssd1 vccd1 vccd1 _0899_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA__0727__C1 _0714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0432__A _0668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput26 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _0670_/A sky130_fd_sc_hd__clkbuf_1
X_0670_ _0670_/A _0670_/B vssd1 vssd1 vccd1 vccd1 _0758_/A sky130_fd_sc_hd__and2_1
Xinput15 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 _0678_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0868_ _0868_/D _0429_/X vssd1 vssd1 vccd1 vccd1 _0908_/Q sky130_fd_sc_hd__dlxtn_1
X_0799_ _0838_/CLK _0799_/D vssd1 vssd1 vccd1 vccd1 _0799_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__0412__A1 _0756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0820__CLK _0921_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0427__A _0486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0653_ _0655_/A _0653_/B vssd1 vssd1 vccd1 vccd1 _0654_/A sky130_fd_sc_hd__and2_1
X_0722_ _0736_/A vssd1 vssd1 vccd1 vccd1 _0722_/X sky130_fd_sc_hd__clkbuf_2
X_0584_ _0584_/A vssd1 vssd1 vccd1 vccd1 _0878_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0620__A _0622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0530__A _0538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0636_ _0640_/A _0636_/B vssd1 vssd1 vccd1 vccd1 _0637_/A sky130_fd_sc_hd__and2_1
X_0705_ _0705_/A vssd1 vssd1 vccd1 vccd1 _0705_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0567_ _0567_/A vssd1 vssd1 vccd1 vccd1 _0874_/D sky130_fd_sc_hd__clkbuf_1
X_0498_ _0498_/A vssd1 vssd1 vccd1 vccd1 _0841_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0705__A _0705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xpixel_macro_94 vssd1 vssd1 vccd1 vccd1 pixel_macro_94/HI io_oeb[4] sky130_fd_sc_hd__conb_1
XFILLER_5_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0421_ _0503_/B _0446_/A vssd1 vssd1 vccd1 vccd1 _0640_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0525__A _0525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0619_ _0619_/A vssd1 vssd1 vccd1 vccd1 _0893_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0419__B _0433_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0435__A _0560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_69 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0404_ _0514_/A _0510_/A vssd1 vssd1 vccd1 vccd1 _0634_/B sky130_fd_sc_hd__nor2_1
Xpixel_macro_122 vssd1 vssd1 vccd1 vccd1 pixel_macro_122/HI io_oeb[32] sky130_fd_sc_hd__conb_1
Xpixel_macro_111 vssd1 vssd1 vccd1 vccd1 pixel_macro_111/HI io_oeb[21] sky130_fd_sc_hd__conb_1
Xpixel_macro_100 vssd1 vssd1 vccd1 vccd1 pixel_macro_100/HI io_oeb[10] sky130_fd_sc_hd__conb_1
Xpixel_macro_155 vssd1 vssd1 vccd1 vccd1 pixel_macro_155/HI io_out[27] sky130_fd_sc_hd__conb_1
Xpixel_macro_144 vssd1 vssd1 vccd1 vccd1 pixel_macro_144/HI io_out[16] sky130_fd_sc_hd__conb_1
Xpixel_macro_133 vssd1 vssd1 vccd1 vccd1 pixel_macro_133/HI io_out[5] sky130_fd_sc_hd__conb_1
Xpixel_macro_199 vssd1 vssd1 vccd1 vccd1 pixel_macro_199/HI la_data_out[48] sky130_fd_sc_hd__conb_1
Xpixel_macro_177 vssd1 vssd1 vccd1 vccd1 pixel_macro_177/HI la_data_out[26] sky130_fd_sc_hd__conb_1
Xpixel_macro_166 vssd1 vssd1 vccd1 vccd1 pixel_macro_166/HI irq[0] sky130_fd_sc_hd__conb_1
Xpixel_macro_188 vssd1 vssd1 vccd1 vccd1 pixel_macro_188/HI la_data_out[37] sky130_fd_sc_hd__conb_1
XFILLER_2_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0681__C1 _0680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0885__GATE_N _0436_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output39_A _0821_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0884_ _0884_/D _0442_/X vssd1 vssd1 vccd1 vccd1 _0910_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_5_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput27 wbs_we_i vssd1 vssd1 vccd1 vccd1 _0684_/A sky130_fd_sc_hd__clkbuf_1
Xinput16 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0412__A2 _0925_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0867_ _0867_/D repeater62/X vssd1 vssd1 vccd1 vccd1 _0907_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_0_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0798_ input1/X vssd1 vssd1 vccd1 vccd1 _0798_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0416__C_N _0821_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0479__A2 _0483_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0443__A _0514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0618__A _0622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0583_ _0926_/Q _0918_/D vssd1 vssd1 vccd1 vccd1 _0584_/A sky130_fd_sc_hd__and2_1
X_0721_ _0735_/A vssd1 vssd1 vccd1 vccd1 _0721_/X sky130_fd_sc_hd__clkbuf_2
X_0652_ _0652_/A vssd1 vssd1 vccd1 vccd1 _0906_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_280 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_0919_ _0921_/CLK _0922_/Q _0796_/Y vssd1 vssd1 vccd1 vccd1 _0919_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0438__A _0438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0810__CLK _0839_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0566_ _0566_/A _0647_/B vssd1 vssd1 vccd1 vccd1 _0567_/A sky130_fd_sc_hd__and2_1
X_0704_ _0704_/A vssd1 vssd1 vccd1 vccd1 _0704_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0635_ _0635_/A vssd1 vssd1 vccd1 vccd1 _0897_/D sky130_fd_sc_hd__clkbuf_1
X_0497_ _0500_/A _0620_/B vssd1 vssd1 vccd1 vccd1 _0498_/A sky130_fd_sc_hd__and2_1
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xpixel_macro_95 vssd1 vssd1 vccd1 vccd1 pixel_macro_95/HI io_oeb[5] sky130_fd_sc_hd__conb_1
XFILLER_12_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0833__CLK _0838_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0631__A _1140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0420_ _0821_/Q _0426_/A vssd1 vssd1 vccd1 vccd1 _0446_/A sky130_fd_sc_hd__or2b_1
XFILLER_23_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0541__A _0549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0549_ _0549_/A _0625_/B vssd1 vssd1 vccd1 vccd1 _0550_/A sky130_fd_sc_hd__and2_1
X_0618_ _0622_/A _0618_/B vssd1 vssd1 vccd1 vccd1 _0619_/A sky130_fd_sc_hd__and2_1
XFILLER_26_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input20_A wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_59 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0403_ _0434_/A _0426_/A vssd1 vssd1 vccd1 vccd1 _0510_/A sky130_fd_sc_hd__nand2_2
Xpixel_macro_123 vssd1 vssd1 vccd1 vccd1 pixel_macro_123/HI io_oeb[33] sky130_fd_sc_hd__conb_1
Xpixel_macro_156 vssd1 vssd1 vccd1 vccd1 pixel_macro_156/HI io_out[28] sky130_fd_sc_hd__conb_1
Xpixel_macro_112 vssd1 vssd1 vccd1 vccd1 pixel_macro_112/HI io_oeb[22] sky130_fd_sc_hd__conb_1
Xpixel_macro_145 vssd1 vssd1 vccd1 vccd1 pixel_macro_145/HI io_out[17] sky130_fd_sc_hd__conb_1
Xpixel_macro_101 vssd1 vssd1 vccd1 vccd1 pixel_macro_101/HI io_oeb[11] sky130_fd_sc_hd__conb_1
Xpixel_macro_134 vssd1 vssd1 vccd1 vccd1 pixel_macro_134/HI io_out[6] sky130_fd_sc_hd__conb_1
XFILLER_23_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0536__A _0538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xpixel_macro_167 vssd1 vssd1 vccd1 vccd1 pixel_macro_167/HI irq[1] sky130_fd_sc_hd__conb_1
Xpixel_macro_189 vssd1 vssd1 vccd1 vccd1 pixel_macro_189/HI la_data_out[38] sky130_fd_sc_hd__conb_1
Xpixel_macro_178 vssd1 vssd1 vccd1 vccd1 pixel_macro_178/HI la_data_out[27] sky130_fd_sc_hd__conb_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_175 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0446__A _0446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0727__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0883_ _0883_/D _0435_/Y vssd1 vssd1 vccd1 vccd1 _0897_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_24_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput17 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_159 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0866_ _0866_/D _0417_/Y vssd1 vssd1 vccd1 vccd1 _0916_/Q sky130_fd_sc_hd__dlxtn_1
X_0797_ _0797_/A vssd1 vssd1 vccd1 vccd1 _0797_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0443__B _0446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0634__A _0640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0720_ _0736_/A _0737_/A vssd1 vssd1 vccd1 vccd1 _0735_/A sky130_fd_sc_hd__nand2_1
XFILLER_7_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0651_ _0929_/Q _0651_/B vssd1 vssd1 vccd1 vccd1 _0652_/A sky130_fd_sc_hd__and2_1
XFILLER_6_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0582_ _0582_/A vssd1 vssd1 vccd1 vccd1 _0875_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_292 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0918_ _0921_/CLK _0918_/D vssd1 vssd1 vccd1 vccd1 _0918_/Q sky130_fd_sc_hd__dfxtp_2
X_0849_ _0849_/D repeater69/X vssd1 vssd1 vccd1 vccd1 _0913_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_0_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0927__GATE_N repeater82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0793__C1 _0731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0629__A _0649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0703_ input19/X _0689_/X _0702_/X _0700_/X vssd1 vssd1 vccd1 vccd1 _0804_/D sky130_fd_sc_hd__o211a_1
X_0565_ _0565_/A vssd1 vssd1 vccd1 vccd1 _0867_/D sky130_fd_sc_hd__clkbuf_1
X_0496_ _0638_/B vssd1 vssd1 vccd1 vccd1 _0620_/B sky130_fd_sc_hd__clkbuf_1
X_0634_ _0640_/A _0634_/B vssd1 vssd1 vccd1 vccd1 _0635_/A sky130_fd_sc_hd__and2_1
XFILLER_0_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0449__A _0668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xpixel_macro_96 vssd1 vssd1 vccd1 vccd1 pixel_macro_96/HI io_oeb[6] sky130_fd_sc_hd__conb_1
XFILLER_17_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0766__C1 _0745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0479_ _0483_/A _0483_/C _0483_/B vssd1 vssd1 vccd1 vccd1 _0479_/Y sky130_fd_sc_hd__a21boi_1
X_0548_ _0548_/A vssd1 vssd1 vccd1 vccd1 _0858_/D sky130_fd_sc_hd__clkbuf_1
X_0617_ _0617_/A vssd1 vssd1 vccd1 vccd1 _0892_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0748__C1 _0745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0800__CLK _0838_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input13_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_574 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0739__C1 _0731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0402_ _0820_/Q vssd1 vssd1 vccd1 vccd1 _0426_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xpixel_macro_124 vssd1 vssd1 vccd1 vccd1 pixel_macro_124/HI io_oeb[34] sky130_fd_sc_hd__conb_1
Xpixel_macro_157 vssd1 vssd1 vccd1 vccd1 pixel_macro_157/HI io_out[29] sky130_fd_sc_hd__conb_1
Xpixel_macro_113 vssd1 vssd1 vccd1 vccd1 pixel_macro_113/HI io_oeb[23] sky130_fd_sc_hd__conb_1
Xpixel_macro_146 vssd1 vssd1 vccd1 vccd1 pixel_macro_146/HI io_out[18] sky130_fd_sc_hd__conb_1
Xpixel_macro_102 vssd1 vssd1 vccd1 vccd1 pixel_macro_102/HI io_oeb[12] sky130_fd_sc_hd__conb_1
Xpixel_macro_135 vssd1 vssd1 vccd1 vccd1 pixel_macro_135/HI io_out[7] sky130_fd_sc_hd__conb_1
XFILLER_23_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xpixel_macro_168 vssd1 vssd1 vccd1 vccd1 pixel_macro_168/HI irq[2] sky130_fd_sc_hd__conb_1
Xpixel_macro_179 vssd1 vssd1 vccd1 vccd1 pixel_macro_179/HI la_data_out[28] sky130_fd_sc_hd__conb_1
XFILLER_23_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0823__CLK _0921_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input5_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0681__A1 _0799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_327 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0882_ _0882_/D repeater87/X vssd1 vssd1 vccd1 vccd1 _0917_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA__0547__A _0549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0415__A1 _0756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0865_ _0865_/D repeater63/X vssd1 vssd1 vccd1 vccd1 _0915_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_9_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0796_ _0797_/A vssd1 vssd1 vccd1 vccd1 _0796_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0923__GATE_N repeater82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0650_ _0650_/A vssd1 vssd1 vccd1 vccd1 _0908_/D sky130_fd_sc_hd__clkbuf_1
X_0581_ _0926_/Q _0645_/B vssd1 vssd1 vccd1 vccd1 _0582_/A sky130_fd_sc_hd__and2_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0560__A _0566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0848_ _0848_/D repeater66/X vssd1 vssd1 vccd1 vccd1 _0912_/Q sky130_fd_sc_hd__dlxtn_1
X_0917_ _0917_/D repeater88/X vssd1 vssd1 vccd1 vccd1 _0917_/Q sky130_fd_sc_hd__dlxtn_1
X_0779_ _0914_/Q _0777_/X _0778_/X _0768_/X vssd1 vssd1 vccd1 vccd1 _0832_/D sky130_fd_sc_hd__o211a_1
XFILLER_17_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0629__B _0668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0645__A _0661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0633_ _0633_/A vssd1 vssd1 vccd1 vccd1 _0904_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0702_ _0690_/X _0691_/X _0804_/Q vssd1 vssd1 vccd1 vccd1 _0702_/X sky130_fd_sc_hd__a21o_1
XFILLER_7_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0564_ _0566_/A _0620_/B vssd1 vssd1 vccd1 vccd1 _0565_/A sky130_fd_sc_hd__and2_1
X_0495_ _0510_/A _0495_/B vssd1 vssd1 vccd1 vccd1 _0638_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_97 vssd1 vssd1 vccd1 vccd1 pixel_macro_97/HI io_oeb[7] sky130_fd_sc_hd__conb_1
XFILLER_25_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0616_ _0622_/A _0634_/B vssd1 vssd1 vccd1 vccd1 _0617_/A sky130_fd_sc_hd__and2_1
X_0478_ _0466_/A _0476_/Y _0477_/X vssd1 vssd1 vccd1 vccd1 _0478_/X sky130_fd_sc_hd__a21o_1
X_0547_ _0549_/A _0653_/B vssd1 vssd1 vccd1 vccd1 _0548_/A sky130_fd_sc_hd__and2_1
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0693__C1 _0680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_586 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0401_ _0821_/Q vssd1 vssd1 vccd1 vccd1 _0434_/A sky130_fd_sc_hd__clkbuf_2
Xpixel_macro_125 vssd1 vssd1 vccd1 vccd1 pixel_macro_125/HI io_oeb[35] sky130_fd_sc_hd__conb_1
Xpixel_macro_158 vssd1 vssd1 vccd1 vccd1 pixel_macro_158/HI io_out[30] sky130_fd_sc_hd__conb_1
Xpixel_macro_114 vssd1 vssd1 vccd1 vccd1 pixel_macro_114/HI io_oeb[24] sky130_fd_sc_hd__conb_1
Xpixel_macro_147 vssd1 vssd1 vccd1 vccd1 pixel_macro_147/HI io_out[19] sky130_fd_sc_hd__conb_1
Xpixel_macro_103 vssd1 vssd1 vccd1 vccd1 pixel_macro_103/HI io_oeb[13] sky130_fd_sc_hd__conb_1
Xpixel_macro_136 vssd1 vssd1 vccd1 vccd1 pixel_macro_136/HI io_out[8] sky130_fd_sc_hd__conb_1
XFILLER_23_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xpixel_macro_169 vssd1 vssd1 vccd1 vccd1 pixel_macro_169/HI la_data_out[4] sky130_fd_sc_hd__conb_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0881_ _0881_/D repeater64/X vssd1 vssd1 vccd1 vccd1 _0908_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0547__B _0653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput19 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0813__CLK _0839_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0864_ _0864_/D repeater65/X vssd1 vssd1 vccd1 vccd1 _0904_/Q sky130_fd_sc_hd__dlxtn_1
X_0795_ _0897_/Q _0764_/A _0794_/X _0731_/A vssd1 vssd1 vccd1 vccd1 _0839_/D sky130_fd_sc_hd__o211a_1
XANTENNA__0558__A _0566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0836__CLK _0838_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0580_ _0580_/A vssd1 vssd1 vccd1 vccd1 _0869_/D sky130_fd_sc_hd__clkbuf_1
X_0916_ _0916_/D _0417_/Y vssd1 vssd1 vccd1 vccd1 _0916_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA__0560__B _0560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0847_ _0847_/D _0452_/X vssd1 vssd1 vccd1 vccd1 _0911_/Q sky130_fd_sc_hd__dlxtn_1
X_0778_ _0832_/Q _0780_/B vssd1 vssd1 vccd1 vccd1 _0778_/X sky130_fd_sc_hd__or2_1
XFILLER_24_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0661__A _0661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0632_ _0640_/A _0632_/B vssd1 vssd1 vccd1 vccd1 _0633_/A sky130_fd_sc_hd__and2_1
X_0701_ input18/X _0689_/X _0698_/X _0700_/X vssd1 vssd1 vccd1 vccd1 _0803_/D sky130_fd_sc_hd__o211a_1
XFILLER_7_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0563_ _0563_/A vssd1 vssd1 vccd1 vccd1 _0872_/D sky130_fd_sc_hd__clkbuf_1
X_0494_ _0494_/A vssd1 vssd1 vccd1 vccd1 _0846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0571__A _0577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xpixel_macro_98 vssd1 vssd1 vccd1 vccd1 pixel_macro_98/HI io_oeb[8] sky130_fd_sc_hd__conb_1
XFILLER_25_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0656__A _0656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0615_ _0615_/A vssd1 vssd1 vccd1 vccd1 _0894_/D sky130_fd_sc_hd__clkbuf_1
X_0546_ _0546_/A vssd1 vssd1 vccd1 vccd1 _0853_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__0566__A _0566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0477_ _0920_/Q _0919_/Q _0476_/B vssd1 vssd1 vccd1 vccd1 _0477_/X sky130_fd_sc_hd__o21a_1
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0748__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_598 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0739__A1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0400_ _0433_/A _0400_/B vssd1 vssd1 vccd1 vccd1 _0514_/A sky130_fd_sc_hd__nand2_1
Xpixel_macro_104 vssd1 vssd1 vccd1 vccd1 pixel_macro_104/HI io_oeb[14] sky130_fd_sc_hd__conb_1
XFILLER_0_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_126 vssd1 vssd1 vccd1 vccd1 pixel_macro_126/HI io_oeb[36] sky130_fd_sc_hd__conb_1
Xpixel_macro_159 vssd1 vssd1 vccd1 vccd1 pixel_macro_159/HI io_out[31] sky130_fd_sc_hd__conb_1
Xpixel_macro_115 vssd1 vssd1 vccd1 vccd1 pixel_macro_115/HI io_oeb[25] sky130_fd_sc_hd__conb_1
Xpixel_macro_148 vssd1 vssd1 vccd1 vccd1 pixel_macro_148/HI io_out[20] sky130_fd_sc_hd__conb_1
Xpixel_macro_137 vssd1 vssd1 vccd1 vccd1 pixel_macro_137/HI io_out[9] sky130_fd_sc_hd__conb_1
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0529_ _0551_/A vssd1 vssd1 vccd1 vccd1 _0538_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0409__B1 _0918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0653__B _0653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0880_ _0880_/D repeater62/X vssd1 vssd1 vccd1 vccd1 _0907_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_23_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0664__A _0756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0863_ _0863_/D repeater85/X vssd1 vssd1 vccd1 vccd1 _0914_/Q sky130_fd_sc_hd__dlxtn_1
X_0794_ _0839_/Q _0794_/B vssd1 vssd1 vccd1 vccd1 _0794_/X sky130_fd_sc_hd__or2_1
XFILLER_3_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0749__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0659__A _0661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0915_ _0915_/D _0448_/X vssd1 vssd1 vccd1 vccd1 _0915_/Q sky130_fd_sc_hd__dlxtn_2
XANTENNA__0569__A _0577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0777_ _0777_/A vssd1 vssd1 vccd1 vccd1 _0777_/X sky130_fd_sc_hd__clkbuf_2
X_0846_ _0846_/D _0444_/A vssd1 vssd1 vccd1 vccd1 _0899_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_24_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0470__C _0470_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0803__CLK _0829_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0700_ _0731_/A vssd1 vssd1 vccd1 vccd1 _0700_/X sky130_fd_sc_hd__clkbuf_2
X_0562_ _0566_/A _0618_/B vssd1 vssd1 vccd1 vccd1 _0563_/A sky130_fd_sc_hd__and2_1
X_0631_ _1140_/A vssd1 vssd1 vccd1 vccd1 _0640_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0493_ _0500_/A _0618_/B vssd1 vssd1 vccd1 vccd1 _0494_/A sky130_fd_sc_hd__and2_1
XFILLER_21_202 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0829_ _0829_/CLK _0829_/D vssd1 vssd1 vccd1 vccd1 _0829_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0826__CLK _0839_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xpixel_macro_99 vssd1 vssd1 vccd1 vccd1 pixel_macro_99/HI io_oeb[9] sky130_fd_sc_hd__conb_1
XFILLER_25_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0614_ _0622_/A _0614_/B vssd1 vssd1 vccd1 vccd1 _0615_/A sky130_fd_sc_hd__and2_1
X_0545_ _0549_/A _0643_/B vssd1 vssd1 vccd1 vccd1 _0546_/A sky130_fd_sc_hd__and2_1
X_0476_ _0483_/A _0476_/B vssd1 vssd1 vccd1 vccd1 _0476_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0693__A1 _0678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_127 vssd1 vssd1 vccd1 vccd1 pixel_macro_127/HI io_oeb[37] sky130_fd_sc_hd__conb_1
Xpixel_macro_116 vssd1 vssd1 vccd1 vccd1 pixel_macro_116/HI io_oeb[26] sky130_fd_sc_hd__conb_1
Xpixel_macro_105 vssd1 vssd1 vccd1 vccd1 pixel_macro_105/HI io_oeb[15] sky130_fd_sc_hd__conb_1
Xpixel_macro_138 vssd1 vssd1 vccd1 vccd1 pixel_macro_138/HI io_out[10] sky130_fd_sc_hd__conb_1
Xpixel_macro_149 vssd1 vssd1 vccd1 vccd1 pixel_macro_149/HI io_out[21] sky130_fd_sc_hd__conb_1
XFILLER_16_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0577__A _0577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0528_ _0528_/A vssd1 vssd1 vccd1 vccd1 _0852_/D sky130_fd_sc_hd__clkbuf_1
X_0459_ _0929_/D vssd1 vssd1 vccd1 vccd1 _0926_/D sky130_fd_sc_hd__clkinv_2
XFILLER_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input11_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0409__A1 _0400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input3_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0931_ _0931_/D repeater84/X vssd1 vssd1 vccd1 vccd1 _0931_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0862_ _0862_/D repeater69/X vssd1 vssd1 vccd1 vccd1 _0913_/Q sky130_fd_sc_hd__dlxtn_1
X_0793_ _0904_/Q _0764_/A _0792_/X _0731_/A vssd1 vssd1 vccd1 vccd1 _0838_/D sky130_fd_sc_hd__o211a_1
XFILLER_9_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output42_A _0433_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0914_ _0914_/D _0439_/B vssd1 vssd1 vccd1 vccd1 _0914_/Q sky130_fd_sc_hd__dlxtn_1
X_0845_ _0845_/D repeater71/X vssd1 vssd1 vccd1 vccd1 _0910_/Q sky130_fd_sc_hd__dlxtn_1
X_0776_ _0908_/Q _0764_/X _0775_/X _0768_/X vssd1 vssd1 vccd1 vccd1 _0831_/D sky130_fd_sc_hd__o211a_1
XANTENNA__0585__A _0609_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0495__A _0510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0630_ _0630_/A vssd1 vssd1 vccd1 vccd1 _0915_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0492_ _0636_/B vssd1 vssd1 vccd1 vccd1 _0618_/B sky130_fd_sc_hd__clkbuf_1
X_0561_ _0561_/A vssd1 vssd1 vccd1 vccd1 _0870_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0759_ _0794_/B vssd1 vssd1 vccd1 vccd1 _0767_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_0828_ _0839_/CLK _0828_/D vssd1 vssd1 vccd1 vccd1 _0828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0920__CLK _0921_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0672__B _0758_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0613_ _1141_/A vssd1 vssd1 vccd1 vccd1 _0622_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0544_ _0544_/A vssd1 vssd1 vccd1 vccd1 _0860_/D sky130_fd_sc_hd__clkbuf_1
X_0475_ _0799_/Q vssd1 vssd1 vccd1 vccd1 _0475_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_22_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0773__A _0830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0436__A2 _0400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xpixel_macro_117 vssd1 vssd1 vccd1 vccd1 pixel_macro_117/HI io_oeb[27] sky130_fd_sc_hd__conb_1
Xpixel_macro_106 vssd1 vssd1 vccd1 vccd1 pixel_macro_106/HI io_oeb[16] sky130_fd_sc_hd__conb_1
Xpixel_macro_139 vssd1 vssd1 vccd1 vccd1 pixel_macro_139/HI io_out[11] sky130_fd_sc_hd__conb_1
Xpixel_macro_128 vssd1 vssd1 vccd1 vccd1 pixel_macro_128/HI io_out[0] sky130_fd_sc_hd__conb_1
XFILLER_16_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0816__CLK _0829_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0527_ _0930_/Q _0918_/D vssd1 vssd1 vccd1 vccd1 _0528_/A sky130_fd_sc_hd__and2_1
X_0458_ _0458_/A vssd1 vssd1 vccd1 vccd1 _0929_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_26_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0839__CLK _0839_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0678__A _0678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0419__A_N _0823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0861_ _0861_/D repeater66/X vssd1 vssd1 vccd1 vccd1 _0912_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_13_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0792_ _0838_/Q _0792_/B vssd1 vssd1 vccd1 vccd1 _0792_/X sky130_fd_sc_hd__or2_1
X_0930_ _0930_/D repeater83/X vssd1 vssd1 vccd1 vccd1 _0930_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_9_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output35_A _0525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0844_ _0844_/D repeater68/X vssd1 vssd1 vccd1 vccd1 _0897_/Q sky130_fd_sc_hd__dlxtn_1
X_0775_ _0831_/Q _0780_/B vssd1 vssd1 vccd1 vccd1 _0775_/X sky130_fd_sc_hd__or2_1
X_0913_ _0913_/D _0428_/A vssd1 vssd1 vccd1 vccd1 _0913_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0769__A1 _0917_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0491_ _0491_/A vssd1 vssd1 vccd1 vccd1 _0844_/D sky130_fd_sc_hd__clkbuf_1
X_0560_ _0566_/A _0560_/B vssd1 vssd1 vccd1 vccd1 _0561_/A sky130_fd_sc_hd__and2_1
XFILLER_19_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0758_ _0758_/A _0758_/B _0758_/C _0758_/D vssd1 vssd1 vccd1 vccd1 _0794_/B sky130_fd_sc_hd__and4_1
XFILLER_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0827_ _0839_/CLK _0827_/D vssd1 vssd1 vccd1 vccd1 _0827_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0596__A _0609_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0689_ _0704_/A vssd1 vssd1 vccd1 vccd1 _0689_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0612_ _0612_/A vssd1 vssd1 vccd1 vccd1 _0891_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0543_ _0549_/A _0622_/B vssd1 vssd1 vccd1 vccd1 _0544_/A sky130_fd_sc_hd__and2_1
X_0474_ _0474_/A vssd1 vssd1 vccd1 vccd1 _0474_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_118 vssd1 vssd1 vccd1 vccd1 pixel_macro_118/HI io_oeb[28] sky130_fd_sc_hd__conb_1
Xpixel_macro_107 vssd1 vssd1 vccd1 vccd1 pixel_macro_107/HI io_oeb[17] sky130_fd_sc_hd__conb_1
Xpixel_macro_129 vssd1 vssd1 vccd1 vccd1 pixel_macro_129/HI io_out[1] sky130_fd_sc_hd__conb_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0526_ _0526_/A vssd1 vssd1 vccd1 vccd1 _0849_/D sky130_fd_sc_hd__clkbuf_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0457_ _0483_/A _0483_/B vssd1 vssd1 vccd1 vccd1 _0458_/A sky130_fd_sc_hd__and2_1
XFILLER_25_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0741__C1 _0731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0509_ _0509_/A vssd1 vssd1 vccd1 vccd1 _0847_/D sky130_fd_sc_hd__clkbuf_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0806__CLK _0921_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0732__C1 _0731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0929__D _0929_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0860_ _0860_/D repeater70/X vssd1 vssd1 vccd1 vccd1 _0911_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_13_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0791_ _0899_/Q _0764_/A _0790_/X _0781_/X vssd1 vssd1 vccd1 vccd1 _0837_/D sky130_fd_sc_hd__o211a_1
XFILLER_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0599__A _0605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0829__CLK _0829_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_290 vssd1 vssd1 vccd1 vccd1 pixel_macro_290/HI wbs_dat_o[26] sky130_fd_sc_hd__conb_1
XFILLER_12_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output28_A _0820_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0912_ _0912_/D _0449_/B vssd1 vssd1 vccd1 vccd1 _0912_/Q sky130_fd_sc_hd__dlxtn_1
X_0774_ _0913_/Q _0764_/X _0773_/X _0768_/X vssd1 vssd1 vccd1 vccd1 _0830_/D sky130_fd_sc_hd__o211a_1
X_0843_ _0843_/D repeater87/X vssd1 vssd1 vccd1 vccd1 _0917_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0686__B _0758_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0490_ _0500_/A _0560_/B vssd1 vssd1 vccd1 vccd1 _0491_/A sky130_fd_sc_hd__and2_1
XFILLER_19_585 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0757_ input3/X input2/X input9/X input6/X vssd1 vssd1 vccd1 vccd1 _0758_/D sky130_fd_sc_hd__and4bb_1
X_0688_ _0705_/A _0736_/A vssd1 vssd1 vccd1 vccd1 _0704_/A sky130_fd_sc_hd__nand2_1
X_0826_ _0839_/CLK _0826_/D vssd1 vssd1 vccd1 vccd1 _0826_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0893__GATE_N _0436_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input27_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0611_ _0928_/Q _0918_/D vssd1 vssd1 vccd1 vccd1 _0612_/A sky130_fd_sc_hd__and2_1
X_0542_ _0542_/A vssd1 vssd1 vccd1 vccd1 _0855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0473_ _0809_/Q _0808_/Q _0473_/C _0473_/D vssd1 vssd1 vccd1 vccd1 _0474_/A sky130_fd_sc_hd__or4_2
XFILLER_22_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0809_ _0921_/CLK _0809_/D vssd1 vssd1 vccd1 vccd1 _0809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_119 vssd1 vssd1 vccd1 vccd1 pixel_macro_119/HI io_oeb[29] sky130_fd_sc_hd__conb_1
Xpixel_macro_108 vssd1 vssd1 vccd1 vccd1 pixel_macro_108/HI io_oeb[18] sky130_fd_sc_hd__conb_1
XANTENNA__1141__A _1141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0456_ _0466_/A _0476_/B vssd1 vssd1 vccd1 vccd1 _0483_/B sky130_fd_sc_hd__nor2_1
X_0525_ _0525_/A _0645_/B vssd1 vssd1 vccd1 vccd1 _0526_/A sky130_fd_sc_hd__and2_1
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput60 _0833_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
XANTENNA_output58_A _0831_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater80_A _0925_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0508_ _0519_/A _0622_/B vssd1 vssd1 vccd1 vccd1 _0509_/A sky130_fd_sc_hd__and2_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0439_ _0664_/B _0439_/B vssd1 vssd1 vccd1 vccd1 _0440_/A sky130_fd_sc_hd__or2_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_60 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0790_ _0837_/Q _0792_/B vssd1 vssd1 vccd1 vccd1 _0790_/X sky130_fd_sc_hd__or2_1
XFILLER_5_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input1_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xpixel_macro_291 vssd1 vssd1 vccd1 vccd1 pixel_macro_291/HI wbs_dat_o[27] sky130_fd_sc_hd__conb_1
Xpixel_macro_280 vssd1 vssd1 vccd1 vccd1 pixel_macro_280/HI wbs_dat_o[16] sky130_fd_sc_hd__conb_1
XFILLER_18_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0842_ _0842_/D repeater64/X vssd1 vssd1 vccd1 vccd1 _0908_/Q sky130_fd_sc_hd__dlxtn_1
X_0911_ _0911_/D repeater70/X vssd1 vssd1 vccd1 vccd1 _0911_/Q sky130_fd_sc_hd__dlxtn_1
X_0773_ _0830_/Q _0780_/B vssd1 vssd1 vccd1 vccd1 _0773_/X sky130_fd_sc_hd__or2_1
XFILLER_17_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output40_A _0483_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0819__CLK _0829_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0825_ _0838_/CLK _0825_/D vssd1 vssd1 vccd1 vccd1 _0825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0687_ _0706_/A vssd1 vssd1 vccd1 vccd1 _0736_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_0756_ _0756_/A _0756_/B _0756_/C vssd1 vssd1 vccd1 vccd1 _0756_/X sky130_fd_sc_hd__and3_1
XFILLER_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1139__A _1141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0541_ _0549_/A _0649_/B vssd1 vssd1 vccd1 vccd1 _0542_/A sky130_fd_sc_hd__and2_1
XFILLER_3_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0472_ _0807_/Q _0806_/Q _0805_/Q _0804_/Q vssd1 vssd1 vccd1 vccd1 _0473_/D sky130_fd_sc_hd__or4_1
XFILLER_7_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0610_ _0610_/A vssd1 vssd1 vccd1 vccd1 _0888_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0808_ _0921_/CLK _0808_/D vssd1 vssd1 vccd1 vccd1 _0808_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0400__B _0400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0739_ input20/X _0735_/X _0738_/X _0731_/X vssd1 vssd1 vccd1 vccd1 _0815_/D sky130_fd_sc_hd__o211a_1
XFILLER_4_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0798__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xpixel_macro_109 vssd1 vssd1 vccd1 vccd1 pixel_macro_109/HI io_oeb[19] sky130_fd_sc_hd__conb_1
XFILLER_0_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0455_ _0921_/Q vssd1 vssd1 vccd1 vccd1 _0476_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_0524_ _0655_/B vssd1 vssd1 vccd1 vccd1 _0645_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput50 _0837_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
Xoutput61 _0834_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0438_ _0438_/A _0503_/B vssd1 vssd1 vccd1 vccd1 _0441_/A sky130_fd_sc_hd__nand2_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0507_ _0640_/B vssd1 vssd1 vccd1 vccd1 _0622_/B sky130_fd_sc_hd__clkbuf_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0741__A1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0732__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_72 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_613 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater80 _0925_/Q vssd1 vssd1 vccd1 vccd1 _0406_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_15_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xpixel_macro_281 vssd1 vssd1 vccd1 vccd1 pixel_macro_281/HI wbs_dat_o[17] sky130_fd_sc_hd__conb_1
Xpixel_macro_292 vssd1 vssd1 vccd1 vccd1 pixel_macro_292/HI wbs_dat_o[28] sky130_fd_sc_hd__conb_1
Xpixel_macro_270 vssd1 vssd1 vccd1 vccd1 pixel_macro_270/HI la_data_out[119] sky130_fd_sc_hd__conb_1
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0841_ _0841_/D _0450_/X vssd1 vssd1 vccd1 vccd1 _0907_/Q sky130_fd_sc_hd__dlxtn_1
X_0772_ _0911_/Q _0764_/X _0771_/X _0768_/X vssd1 vssd1 vccd1 vccd1 _0829_/D sky130_fd_sc_hd__o211a_1
X_0910_ _0910_/D repeater71/X vssd1 vssd1 vccd1 vccd1 _0910_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_20_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output33_A _0609_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0824_ _0839_/CLK _0824_/D vssd1 vssd1 vccd1 vccd1 _0824_/Q sky130_fd_sc_hd__dfxtp_1
X_0755_ _0777_/A vssd1 vssd1 vccd1 vccd1 _0764_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0686_ _0758_/A _0758_/B _0686_/C _0758_/C vssd1 vssd1 vccd1 vccd1 _0706_/A sky130_fd_sc_hd__and4_1
XFILLER_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0540_ _0551_/A vssd1 vssd1 vccd1 vccd1 _0549_/A sky130_fd_sc_hd__clkbuf_2
X_0471_ _0803_/Q _0802_/Q _0801_/Q _0800_/Q vssd1 vssd1 vccd1 vccd1 _0473_/C sky130_fd_sc_hd__or4_1
XFILLER_19_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0738_ _0736_/X _0737_/X _0815_/Q vssd1 vssd1 vccd1 vccd1 _0738_/X sky130_fd_sc_hd__a21o_1
X_0807_ _0921_/CLK _0807_/D vssd1 vssd1 vccd1 vccd1 _0807_/Q sky130_fd_sc_hd__dfxtp_1
X_0669_ _0669_/A vssd1 vssd1 vccd1 vccd1 _0905_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_63 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0809__CLK _0921_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0454_ _0920_/Q vssd1 vssd1 vccd1 vccd1 _0466_/A sky130_fd_sc_hd__inv_2
X_0523_ _0523_/A vssd1 vssd1 vccd1 vccd1 _0843_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput40 _0483_/C vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
Xoutput51 _0838_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
XFILLER_16_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0512__A _0519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0506_ _0506_/A vssd1 vssd1 vccd1 vccd1 _0842_/D sky130_fd_sc_hd__clkbuf_1
XTAP_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0437_ _0514_/B _0495_/B vssd1 vssd1 vccd1 vccd1 _0664_/B sky130_fd_sc_hd__nor2_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0422__A _0821_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0717__C1 _0714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0708__C1 _0700_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater70 _0452_/X vssd1 vssd1 vccd1 vccd1 repeater70/X sky130_fd_sc_hd__clkbuf_1
Xrepeater81 _0417_/Y vssd1 vssd1 vccd1 vccd1 _0762_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_15_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xpixel_macro_260 vssd1 vssd1 vccd1 vccd1 pixel_macro_260/HI la_data_out[109] sky130_fd_sc_hd__conb_1
XFILLER_23_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0417__A _0756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xpixel_macro_282 vssd1 vssd1 vccd1 vccd1 pixel_macro_282/HI wbs_dat_o[18] sky130_fd_sc_hd__conb_1
Xpixel_macro_293 vssd1 vssd1 vccd1 vccd1 pixel_macro_293/HI wbs_dat_o[29] sky130_fd_sc_hd__conb_1
Xpixel_macro_271 vssd1 vssd1 vccd1 vccd1 pixel_macro_271/HI la_data_out[120] sky130_fd_sc_hd__conb_1
XFILLER_10_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_268 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0771_ _0829_/Q _0780_/B vssd1 vssd1 vccd1 vccd1 _0771_/X sky130_fd_sc_hd__or2_1
X_0840_ _0840_/D _0762_/A2 vssd1 vssd1 vccd1 vccd1 _0916_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_5_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0700__A _0731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0754_ _0754_/A _0754_/B _0754_/C _0758_/C vssd1 vssd1 vccd1 vccd1 _0777_/A sky130_fd_sc_hd__or4b_1
X_0685_ _0685_/A _0685_/B _0685_/C _0676_/B vssd1 vssd1 vccd1 vccd1 _0758_/C sky130_fd_sc_hd__nor4b_1
X_0823_ _0921_/CLK _0823_/D _0752_/Y vssd1 vssd1 vccd1 vccd1 _0823_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0926__GATE_N repeater82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_503 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0605__A _0605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0470_ _0819_/Q _0818_/Q _0470_/C _0470_/D vssd1 vssd1 vccd1 vccd1 _0483_/C sky130_fd_sc_hd__nor4_4
XFILLER_3_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0668_ _0756_/B _0668_/B vssd1 vssd1 vccd1 vccd1 _0669_/A sky130_fd_sc_hd__and2_1
X_0737_ _0737_/A vssd1 vssd1 vccd1 vccd1 _0737_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0806_ _0921_/CLK _0806_/D vssd1 vssd1 vccd1 vccd1 _0806_/Q sky130_fd_sc_hd__dfxtp_1
X_0599_ _0605_/A _0622_/B vssd1 vssd1 vccd1 vccd1 _0600_/A sky130_fd_sc_hd__and2_1
XFILLER_13_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input25_A wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0522_ _0930_/Q _0627_/B vssd1 vssd1 vccd1 vccd1 _0523_/A sky130_fd_sc_hd__and2_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0453_ _0919_/Q vssd1 vssd1 vccd1 vccd1 _0483_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput41 _0918_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
Xoutput30 _1141_/X vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
Xoutput52 _0839_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0505_ _0519_/A _0649_/B vssd1 vssd1 vccd1 vccd1 _0506_/A sky130_fd_sc_hd__and2_1
XTAP_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0436_ _0433_/A _0400_/B _0514_/B _0756_/C vssd1 vssd1 vccd1 vccd1 _0436_/Y sky130_fd_sc_hd__a31oi_4
.ends

