magic
tech sky130B
magscale 1 2
timestamp 1662149815
<< obsli1 >>
rect 1104 2159 38824 33745
<< obsm1 >>
rect 1104 2128 39178 33776
<< metal2 >>
rect 2870 35200 2926 36000
rect 8574 35200 8630 36000
rect 14278 35200 14334 36000
rect 19982 35200 20038 36000
rect 25686 35200 25742 36000
rect 31390 35200 31446 36000
rect 37094 35200 37150 36000
rect 846 0 902 800
rect 2042 0 2098 800
rect 3238 0 3294 800
rect 4434 0 4490 800
rect 5630 0 5686 800
rect 6826 0 6882 800
rect 8022 0 8078 800
rect 9218 0 9274 800
rect 10414 0 10470 800
rect 11610 0 11666 800
rect 12806 0 12862 800
rect 14002 0 14058 800
rect 15198 0 15254 800
rect 16394 0 16450 800
rect 17590 0 17646 800
rect 18786 0 18842 800
rect 19982 0 20038 800
rect 21178 0 21234 800
rect 22374 0 22430 800
rect 23570 0 23626 800
rect 24766 0 24822 800
rect 25962 0 26018 800
rect 27158 0 27214 800
rect 28354 0 28410 800
rect 29550 0 29606 800
rect 30746 0 30802 800
rect 31942 0 31998 800
rect 33138 0 33194 800
rect 34334 0 34390 800
rect 35530 0 35586 800
rect 36726 0 36782 800
rect 37922 0 37978 800
rect 39118 0 39174 800
<< obsm2 >>
rect 1398 35144 2814 35306
rect 2982 35144 8518 35306
rect 8686 35144 14222 35306
rect 14390 35144 19926 35306
rect 20094 35144 25630 35306
rect 25798 35144 31334 35306
rect 31502 35144 37038 35306
rect 37206 35144 39172 35306
rect 1398 856 39172 35144
rect 1398 734 1986 856
rect 2154 734 3182 856
rect 3350 734 4378 856
rect 4546 734 5574 856
rect 5742 734 6770 856
rect 6938 734 7966 856
rect 8134 734 9162 856
rect 9330 734 10358 856
rect 10526 734 11554 856
rect 11722 734 12750 856
rect 12918 734 13946 856
rect 14114 734 15142 856
rect 15310 734 16338 856
rect 16506 734 17534 856
rect 17702 734 18730 856
rect 18898 734 19926 856
rect 20094 734 21122 856
rect 21290 734 22318 856
rect 22486 734 23514 856
rect 23682 734 24710 856
rect 24878 734 25906 856
rect 26074 734 27102 856
rect 27270 734 28298 856
rect 28466 734 29494 856
rect 29662 734 30690 856
rect 30858 734 31886 856
rect 32054 734 33082 856
rect 33250 734 34278 856
rect 34446 734 35474 856
rect 35642 734 36670 856
rect 36838 734 37866 856
rect 38034 734 39062 856
<< metal3 >>
rect 0 34280 800 34400
rect 0 32920 800 33040
rect 0 31560 800 31680
rect 0 30200 800 30320
rect 0 28840 800 28960
rect 0 27480 800 27600
rect 0 26120 800 26240
rect 0 24760 800 24880
rect 0 23400 800 23520
rect 0 22040 800 22160
rect 0 20680 800 20800
rect 0 19320 800 19440
rect 0 17960 800 18080
rect 0 16600 800 16720
rect 0 15240 800 15360
rect 0 13880 800 14000
rect 0 12520 800 12640
rect 0 11160 800 11280
rect 0 9800 800 9920
rect 0 8440 800 8560
rect 0 7080 800 7200
rect 0 5720 800 5840
rect 0 4360 800 4480
rect 0 3000 800 3120
rect 0 1640 800 1760
<< obsm3 >>
rect 880 34200 34330 34373
rect 800 33120 34330 34200
rect 880 32840 34330 33120
rect 800 31760 34330 32840
rect 880 31480 34330 31760
rect 800 30400 34330 31480
rect 880 30120 34330 30400
rect 800 29040 34330 30120
rect 880 28760 34330 29040
rect 800 27680 34330 28760
rect 880 27400 34330 27680
rect 800 26320 34330 27400
rect 880 26040 34330 26320
rect 800 24960 34330 26040
rect 880 24680 34330 24960
rect 800 23600 34330 24680
rect 880 23320 34330 23600
rect 800 22240 34330 23320
rect 880 21960 34330 22240
rect 800 20880 34330 21960
rect 880 20600 34330 20880
rect 800 19520 34330 20600
rect 880 19240 34330 19520
rect 800 18160 34330 19240
rect 880 17880 34330 18160
rect 800 16800 34330 17880
rect 880 16520 34330 16800
rect 800 15440 34330 16520
rect 880 15160 34330 15440
rect 800 14080 34330 15160
rect 880 13800 34330 14080
rect 800 12720 34330 13800
rect 880 12440 34330 12720
rect 800 11360 34330 12440
rect 880 11080 34330 11360
rect 800 10000 34330 11080
rect 880 9720 34330 10000
rect 800 8640 34330 9720
rect 880 8360 34330 8640
rect 800 7280 34330 8360
rect 880 7000 34330 7280
rect 800 5920 34330 7000
rect 880 5640 34330 5920
rect 800 4560 34330 5640
rect 880 4280 34330 4560
rect 800 3200 34330 4280
rect 880 2920 34330 3200
rect 800 1840 34330 2920
rect 880 1667 34330 1840
<< metal4 >>
rect 5668 2128 5988 33776
rect 10392 2128 10712 33776
rect 15116 2128 15436 33776
rect 19840 2128 20160 33776
rect 24564 2128 24884 33776
rect 29288 2128 29608 33776
rect 34012 2128 34332 33776
<< labels >>
rlabel metal2 s 28354 0 28410 800 6 adj_max_clk[0]
port 1 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 adj_max_clk[1]
port 2 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 adj_max_clk[2]
port 3 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 adj_max_clk[3]
port 4 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 adj_max_clk[4]
port 5 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 adj_max_clk[5]
port 6 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 adj_max_clk[6]
port 7 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 adj_max_clk[7]
port 8 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 adj_max_clk[8]
port 9 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 adj_max_clk[9]
port 10 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 adj_timer_en
port 11 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 adj_timer_m_i
port 12 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 adj_timer_max
port 13 nsew signal output
rlabel metal2 s 2870 35200 2926 36000 6 clk
port 14 nsew signal input
rlabel metal2 s 14278 35200 14334 36000 6 data_in
port 15 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 data_out[0]
port 16 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 data_out[10]
port 17 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 data_out[11]
port 18 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 data_out[12]
port 19 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 data_out[13]
port 20 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 data_out[14]
port 21 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 data_out[15]
port 22 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 data_out[1]
port 23 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 data_out[2]
port 24 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 data_out[3]
port 25 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 data_out[4]
port 26 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 data_out[5]
port 27 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 data_out[6]
port 28 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 data_out[7]
port 29 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 data_out[8]
port 30 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 data_out[9]
port 31 nsew signal output
rlabel metal2 s 19982 35200 20038 36000 6 data_sel[0]
port 32 nsew signal output
rlabel metal2 s 25686 35200 25742 36000 6 data_sel[1]
port 33 nsew signal output
rlabel metal2 s 31390 35200 31446 36000 6 data_sel[2]
port 34 nsew signal output
rlabel metal2 s 37094 35200 37150 36000 6 data_sel[3]
port 35 nsew signal output
rlabel metal3 s 0 34280 800 34400 6 kernel_done_o
port 36 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 loc_max_clk[0]
port 37 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 loc_max_clk[1]
port 38 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 loc_max_clk[2]
port 39 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 loc_max_clk[3]
port 40 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 loc_max_clk[4]
port 41 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 loc_max_clk[5]
port 42 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 loc_max_clk[6]
port 43 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 loc_max_clk[7]
port 44 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 loc_max_clk[8]
port 45 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 loc_max_clk[9]
port 46 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 loc_timer_en
port 47 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 loc_timer_m_i
port 48 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 loc_timer_max
port 49 nsew signal output
rlabel metal2 s 846 0 902 800 6 pxl_done_i
port 50 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 pxl_done_o
port 51 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 pxl_q[0]
port 52 nsew signal output
rlabel metal2 s 5630 0 5686 800 6 pxl_q[1]
port 53 nsew signal output
rlabel metal2 s 6826 0 6882 800 6 pxl_q[2]
port 54 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 pxl_q[3]
port 55 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 pxl_start_i
port 56 nsew signal input
rlabel metal2 s 8574 35200 8630 36000 6 reset
port 57 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 s1
port 58 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 s1_inv
port 59 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 s2
port 60 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 s2_inv
port 61 nsew signal output
rlabel metal3 s 0 28840 800 28960 6 s_p1
port 62 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 s_p2
port 63 nsew signal output
rlabel metal3 s 0 31560 800 31680 6 v_b0
port 64 nsew signal output
rlabel metal3 s 0 32920 800 33040 6 v_b1
port 65 nsew signal output
rlabel metal4 s 5668 2128 5988 33776 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 15116 2128 15436 33776 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 24564 2128 24884 33776 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 34012 2128 34332 33776 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 10392 2128 10712 33776 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 19840 2128 20160 33776 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 29288 2128 29608 33776 6 vssd1
port 67 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 36000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1681916
string GDS_FILE /home/mxmont/Documents/Universidad/IC-UBB/MixPix/CARAVEL_WRAPPER/MixPix/openlane/pixel/runs/22_09_02_16_15/results/signoff/pixel.magic.gds
string GDS_START 322244
<< end >>

