magic
tech sky130A
magscale 1 2
timestamp 1669402136
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 410518 700476 410524 700528
rect 410576 700516 410582 700528
rect 429838 700516 429844 700528
rect 410576 700488 429844 700516
rect 410576 700476 410582 700488
rect 429838 700476 429844 700488
rect 429896 700476 429902 700528
rect 399478 700408 399484 700460
rect 399536 700448 399542 700460
rect 446122 700448 446128 700460
rect 399536 700420 446128 700448
rect 399536 700408 399542 700420
rect 446122 700408 446128 700420
rect 446180 700408 446186 700460
rect 409138 700340 409144 700392
rect 409196 700380 409202 700392
rect 494790 700380 494796 700392
rect 409196 700352 494796 700380
rect 409196 700340 409202 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 33778 700312 33784 700324
rect 24360 700284 33784 700312
rect 24360 700272 24366 700284
rect 33778 700272 33784 700284
rect 33836 700272 33842 700324
rect 407758 700272 407764 700324
rect 407816 700312 407822 700324
rect 559650 700312 559656 700324
rect 407816 700284 559656 700312
rect 407816 700272 407822 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 196618 699660 196624 699712
rect 196676 699700 196682 699712
rect 202782 699700 202788 699712
rect 196676 699672 202788 699700
rect 196676 699660 196682 699672
rect 202782 699660 202788 699672
rect 202840 699660 202846 699712
rect 229738 699660 229744 699712
rect 229796 699700 229802 699712
rect 235166 699700 235172 699712
rect 229796 699672 235172 699700
rect 229796 699660 229802 699672
rect 235166 699660 235172 699672
rect 235224 699660 235230 699712
rect 364978 699660 364984 699712
rect 365036 699700 365042 699712
rect 369118 699700 369124 699712
rect 365036 699672 369124 699700
rect 365036 699660 365042 699672
rect 369118 699660 369124 699672
rect 369176 699660 369182 699712
rect 300118 697688 300124 697740
rect 300176 697728 300182 697740
rect 307018 697728 307024 697740
rect 300176 697700 307024 697728
rect 300176 697688 300182 697700
rect 307018 697688 307024 697700
rect 307076 697688 307082 697740
rect 260098 697280 260104 697332
rect 260156 697320 260162 697332
rect 267642 697320 267648 697332
rect 260156 697292 267648 697320
rect 260156 697280 260162 697292
rect 267642 697280 267648 697292
rect 267700 697280 267706 697332
rect 152826 696940 152832 696992
rect 152884 696980 152890 696992
rect 154114 696980 154120 696992
rect 152884 696952 154120 696980
rect 152884 696940 152890 696952
rect 154114 696940 154120 696952
rect 154172 696940 154178 696992
rect 504358 696940 504364 696992
rect 504416 696980 504422 696992
rect 580166 696980 580172 696992
rect 504416 696952 580172 696980
rect 504416 696940 504422 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 150434 692792 150440 692844
rect 150492 692832 150498 692844
rect 152826 692832 152832 692844
rect 150492 692804 152832 692832
rect 150492 692792 150498 692804
rect 152826 692792 152832 692804
rect 152884 692792 152890 692844
rect 185578 692044 185584 692096
rect 185636 692084 185642 692096
rect 196618 692084 196624 692096
rect 185636 692056 196624 692084
rect 185636 692044 185642 692056
rect 196618 692044 196624 692056
rect 196676 692044 196682 692096
rect 210418 690616 210424 690668
rect 210476 690656 210482 690668
rect 229738 690656 229744 690668
rect 210476 690628 229744 690656
rect 210476 690616 210482 690628
rect 229738 690616 229744 690628
rect 229796 690616 229802 690668
rect 180058 689256 180064 689308
rect 180116 689296 180122 689308
rect 185578 689296 185584 689308
rect 180116 689268 185584 689296
rect 180116 689256 180122 689268
rect 185578 689256 185584 689268
rect 185636 689256 185642 689308
rect 369118 688576 369124 688628
rect 369176 688616 369182 688628
rect 374638 688616 374644 688628
rect 369176 688588 374644 688616
rect 369176 688576 369182 688588
rect 374638 688576 374644 688588
rect 374696 688576 374702 688628
rect 347774 688440 347780 688492
rect 347832 688480 347838 688492
rect 351914 688480 351920 688492
rect 347832 688452 351920 688480
rect 347832 688440 347838 688452
rect 351914 688440 351920 688452
rect 351972 688440 351978 688492
rect 150342 687256 150348 687268
rect 147692 687228 150348 687256
rect 146938 687148 146944 687200
rect 146996 687188 147002 687200
rect 147692 687188 147720 687228
rect 150342 687216 150348 687228
rect 150400 687216 150406 687268
rect 146996 687160 147720 687188
rect 146996 687148 147002 687160
rect 307018 684428 307024 684480
rect 307076 684468 307082 684480
rect 310238 684468 310244 684480
rect 307076 684440 310244 684468
rect 307076 684428 307082 684440
rect 310238 684428 310244 684440
rect 310296 684428 310302 684480
rect 351914 683748 351920 683800
rect 351972 683788 351978 683800
rect 362218 683788 362224 683800
rect 351972 683760 362224 683788
rect 351972 683748 351978 683760
rect 362218 683748 362224 683760
rect 362276 683748 362282 683800
rect 374638 682252 374644 682304
rect 374696 682292 374702 682304
rect 380250 682292 380256 682304
rect 374696 682264 380256 682292
rect 374696 682252 374702 682264
rect 380250 682252 380256 682264
rect 380308 682252 380314 682304
rect 362218 680960 362224 681012
rect 362276 681000 362282 681012
rect 371234 681000 371240 681012
rect 362276 680972 371240 681000
rect 362276 680960 362282 680972
rect 371234 680960 371240 680972
rect 371292 680960 371298 681012
rect 217318 680348 217324 680400
rect 217376 680388 217382 680400
rect 218054 680388 218060 680400
rect 217376 680360 218060 680388
rect 217376 680348 217382 680360
rect 218054 680348 218060 680360
rect 218112 680348 218118 680400
rect 310238 678716 310244 678768
rect 310296 678756 310302 678768
rect 315298 678756 315304 678768
rect 310296 678728 315304 678756
rect 310296 678716 310302 678728
rect 315298 678716 315304 678728
rect 315356 678716 315362 678768
rect 253566 678444 253572 678496
rect 253624 678484 253630 678496
rect 260098 678484 260104 678496
rect 253624 678456 260104 678484
rect 253624 678444 253630 678456
rect 260098 678444 260104 678456
rect 260156 678444 260162 678496
rect 144914 678240 144920 678292
rect 144972 678280 144978 678292
rect 146938 678280 146944 678292
rect 144972 678252 146944 678280
rect 144972 678240 144978 678252
rect 146938 678240 146944 678252
rect 146996 678240 147002 678292
rect 135990 676812 135996 676864
rect 136048 676852 136054 676864
rect 144914 676852 144920 676864
rect 136048 676824 144920 676852
rect 136048 676812 136054 676824
rect 144914 676812 144920 676824
rect 144972 676812 144978 676864
rect 371234 675452 371240 675504
rect 371292 675492 371298 675504
rect 380158 675492 380164 675504
rect 371292 675464 380164 675492
rect 371292 675452 371298 675464
rect 380158 675452 380164 675464
rect 380216 675452 380222 675504
rect 380250 675452 380256 675504
rect 380308 675492 380314 675504
rect 396442 675492 396448 675504
rect 380308 675464 396448 675492
rect 380308 675452 380314 675464
rect 396442 675452 396448 675464
rect 396500 675452 396506 675504
rect 278406 674772 278412 674824
rect 278464 674812 278470 674824
rect 282822 674812 282828 674824
rect 278464 674784 282828 674812
rect 278464 674772 278470 674784
rect 282822 674772 282828 674784
rect 282880 674772 282886 674824
rect 331214 674772 331220 674824
rect 331272 674812 331278 674824
rect 334618 674812 334624 674824
rect 331272 674784 334624 674812
rect 331272 674772 331278 674784
rect 334618 674772 334624 674784
rect 334676 674772 334682 674824
rect 133874 674432 133880 674484
rect 133932 674472 133938 674484
rect 135990 674472 135996 674484
rect 133932 674444 135996 674472
rect 133932 674432 133938 674444
rect 135990 674432 135996 674444
rect 136048 674432 136054 674484
rect 250438 674024 250444 674076
rect 250496 674064 250502 674076
rect 253566 674064 253572 674076
rect 250496 674036 253572 674064
rect 250496 674024 250502 674036
rect 253566 674024 253572 674036
rect 253624 674024 253630 674076
rect 2774 670692 2780 670744
rect 2832 670732 2838 670744
rect 6178 670732 6184 670744
rect 2832 670704 6184 670732
rect 2832 670692 2838 670704
rect 6178 670692 6184 670704
rect 6236 670692 6242 670744
rect 544378 670692 544384 670744
rect 544436 670732 544442 670744
rect 580166 670732 580172 670744
rect 544436 670704 580172 670732
rect 544436 670692 544442 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 276658 669060 276664 669112
rect 276716 669100 276722 669112
rect 278406 669100 278412 669112
rect 276716 669072 278412 669100
rect 276716 669060 276722 669072
rect 278406 669060 278412 669072
rect 278464 669060 278470 669112
rect 131758 667496 131764 667548
rect 131816 667536 131822 667548
rect 133874 667536 133880 667548
rect 131816 667508 133880 667536
rect 131816 667496 131822 667508
rect 133874 667496 133880 667508
rect 133932 667496 133938 667548
rect 202138 667156 202144 667208
rect 202196 667196 202202 667208
rect 210418 667196 210424 667208
rect 202196 667168 210424 667196
rect 202196 667156 202202 667168
rect 210418 667156 210424 667168
rect 210476 667156 210482 667208
rect 177298 666408 177304 666460
rect 177356 666448 177362 666460
rect 180058 666448 180064 666460
rect 177356 666420 180064 666448
rect 177356 666408 177362 666420
rect 180058 666408 180064 666420
rect 180116 666408 180122 666460
rect 247678 663756 247684 663808
rect 247736 663796 247742 663808
rect 250438 663796 250444 663808
rect 247736 663768 250444 663796
rect 247736 663756 247742 663768
rect 250438 663756 250444 663768
rect 250496 663756 250502 663808
rect 334618 663008 334624 663060
rect 334676 663048 334682 663060
rect 358078 663048 358084 663060
rect 334676 663020 358084 663048
rect 334676 663008 334682 663020
rect 358078 663008 358084 663020
rect 358136 663008 358142 663060
rect 127618 662396 127624 662448
rect 127676 662436 127682 662448
rect 131758 662436 131764 662448
rect 127676 662408 131764 662436
rect 127676 662396 127682 662408
rect 131758 662396 131764 662408
rect 131816 662396 131822 662448
rect 174538 662396 174544 662448
rect 174596 662436 174602 662448
rect 177298 662436 177304 662448
rect 174596 662408 177304 662436
rect 174596 662396 174602 662408
rect 177298 662396 177304 662408
rect 177356 662396 177362 662448
rect 273898 661036 273904 661088
rect 273956 661076 273962 661088
rect 276658 661076 276664 661088
rect 273956 661048 276664 661076
rect 273956 661036 273962 661048
rect 276658 661036 276664 661048
rect 276716 661036 276722 661088
rect 214558 658792 214564 658844
rect 214616 658832 214622 658844
rect 217318 658832 217324 658844
rect 214616 658804 217324 658832
rect 214616 658792 214622 658804
rect 217318 658792 217324 658804
rect 217376 658792 217382 658844
rect 315298 653352 315304 653404
rect 315356 653392 315362 653404
rect 319806 653392 319812 653404
rect 315356 653364 319812 653392
rect 315356 653352 315362 653364
rect 319806 653352 319812 653364
rect 319864 653352 319870 653404
rect 171686 651380 171692 651432
rect 171744 651420 171750 651432
rect 174538 651420 174544 651432
rect 171744 651392 174544 651420
rect 171744 651380 171750 651392
rect 174538 651380 174544 651392
rect 174596 651380 174602 651432
rect 195238 650700 195244 650752
rect 195296 650740 195302 650752
rect 202138 650740 202144 650752
rect 195296 650712 202144 650740
rect 195296 650700 195302 650712
rect 202138 650700 202144 650712
rect 202196 650700 202202 650752
rect 273898 650060 273904 650072
rect 270788 650032 273904 650060
rect 269758 649952 269764 650004
rect 269816 649992 269822 650004
rect 270788 649992 270816 650032
rect 273898 650020 273904 650032
rect 273956 650020 273962 650072
rect 269816 649964 270816 649992
rect 269816 649952 269822 649964
rect 358078 649952 358084 650004
rect 358136 649992 358142 650004
rect 366358 649992 366364 650004
rect 358136 649964 366364 649992
rect 358136 649952 358142 649964
rect 366358 649952 366364 649964
rect 366416 649952 366422 650004
rect 163498 649272 163504 649324
rect 163556 649312 163562 649324
rect 171686 649312 171692 649324
rect 163556 649284 171692 649312
rect 163556 649272 163562 649284
rect 171686 649272 171692 649284
rect 171744 649272 171750 649324
rect 380158 649272 380164 649324
rect 380216 649312 380222 649324
rect 387058 649312 387064 649324
rect 380216 649284 387064 649312
rect 380216 649272 380222 649284
rect 387058 649272 387064 649284
rect 387116 649272 387122 649324
rect 319806 648864 319812 648916
rect 319864 648904 319870 648916
rect 324958 648904 324964 648916
rect 319864 648876 324964 648904
rect 319864 648864 319870 648876
rect 324958 648864 324964 648876
rect 325016 648864 325022 648916
rect 127618 648632 127624 648644
rect 125612 648604 127624 648632
rect 124858 648524 124864 648576
rect 124916 648564 124922 648576
rect 125612 648564 125640 648604
rect 127618 648592 127624 648604
rect 127676 648592 127682 648644
rect 124916 648536 125640 648564
rect 124916 648524 124922 648536
rect 265618 647912 265624 647964
rect 265676 647952 265682 647964
rect 269758 647952 269764 647964
rect 265676 647924 269764 647952
rect 265676 647912 265682 647924
rect 269758 647912 269764 647924
rect 269816 647912 269822 647964
rect 366358 647164 366364 647216
rect 366416 647204 366422 647216
rect 371878 647204 371884 647216
rect 366416 647176 371884 647204
rect 366416 647164 366422 647176
rect 371878 647164 371884 647176
rect 371936 647164 371942 647216
rect 244918 645804 244924 645856
rect 244976 645844 244982 645856
rect 247678 645844 247684 645856
rect 244976 645816 247684 645844
rect 244976 645804 244982 645816
rect 247678 645804 247684 645816
rect 247736 645804 247742 645856
rect 324958 640228 324964 640280
rect 325016 640268 325022 640280
rect 327718 640268 327724 640280
rect 325016 640240 327724 640268
rect 325016 640228 325022 640240
rect 327718 640228 327724 640240
rect 327776 640228 327782 640280
rect 156598 638460 156604 638512
rect 156656 638500 156662 638512
rect 163498 638500 163504 638512
rect 156656 638472 163504 638500
rect 156656 638460 156662 638472
rect 163498 638460 163504 638472
rect 163556 638460 163562 638512
rect 371878 635468 371884 635520
rect 371936 635508 371942 635520
rect 388898 635508 388904 635520
rect 371936 635480 388904 635508
rect 371936 635468 371942 635480
rect 388898 635468 388904 635480
rect 388956 635468 388962 635520
rect 327718 632476 327724 632528
rect 327776 632516 327782 632528
rect 329926 632516 329932 632528
rect 327776 632488 329932 632516
rect 327776 632476 327782 632488
rect 329926 632476 329932 632488
rect 329984 632476 329990 632528
rect 388898 631660 388904 631712
rect 388956 631700 388962 631712
rect 395338 631700 395344 631712
rect 388956 631672 395344 631700
rect 388956 631660 388962 631672
rect 395338 631660 395344 631672
rect 395396 631660 395402 631712
rect 329926 629892 329932 629944
rect 329984 629932 329990 629944
rect 339494 629932 339500 629944
rect 329984 629904 339500 629932
rect 329984 629892 329990 629904
rect 339494 629892 339500 629904
rect 339552 629892 339558 629944
rect 339494 626492 339500 626544
rect 339552 626532 339558 626544
rect 344002 626532 344008 626544
rect 339552 626504 344008 626532
rect 339552 626492 339558 626504
rect 344002 626492 344008 626504
rect 344060 626492 344066 626544
rect 186958 623024 186964 623076
rect 187016 623064 187022 623076
rect 195238 623064 195244 623076
rect 187016 623036 195244 623064
rect 187016 623024 187022 623036
rect 195238 623024 195244 623036
rect 195296 623024 195302 623076
rect 152458 622412 152464 622464
rect 152516 622452 152522 622464
rect 156598 622452 156604 622464
rect 152516 622424 156604 622452
rect 152516 622412 152522 622424
rect 156598 622412 156604 622424
rect 156656 622412 156662 622464
rect 344002 620236 344008 620288
rect 344060 620276 344066 620288
rect 353294 620276 353300 620288
rect 344060 620248 353300 620276
rect 344060 620236 344066 620248
rect 353294 620236 353300 620248
rect 353352 620236 353358 620288
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 15838 618304 15844 618316
rect 3568 618276 15844 618304
rect 3568 618264 3574 618276
rect 15838 618264 15844 618276
rect 15896 618264 15902 618316
rect 353294 617516 353300 617568
rect 353352 617556 353358 617568
rect 395430 617556 395436 617568
rect 353352 617528 395436 617556
rect 353352 617516 353358 617528
rect 395430 617516 395436 617528
rect 395488 617516 395494 617568
rect 406378 616836 406384 616888
rect 406436 616876 406442 616888
rect 579706 616876 579712 616888
rect 406436 616848 579712 616876
rect 406436 616836 406442 616848
rect 579706 616836 579712 616848
rect 579764 616836 579770 616888
rect 184198 612756 184204 612808
rect 184256 612796 184262 612808
rect 186958 612796 186964 612808
rect 184256 612768 186964 612796
rect 184256 612756 184262 612768
rect 186958 612756 186964 612768
rect 187016 612756 187022 612808
rect 211798 609696 211804 609748
rect 211856 609736 211862 609748
rect 214558 609736 214564 609748
rect 211856 609708 214564 609736
rect 211856 609696 211862 609708
rect 214558 609696 214564 609708
rect 214616 609696 214622 609748
rect 138658 603712 138664 603764
rect 138716 603752 138722 603764
rect 152458 603752 152464 603764
rect 138716 603724 152464 603752
rect 138716 603712 138722 603724
rect 152458 603712 152464 603724
rect 152516 603712 152522 603764
rect 178034 603712 178040 603764
rect 178092 603752 178098 603764
rect 184198 603752 184204 603764
rect 178092 603724 184204 603752
rect 178092 603712 178098 603724
rect 184198 603712 184204 603724
rect 184256 603712 184262 603764
rect 124858 603140 124864 603152
rect 122806 603112 124864 603140
rect 121454 603032 121460 603084
rect 121512 603072 121518 603084
rect 122806 603072 122834 603112
rect 124858 603100 124864 603112
rect 124916 603100 124922 603152
rect 121512 603044 122834 603072
rect 121512 603032 121518 603044
rect 171778 600312 171784 600364
rect 171836 600352 171842 600364
rect 178034 600352 178040 600364
rect 171836 600324 178040 600352
rect 171836 600312 171842 600324
rect 178034 600312 178040 600324
rect 178092 600312 178098 600364
rect 119982 599564 119988 599616
rect 120040 599604 120046 599616
rect 121454 599604 121460 599616
rect 120040 599576 121460 599604
rect 120040 599564 120046 599576
rect 121454 599564 121460 599576
rect 121512 599564 121518 599616
rect 263594 598748 263600 598800
rect 263652 598788 263658 598800
rect 265618 598788 265624 598800
rect 263652 598760 265624 598788
rect 263652 598748 263658 598760
rect 265618 598748 265624 598760
rect 265676 598748 265682 598800
rect 117682 597184 117688 597236
rect 117740 597224 117746 597236
rect 119982 597224 119988 597236
rect 117740 597196 119988 597224
rect 117740 597184 117746 597196
rect 119982 597184 119988 597196
rect 120040 597184 120046 597236
rect 249058 595416 249064 595468
rect 249116 595456 249122 595468
rect 263594 595456 263600 595468
rect 249116 595428 263600 595456
rect 249116 595416 249122 595428
rect 263594 595416 263600 595428
rect 263652 595416 263658 595468
rect 210418 592016 210424 592068
rect 210476 592056 210482 592068
rect 211798 592056 211804 592068
rect 210476 592028 211804 592056
rect 210476 592016 210482 592028
rect 211798 592016 211804 592028
rect 211856 592016 211862 592068
rect 115198 590588 115204 590640
rect 115256 590628 115262 590640
rect 117682 590628 117688 590640
rect 115256 590600 117688 590628
rect 115256 590588 115262 590600
rect 117682 590588 117688 590600
rect 117740 590588 117746 590640
rect 241606 581136 241612 581188
rect 241664 581176 241670 581188
rect 244918 581176 244924 581188
rect 241664 581148 244924 581176
rect 241664 581136 241670 581148
rect 244918 581136 244924 581148
rect 244976 581136 244982 581188
rect 112438 580932 112444 580984
rect 112496 580972 112502 580984
rect 115198 580972 115204 580984
rect 112496 580944 115204 580972
rect 112496 580932 112502 580944
rect 115198 580932 115204 580944
rect 115256 580932 115262 580984
rect 135898 580660 135904 580712
rect 135956 580700 135962 580712
rect 138658 580700 138664 580712
rect 135956 580672 138664 580700
rect 135956 580660 135962 580672
rect 138658 580660 138664 580672
rect 138716 580660 138722 580712
rect 157978 580252 157984 580304
rect 158036 580292 158042 580304
rect 171778 580292 171784 580304
rect 158036 580264 171784 580292
rect 158036 580252 158042 580264
rect 171778 580252 171784 580264
rect 171836 580252 171842 580304
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 19978 579680 19984 579692
rect 3384 579652 19984 579680
rect 3384 579640 3390 579652
rect 19978 579640 19984 579652
rect 20036 579640 20042 579692
rect 238754 577600 238760 577652
rect 238812 577640 238818 577652
rect 241606 577640 241612 577652
rect 238812 577612 241612 577640
rect 238812 577600 238818 577612
rect 241606 577600 241612 577612
rect 241664 577600 241670 577652
rect 236638 574064 236644 574116
rect 236696 574104 236702 574116
rect 238754 574104 238760 574116
rect 236696 574076 238760 574104
rect 236696 574064 236702 574076
rect 238754 574064 238760 574076
rect 238812 574064 238818 574116
rect 126238 571956 126244 572008
rect 126296 571996 126302 572008
rect 135898 571996 135904 572008
rect 126296 571968 135904 571996
rect 126296 571956 126302 571968
rect 135898 571956 135904 571968
rect 135956 571956 135962 572008
rect 3050 565836 3056 565888
rect 3108 565876 3114 565888
rect 43438 565876 43444 565888
rect 3108 565848 43444 565876
rect 3108 565836 3114 565848
rect 43438 565836 43444 565848
rect 43496 565836 43502 565888
rect 404998 563048 405004 563100
rect 405056 563088 405062 563100
rect 580166 563088 580172 563100
rect 405056 563060 580172 563088
rect 405056 563048 405062 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 233234 562096 233240 562148
rect 233292 562136 233298 562148
rect 236638 562136 236644 562148
rect 233292 562108 236644 562136
rect 233292 562096 233298 562108
rect 236638 562096 236644 562108
rect 236696 562096 236702 562148
rect 209038 558152 209044 558204
rect 209096 558192 209102 558204
rect 233234 558192 233240 558204
rect 209096 558164 233240 558192
rect 209096 558152 209102 558164
rect 233234 558152 233240 558164
rect 233292 558152 233298 558204
rect 207658 554412 207664 554464
rect 207716 554452 207722 554464
rect 210418 554452 210424 554464
rect 207716 554424 210424 554452
rect 207716 554412 207722 554424
rect 210418 554412 210424 554424
rect 210476 554412 210482 554464
rect 149698 545708 149704 545760
rect 149756 545748 149762 545760
rect 157978 545748 157984 545760
rect 149756 545720 157984 545748
rect 149756 545708 149762 545720
rect 157978 545708 157984 545720
rect 158036 545708 158042 545760
rect 206278 543736 206284 543788
rect 206336 543776 206342 543788
rect 207658 543776 207664 543788
rect 206336 543748 207664 543776
rect 206336 543736 206342 543748
rect 207658 543736 207664 543748
rect 207716 543736 207722 543788
rect 204898 536800 204904 536852
rect 204956 536840 204962 536852
rect 209038 536840 209044 536852
rect 204956 536812 209044 536840
rect 204956 536800 204962 536812
rect 209038 536800 209044 536812
rect 209096 536800 209102 536852
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 20070 527184 20076 527196
rect 3016 527156 20076 527184
rect 3016 527144 3022 527156
rect 20070 527144 20076 527156
rect 20128 527144 20134 527196
rect 112438 525824 112444 525836
rect 109696 525796 112444 525824
rect 108942 525716 108948 525768
rect 109000 525756 109006 525768
rect 109696 525756 109724 525796
rect 112438 525784 112444 525796
rect 112496 525784 112502 525836
rect 123478 525784 123484 525836
rect 123536 525824 123542 525836
rect 126238 525824 126244 525836
rect 123536 525796 126244 525824
rect 123536 525784 123542 525796
rect 126238 525784 126244 525796
rect 126296 525784 126302 525836
rect 109000 525728 109724 525756
rect 109000 525716 109006 525728
rect 106918 522520 106924 522572
rect 106976 522560 106982 522572
rect 108942 522560 108948 522572
rect 106976 522532 108948 522560
rect 106976 522520 106982 522532
rect 108942 522520 108948 522532
rect 109000 522520 109006 522572
rect 2774 514768 2780 514820
rect 2832 514808 2838 514820
rect 4798 514808 4804 514820
rect 2832 514780 4804 514808
rect 2832 514768 2838 514780
rect 4798 514768 4804 514780
rect 4856 514768 4862 514820
rect 105538 514768 105544 514820
rect 105596 514808 105602 514820
rect 106918 514808 106924 514820
rect 105596 514780 106924 514808
rect 105596 514768 105602 514780
rect 106918 514768 106924 514780
rect 106976 514768 106982 514820
rect 115198 514020 115204 514072
rect 115256 514060 115262 514072
rect 123478 514060 123484 514072
rect 115256 514032 123484 514060
rect 115256 514020 115262 514032
rect 123478 514020 123484 514032
rect 123536 514020 123542 514072
rect 203518 511912 203524 511964
rect 203576 511952 203582 511964
rect 206278 511952 206284 511964
rect 203576 511924 206284 511952
rect 203576 511912 203582 511924
rect 206278 511912 206284 511924
rect 206336 511912 206342 511964
rect 403618 510620 403624 510672
rect 403676 510660 403682 510672
rect 580166 510660 580172 510672
rect 403676 510632 580172 510660
rect 403676 510620 403682 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 201862 507832 201868 507884
rect 201920 507872 201926 507884
rect 204898 507872 204904 507884
rect 201920 507844 204904 507872
rect 201920 507832 201926 507844
rect 204898 507832 204904 507844
rect 204956 507832 204962 507884
rect 88978 504364 88984 504416
rect 89036 504404 89042 504416
rect 115198 504404 115204 504416
rect 89036 504376 115204 504404
rect 89036 504364 89042 504376
rect 115198 504364 115204 504376
rect 115256 504364 115262 504416
rect 189718 500216 189724 500268
rect 189776 500256 189782 500268
rect 201862 500256 201868 500268
rect 189776 500228 201868 500256
rect 189776 500216 189782 500228
rect 201862 500216 201868 500228
rect 201920 500216 201926 500268
rect 236638 497428 236644 497480
rect 236696 497468 236702 497480
rect 249058 497468 249064 497480
rect 236696 497440 249064 497468
rect 236696 497428 236702 497440
rect 249058 497428 249064 497440
rect 249116 497428 249122 497480
rect 138014 496068 138020 496120
rect 138072 496108 138078 496120
rect 149698 496108 149704 496120
rect 138072 496080 149704 496108
rect 138072 496068 138078 496080
rect 149698 496068 149704 496080
rect 149756 496068 149762 496120
rect 80698 491920 80704 491972
rect 80756 491960 80762 491972
rect 88978 491960 88984 491972
rect 80756 491932 88984 491960
rect 80756 491920 80762 491932
rect 88978 491920 88984 491932
rect 89036 491920 89042 491972
rect 128538 490560 128544 490612
rect 128596 490600 128602 490612
rect 138014 490600 138020 490612
rect 128596 490572 138020 490600
rect 128596 490560 128602 490572
rect 138014 490560 138020 490572
rect 138072 490560 138078 490612
rect 125686 487500 125692 487552
rect 125744 487540 125750 487552
rect 128538 487540 128544 487552
rect 125744 487512 128544 487540
rect 125744 487500 125750 487512
rect 128538 487500 128544 487512
rect 128596 487500 128602 487552
rect 120718 485052 120724 485104
rect 120776 485092 120782 485104
rect 125686 485092 125692 485104
rect 120776 485064 125692 485092
rect 120776 485052 120782 485064
rect 125686 485052 125692 485064
rect 125744 485052 125750 485104
rect 77938 478864 77944 478916
rect 77996 478904 78002 478916
rect 80698 478904 80704 478916
rect 77996 478876 80704 478904
rect 77996 478864 78002 478876
rect 80698 478864 80704 478876
rect 80756 478864 80762 478916
rect 235258 474648 235264 474700
rect 235316 474688 235322 474700
rect 236638 474688 236644 474700
rect 235316 474660 236644 474688
rect 235316 474648 235322 474660
rect 236638 474648 236644 474660
rect 236696 474648 236702 474700
rect 232498 466420 232504 466472
rect 232556 466460 232562 466472
rect 235258 466460 235264 466472
rect 232556 466432 235264 466460
rect 232556 466420 232562 466432
rect 235258 466420 235264 466432
rect 235316 466420 235322 466472
rect 115566 466080 115572 466132
rect 115624 466120 115630 466132
rect 120718 466120 120724 466132
rect 115624 466092 120724 466120
rect 115624 466080 115630 466092
rect 120718 466080 120724 466092
rect 120776 466080 120782 466132
rect 3234 462544 3240 462596
rect 3292 462584 3298 462596
rect 8938 462584 8944 462596
rect 3292 462556 8944 462584
rect 3292 462544 3298 462556
rect 8938 462544 8944 462556
rect 8996 462544 9002 462596
rect 109678 462340 109684 462392
rect 109736 462380 109742 462392
rect 115566 462380 115572 462392
rect 109736 462352 115572 462380
rect 109736 462340 109742 462352
rect 115566 462340 115572 462352
rect 115624 462340 115630 462392
rect 64138 457444 64144 457496
rect 64196 457484 64202 457496
rect 77938 457484 77944 457496
rect 64196 457456 77944 457484
rect 64196 457444 64202 457456
rect 77938 457444 77944 457456
rect 77996 457444 78002 457496
rect 400858 456764 400864 456816
rect 400916 456804 400922 456816
rect 580166 456804 580172 456816
rect 400916 456776 580172 456804
rect 400916 456764 400922 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 226426 446360 226432 446412
rect 226484 446400 226490 446412
rect 232498 446400 232504 446412
rect 226484 446372 232504 446400
rect 226484 446360 226490 446372
rect 232498 446360 232504 446372
rect 232556 446360 232562 446412
rect 201586 445816 201592 445868
rect 201644 445856 201650 445868
rect 203518 445856 203524 445868
rect 201644 445828 203524 445856
rect 201644 445816 201650 445828
rect 203518 445816 203524 445828
rect 203576 445816 203582 445868
rect 199378 445340 199384 445392
rect 199436 445380 199442 445392
rect 201586 445380 201592 445392
rect 199436 445352 201592 445380
rect 199436 445340 199442 445352
rect 201586 445340 201592 445352
rect 201644 445340 201650 445392
rect 48406 445000 48412 445052
rect 48464 445040 48470 445052
rect 64138 445040 64144 445052
rect 48464 445012 64144 445040
rect 48464 445000 48470 445012
rect 64138 445000 64144 445012
rect 64196 445000 64202 445052
rect 104158 442892 104164 442944
rect 104216 442932 104222 442944
rect 105538 442932 105544 442944
rect 104216 442904 105544 442932
rect 104216 442892 104222 442904
rect 105538 442892 105544 442904
rect 105596 442892 105602 442944
rect 225598 442416 225604 442468
rect 225656 442456 225662 442468
rect 226426 442456 226432 442468
rect 225656 442428 226432 442456
rect 225656 442416 225662 442428
rect 226426 442416 226432 442428
rect 226484 442416 226490 442468
rect 46658 442280 46664 442332
rect 46716 442320 46722 442332
rect 48406 442320 48412 442332
rect 46716 442292 48412 442320
rect 46716 442280 46722 442292
rect 48406 442280 48412 442292
rect 48464 442280 48470 442332
rect 184198 438880 184204 438932
rect 184256 438920 184262 438932
rect 189718 438920 189724 438932
rect 184256 438892 189724 438920
rect 184256 438880 184262 438892
rect 189718 438880 189724 438892
rect 189776 438880 189782 438932
rect 199378 437492 199384 437504
rect 197372 437464 199384 437492
rect 196618 437384 196624 437436
rect 196676 437424 196682 437436
rect 197372 437424 197400 437464
rect 199378 437452 199384 437464
rect 199436 437452 199442 437504
rect 196676 437396 197400 437424
rect 196676 437384 196682 437396
rect 45002 436840 45008 436892
rect 45060 436880 45066 436892
rect 46658 436880 46664 436892
rect 45060 436852 46664 436880
rect 45060 436840 45066 436852
rect 46658 436840 46664 436852
rect 46716 436840 46722 436892
rect 174538 435344 174544 435396
rect 174596 435384 174602 435396
rect 184198 435384 184204 435396
rect 174596 435356 184204 435384
rect 174596 435344 174602 435356
rect 184198 435344 184204 435356
rect 184256 435344 184262 435396
rect 396718 430584 396724 430636
rect 396776 430624 396782 430636
rect 579982 430624 579988 430636
rect 396776 430596 579988 430624
rect 396776 430584 396782 430596
rect 579982 430584 579988 430596
rect 580040 430584 580046 430636
rect 169018 429836 169024 429888
rect 169076 429876 169082 429888
rect 174538 429876 174544 429888
rect 169076 429848 174544 429876
rect 169076 429836 169082 429848
rect 174538 429836 174544 429848
rect 174596 429836 174602 429888
rect 193858 426844 193864 426896
rect 193916 426884 193922 426896
rect 196618 426884 196624 426896
rect 193916 426856 196624 426884
rect 193916 426844 193922 426856
rect 196618 426844 196624 426856
rect 196676 426844 196682 426896
rect 106918 423580 106924 423632
rect 106976 423620 106982 423632
rect 109678 423620 109684 423632
rect 106976 423592 109684 423620
rect 106976 423580 106982 423592
rect 109678 423580 109684 423592
rect 109736 423580 109742 423632
rect 3142 422900 3148 422952
rect 3200 422940 3206 422952
rect 6270 422940 6276 422952
rect 3200 422912 6276 422940
rect 3200 422900 3206 422912
rect 6270 422900 6276 422912
rect 6328 422900 6334 422952
rect 3142 409844 3148 409896
rect 3200 409884 3206 409896
rect 10318 409884 10324 409896
rect 3200 409856 10324 409884
rect 3200 409844 3206 409856
rect 10318 409844 10324 409856
rect 10376 409844 10382 409896
rect 166258 407532 166264 407584
rect 166316 407572 166322 407584
rect 169018 407572 169024 407584
rect 166316 407544 169024 407572
rect 166316 407532 166322 407544
rect 169018 407532 169024 407544
rect 169076 407532 169082 407584
rect 224218 407328 224224 407380
rect 224276 407368 224282 407380
rect 225598 407368 225604 407380
rect 224276 407340 225604 407368
rect 224276 407328 224282 407340
rect 225598 407328 225604 407340
rect 225656 407328 225662 407380
rect 193858 404376 193864 404388
rect 191852 404348 193864 404376
rect 191098 404268 191104 404320
rect 191156 404308 191162 404320
rect 191852 404308 191880 404348
rect 193858 404336 193864 404348
rect 193916 404336 193922 404388
rect 418798 404336 418804 404388
rect 418856 404376 418862 404388
rect 580074 404376 580080 404388
rect 418856 404348 580080 404376
rect 418856 404336 418862 404348
rect 580074 404336 580080 404348
rect 580132 404336 580138 404388
rect 191156 404280 191880 404308
rect 191156 404268 191162 404280
rect 69658 396720 69664 396772
rect 69716 396760 69722 396772
rect 136634 396760 136640 396772
rect 69716 396732 136640 396760
rect 69716 396720 69722 396732
rect 136634 396720 136640 396732
rect 136692 396720 136698 396772
rect 223022 395972 223028 396024
rect 223080 396012 223086 396024
rect 224218 396012 224224 396024
rect 223080 395984 224224 396012
rect 223080 395972 223086 395984
rect 224218 395972 224224 395984
rect 224276 395972 224282 396024
rect 95878 392572 95884 392624
rect 95936 392612 95942 392624
rect 106918 392612 106924 392624
rect 95936 392584 106924 392612
rect 95936 392572 95942 392584
rect 106918 392572 106924 392584
rect 106976 392572 106982 392624
rect 163498 391960 163504 392012
rect 163556 392000 163562 392012
rect 166258 392000 166264 392012
rect 163556 391972 166264 392000
rect 163556 391960 163562 391972
rect 166258 391960 166264 391972
rect 166316 391960 166322 392012
rect 209038 387064 209044 387116
rect 209096 387104 209102 387116
rect 223022 387104 223028 387116
rect 209096 387076 223028 387104
rect 209096 387064 209102 387076
rect 223022 387064 223028 387076
rect 223080 387064 223086 387116
rect 191098 385064 191104 385076
rect 190426 385036 191104 385064
rect 68278 384956 68284 385008
rect 68336 384996 68342 385008
rect 69658 384996 69664 385008
rect 68336 384968 69664 384996
rect 68336 384956 68342 384968
rect 69658 384956 69664 384968
rect 69716 384956 69722 385008
rect 186958 384956 186964 385008
rect 187016 384996 187022 385008
rect 190426 384996 190454 385036
rect 191098 385024 191104 385036
rect 191156 385024 191162 385076
rect 187016 384968 190454 384996
rect 187016 384956 187022 384968
rect 78582 382916 78588 382968
rect 78640 382956 78646 382968
rect 95878 382956 95884 382968
rect 78640 382928 95884 382956
rect 78640 382916 78646 382928
rect 95878 382916 95884 382928
rect 95936 382916 95942 382968
rect 205634 382236 205640 382288
rect 205692 382276 205698 382288
rect 209038 382276 209044 382288
rect 205692 382248 209044 382276
rect 205692 382236 205698 382248
rect 209038 382236 209044 382248
rect 209096 382236 209102 382288
rect 102778 381488 102784 381540
rect 102836 381528 102842 381540
rect 163498 381528 163504 381540
rect 102836 381500 163504 381528
rect 102836 381488 102842 381500
rect 163498 381488 163504 381500
rect 163556 381488 163562 381540
rect 64230 380128 64236 380180
rect 64288 380168 64294 380180
rect 78582 380168 78588 380180
rect 64288 380140 78588 380168
rect 64288 380128 64294 380140
rect 78582 380128 78588 380140
rect 78640 380128 78646 380180
rect 102134 379176 102140 379228
rect 102192 379216 102198 379228
rect 104158 379216 104164 379228
rect 102192 379188 104164 379216
rect 102192 379176 102198 379188
rect 104158 379176 104164 379188
rect 104216 379176 104222 379228
rect 396810 378156 396816 378208
rect 396868 378196 396874 378208
rect 580074 378196 580080 378208
rect 396868 378168 580080 378196
rect 396868 378156 396874 378168
rect 580074 378156 580080 378168
rect 580132 378156 580138 378208
rect 202138 378088 202144 378140
rect 202196 378128 202202 378140
rect 205634 378128 205640 378140
rect 202196 378100 205640 378128
rect 202196 378088 202202 378100
rect 205634 378088 205640 378100
rect 205692 378088 205698 378140
rect 101398 374960 101404 375012
rect 101456 375000 101462 375012
rect 102134 375000 102140 375012
rect 101456 374972 102140 375000
rect 101456 374960 101462 374972
rect 102134 374960 102140 374972
rect 102192 374960 102198 375012
rect 202138 372620 202144 372632
rect 200086 372592 202144 372620
rect 197998 372512 198004 372564
rect 198056 372552 198062 372564
rect 200086 372552 200114 372592
rect 202138 372580 202144 372592
rect 202196 372580 202202 372632
rect 198056 372524 200114 372552
rect 198056 372512 198062 372524
rect 3234 371220 3240 371272
rect 3292 371260 3298 371272
rect 24118 371260 24124 371272
rect 3292 371232 24124 371260
rect 3292 371220 3298 371232
rect 24118 371220 24124 371232
rect 24176 371220 24182 371272
rect 95878 369860 95884 369912
rect 95936 369900 95942 369912
rect 102778 369900 102784 369912
rect 95936 369872 102784 369900
rect 95936 369860 95942 369872
rect 102778 369860 102784 369872
rect 102836 369860 102842 369912
rect 398098 364352 398104 364404
rect 398156 364392 398162 364404
rect 579798 364392 579804 364404
rect 398156 364364 579804 364392
rect 398156 364352 398162 364364
rect 579798 364352 579804 364364
rect 579856 364352 579862 364404
rect 100018 362924 100024 362976
rect 100076 362964 100082 362976
rect 101398 362964 101404 362976
rect 100076 362936 101404 362964
rect 100076 362924 100082 362936
rect 101398 362924 101404 362936
rect 101456 362924 101462 362976
rect 65426 358776 65432 358828
rect 65484 358816 65490 358828
rect 68278 358816 68284 358828
rect 65484 358788 68284 358816
rect 65484 358776 65490 358788
rect 68278 358776 68284 358788
rect 68336 358776 68342 358828
rect 64138 358096 64144 358148
rect 64196 358136 64202 358148
rect 65426 358136 65432 358148
rect 64196 358108 65432 358136
rect 64196 358096 64202 358108
rect 65426 358096 65432 358108
rect 65484 358096 65490 358148
rect 3234 357552 3240 357604
rect 3292 357592 3298 357604
rect 6362 357592 6368 357604
rect 3292 357564 6368 357592
rect 3292 357552 3298 357564
rect 6362 357552 6368 357564
rect 6420 357552 6426 357604
rect 60182 356464 60188 356516
rect 60240 356504 60246 356516
rect 64230 356504 64236 356516
rect 60240 356476 64236 356504
rect 60240 356464 60246 356476
rect 64230 356464 64236 356476
rect 64288 356464 64294 356516
rect 49602 353948 49608 354000
rect 49660 353988 49666 354000
rect 60182 353988 60188 354000
rect 49660 353960 60188 353988
rect 49660 353948 49666 353960
rect 60182 353948 60188 353960
rect 60240 353948 60246 354000
rect 93118 352384 93124 352436
rect 93176 352424 93182 352436
rect 95878 352424 95884 352436
rect 93176 352396 95884 352424
rect 93176 352384 93182 352396
rect 95878 352384 95884 352396
rect 95936 352384 95942 352436
rect 417418 351908 417424 351960
rect 417476 351948 417482 351960
rect 580074 351948 580080 351960
rect 417476 351920 580080 351948
rect 417476 351908 417482 351920
rect 580074 351908 580080 351920
rect 580132 351908 580138 351960
rect 46198 350548 46204 350600
rect 46256 350588 46262 350600
rect 49602 350588 49608 350600
rect 46256 350560 49608 350588
rect 46256 350548 46262 350560
rect 49602 350548 49608 350560
rect 49660 350548 49666 350600
rect 185578 350548 185584 350600
rect 185636 350588 185642 350600
rect 186958 350588 186964 350600
rect 185636 350560 186964 350588
rect 185636 350548 185642 350560
rect 186958 350548 186964 350560
rect 187016 350548 187022 350600
rect 195238 346332 195244 346384
rect 195296 346372 195302 346384
rect 197998 346372 198004 346384
rect 195296 346344 198004 346372
rect 195296 346332 195302 346344
rect 197998 346332 198004 346344
rect 198056 346332 198062 346384
rect 45370 342932 45376 342984
rect 45428 342972 45434 342984
rect 46198 342972 46204 342984
rect 45428 342944 46204 342972
rect 45428 342932 45434 342944
rect 46198 342932 46204 342944
rect 46256 342932 46262 342984
rect 184198 338716 184204 338768
rect 184256 338756 184262 338768
rect 185578 338756 185584 338768
rect 184256 338728 185584 338756
rect 184256 338716 184262 338728
rect 185578 338716 185584 338728
rect 185636 338716 185642 338768
rect 94406 332120 94412 332172
rect 94464 332160 94470 332172
rect 100018 332160 100024 332172
rect 94464 332132 100024 332160
rect 94464 332120 94470 332132
rect 100018 332120 100024 332132
rect 100076 332120 100082 332172
rect 62850 331848 62856 331900
rect 62908 331888 62914 331900
rect 88334 331888 88340 331900
rect 62908 331860 88340 331888
rect 62908 331848 62914 331860
rect 88334 331848 88340 331860
rect 88392 331848 88398 331900
rect 91738 329400 91744 329452
rect 91796 329440 91802 329452
rect 94406 329440 94412 329452
rect 91796 329412 94412 329440
rect 91796 329400 91802 329412
rect 94406 329400 94412 329412
rect 94464 329400 94470 329452
rect 182818 329128 182824 329180
rect 182876 329168 182882 329180
rect 184198 329168 184204 329180
rect 182876 329140 184204 329168
rect 182876 329128 182882 329140
rect 184198 329128 184204 329140
rect 184256 329128 184262 329180
rect 194042 328040 194048 328092
rect 194100 328080 194106 328092
rect 195238 328080 195244 328092
rect 194100 328052 195244 328080
rect 194100 328040 194106 328052
rect 195238 328040 195244 328052
rect 195296 328040 195302 328092
rect 396994 324300 397000 324352
rect 397052 324340 397058 324352
rect 580074 324340 580080 324352
rect 397052 324312 580080 324340
rect 397052 324300 397058 324312
rect 580074 324300 580080 324312
rect 580132 324300 580138 324352
rect 183370 322192 183376 322244
rect 183428 322232 183434 322244
rect 194042 322232 194048 322244
rect 183428 322204 194048 322232
rect 183428 322192 183434 322204
rect 194042 322192 194048 322204
rect 194100 322192 194106 322244
rect 181438 320152 181444 320204
rect 181496 320192 181502 320204
rect 183370 320192 183376 320204
rect 181496 320164 183376 320192
rect 181496 320152 181502 320164
rect 183370 320152 183376 320164
rect 183428 320152 183434 320204
rect 62758 319404 62764 319456
rect 62816 319444 62822 319456
rect 64138 319444 64144 319456
rect 62816 319416 64144 319444
rect 62816 319404 62822 319416
rect 64138 319404 64144 319416
rect 64196 319404 64202 319456
rect 3234 318792 3240 318844
rect 3292 318832 3298 318844
rect 24210 318832 24216 318844
rect 3292 318804 24216 318832
rect 3292 318792 3298 318804
rect 24210 318792 24216 318804
rect 24268 318792 24274 318844
rect 61470 318384 61476 318436
rect 61528 318424 61534 318436
rect 62850 318424 62856 318436
rect 61528 318396 62856 318424
rect 61528 318384 61534 318396
rect 62850 318384 62856 318396
rect 62908 318384 62914 318436
rect 84838 315256 84844 315308
rect 84896 315296 84902 315308
rect 104894 315296 104900 315308
rect 84896 315268 104900 315296
rect 84896 315256 84902 315268
rect 104894 315256 104900 315268
rect 104952 315256 104958 315308
rect 179506 314644 179512 314696
rect 179564 314684 179570 314696
rect 181438 314684 181444 314696
rect 179564 314656 181444 314684
rect 179564 314644 179570 314656
rect 181438 314644 181444 314656
rect 181496 314644 181502 314696
rect 398190 311856 398196 311908
rect 398248 311896 398254 311908
rect 580074 311896 580080 311908
rect 398248 311868 580080 311896
rect 398248 311856 398254 311868
rect 580074 311856 580080 311868
rect 580132 311856 580138 311908
rect 59998 311176 60004 311228
rect 60056 311216 60062 311228
rect 61470 311216 61476 311228
rect 60056 311188 61476 311216
rect 60056 311176 60062 311188
rect 61470 311176 61476 311188
rect 61528 311176 61534 311228
rect 178678 309544 178684 309596
rect 178736 309584 178742 309596
rect 179506 309584 179512 309596
rect 178736 309556 179512 309584
rect 178736 309544 178742 309556
rect 179506 309544 179512 309556
rect 179564 309544 179570 309596
rect 176654 305192 176660 305244
rect 176712 305232 176718 305244
rect 178678 305232 178684 305244
rect 176712 305204 178684 305232
rect 176712 305192 176718 305204
rect 178678 305192 178684 305204
rect 178736 305192 178742 305244
rect 170122 304240 170128 304292
rect 170180 304280 170186 304292
rect 176654 304280 176660 304292
rect 170180 304252 176660 304280
rect 170180 304240 170186 304252
rect 176654 304240 176660 304252
rect 176712 304240 176718 304292
rect 180058 302064 180064 302116
rect 180116 302104 180122 302116
rect 182818 302104 182824 302116
rect 180116 302076 182824 302104
rect 180116 302064 180122 302076
rect 182818 302064 182824 302076
rect 182876 302064 182882 302116
rect 169018 300228 169024 300280
rect 169076 300268 169082 300280
rect 170122 300268 170128 300280
rect 169076 300240 170128 300268
rect 169076 300228 169082 300240
rect 170122 300228 170128 300240
rect 170180 300228 170186 300280
rect 60826 299412 60832 299464
rect 60884 299452 60890 299464
rect 62758 299452 62764 299464
rect 60884 299424 62764 299452
rect 60884 299412 60890 299424
rect 62758 299412 62764 299424
rect 62816 299412 62822 299464
rect 414658 298120 414664 298172
rect 414716 298160 414722 298172
rect 580074 298160 580080 298172
rect 414716 298132 580080 298160
rect 414716 298120 414722 298132
rect 580074 298120 580080 298132
rect 580132 298120 580138 298172
rect 90358 298052 90364 298104
rect 90416 298092 90422 298104
rect 93118 298092 93124 298104
rect 90416 298064 93124 298092
rect 90416 298052 90422 298064
rect 93118 298052 93124 298064
rect 93176 298052 93182 298104
rect 167638 295332 167644 295384
rect 167696 295372 167702 295384
rect 169018 295372 169024 295384
rect 167696 295344 169024 295372
rect 167696 295332 167702 295344
rect 169018 295332 169024 295344
rect 169076 295332 169082 295384
rect 60090 293972 60096 294024
rect 60148 294012 60154 294024
rect 60826 294012 60832 294024
rect 60148 293984 60832 294012
rect 60148 293972 60154 293984
rect 60826 293972 60832 293984
rect 60884 293972 60890 294024
rect 2774 292816 2780 292868
rect 2832 292856 2838 292868
rect 4890 292856 4896 292868
rect 2832 292828 4896 292856
rect 2832 292816 2838 292828
rect 4890 292816 4896 292828
rect 4948 292816 4954 292868
rect 58618 291116 58624 291168
rect 58676 291156 58682 291168
rect 59998 291156 60004 291168
rect 58676 291128 60004 291156
rect 58676 291116 58682 291128
rect 59998 291116 60004 291128
rect 60056 291116 60062 291168
rect 175642 290980 175648 291032
rect 175700 291020 175706 291032
rect 180058 291020 180064 291032
rect 175700 290992 180064 291020
rect 175700 290980 175706 290992
rect 180058 290980 180064 290992
rect 180116 290980 180122 291032
rect 169018 289076 169024 289128
rect 169076 289116 169082 289128
rect 175642 289116 175648 289128
rect 169076 289088 175648 289116
rect 169076 289076 169082 289088
rect 175642 289076 175648 289088
rect 175700 289076 175706 289128
rect 57238 287648 57244 287700
rect 57296 287688 57302 287700
rect 71774 287688 71780 287700
rect 57296 287660 71780 287688
rect 57296 287648 57302 287660
rect 71774 287648 71780 287660
rect 71832 287648 71838 287700
rect 58618 284356 58624 284368
rect 56612 284328 58624 284356
rect 56502 284248 56508 284300
rect 56560 284288 56566 284300
rect 56612 284288 56640 284328
rect 58618 284316 58624 284328
rect 58676 284316 58682 284368
rect 84838 284356 84844 284368
rect 84166 284328 84844 284356
rect 56560 284260 56640 284288
rect 56560 284248 56566 284260
rect 82078 284248 82084 284300
rect 82136 284288 82142 284300
rect 84166 284288 84194 284328
rect 84838 284316 84844 284328
rect 84896 284316 84902 284368
rect 82136 284260 84194 284288
rect 82136 284248 82142 284260
rect 57974 282888 57980 282940
rect 58032 282928 58038 282940
rect 60090 282928 60096 282940
rect 58032 282900 60096 282928
rect 58032 282888 58038 282900
rect 60090 282888 60096 282900
rect 60148 282888 60154 282940
rect 54294 281120 54300 281172
rect 54352 281160 54358 281172
rect 56502 281160 56508 281172
rect 54352 281132 56508 281160
rect 54352 281120 54358 281132
rect 56502 281120 56508 281132
rect 56560 281120 56566 281172
rect 59998 280780 60004 280832
rect 60056 280820 60062 280832
rect 169754 280820 169760 280832
rect 60056 280792 169760 280820
rect 60056 280780 60062 280792
rect 169754 280780 169760 280792
rect 169812 280780 169818 280832
rect 53282 278808 53288 278860
rect 53340 278848 53346 278860
rect 54294 278848 54300 278860
rect 53340 278820 54300 278848
rect 53340 278808 53346 278820
rect 54294 278808 54300 278820
rect 54352 278808 54358 278860
rect 54478 278808 54484 278860
rect 54536 278848 54542 278860
rect 57882 278848 57888 278860
rect 54536 278820 57888 278848
rect 54536 278808 54542 278820
rect 57882 278808 57888 278820
rect 57940 278808 57946 278860
rect 167638 278780 167644 278792
rect 164252 278752 167644 278780
rect 162854 278672 162860 278724
rect 162912 278712 162918 278724
rect 164252 278712 164280 278752
rect 167638 278740 167644 278752
rect 167696 278740 167702 278792
rect 162912 278684 164280 278712
rect 162912 278672 162918 278684
rect 57238 277420 57244 277432
rect 55232 277392 57244 277420
rect 53834 277312 53840 277364
rect 53892 277352 53898 277364
rect 55232 277352 55260 277392
rect 57238 277380 57244 277392
rect 57296 277380 57302 277432
rect 53892 277324 55260 277352
rect 53892 277312 53898 277324
rect 55858 276632 55864 276684
rect 55916 276672 55922 276684
rect 82078 276672 82084 276684
rect 55916 276644 82084 276672
rect 55916 276632 55922 276644
rect 82078 276632 82084 276644
rect 82136 276632 82142 276684
rect 53098 274660 53104 274712
rect 53156 274700 53162 274712
rect 53834 274700 53840 274712
rect 53156 274672 53840 274700
rect 53156 274660 53162 274672
rect 53834 274660 53840 274672
rect 53892 274660 53898 274712
rect 159358 274660 159364 274712
rect 159416 274700 159422 274712
rect 162854 274700 162860 274712
rect 159416 274672 162860 274700
rect 159416 274660 159422 274672
rect 162854 274660 162860 274672
rect 162912 274660 162918 274712
rect 169018 273272 169024 273284
rect 167012 273244 169024 273272
rect 166258 273164 166264 273216
rect 166316 273204 166322 273216
rect 167012 273204 167040 273244
rect 169018 273232 169024 273244
rect 169076 273232 169082 273284
rect 166316 273176 167040 273204
rect 166316 273164 166322 273176
rect 51810 272076 51816 272128
rect 51868 272116 51874 272128
rect 53282 272116 53288 272128
rect 51868 272088 53288 272116
rect 51868 272076 51874 272088
rect 53282 272076 53288 272088
rect 53340 272076 53346 272128
rect 396902 271872 396908 271924
rect 396960 271912 396966 271924
rect 579798 271912 579804 271924
rect 396960 271884 579804 271912
rect 396960 271872 396966 271884
rect 579798 271872 579804 271884
rect 579856 271872 579862 271924
rect 86954 270648 86960 270700
rect 87012 270688 87018 270700
rect 90358 270688 90364 270700
rect 87012 270660 90364 270688
rect 87012 270648 87018 270660
rect 90358 270648 90364 270660
rect 90416 270648 90422 270700
rect 77938 268336 77944 268388
rect 77996 268376 78002 268388
rect 86954 268376 86960 268388
rect 77996 268348 86960 268376
rect 77996 268336 78002 268348
rect 86954 268336 86960 268348
rect 87012 268336 87018 268388
rect 56594 268064 56600 268116
rect 56652 268104 56658 268116
rect 59998 268104 60004 268116
rect 56652 268076 60004 268104
rect 56652 268064 56658 268076
rect 59998 268064 60004 268076
rect 60056 268064 60062 268116
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 40678 266404 40684 266416
rect 3108 266376 40684 266404
rect 3108 266364 3114 266376
rect 40678 266364 40684 266376
rect 40736 266364 40742 266416
rect 53190 266364 53196 266416
rect 53248 266404 53254 266416
rect 54478 266404 54484 266416
rect 53248 266376 54484 266404
rect 53248 266364 53254 266376
rect 54478 266364 54484 266376
rect 54536 266364 54542 266416
rect 54570 266364 54576 266416
rect 54628 266404 54634 266416
rect 55858 266404 55864 266416
rect 54628 266376 55864 266404
rect 54628 266364 54634 266376
rect 55858 266364 55864 266376
rect 55916 266364 55922 266416
rect 56502 264976 56508 264988
rect 52472 264948 56508 264976
rect 51718 264868 51724 264920
rect 51776 264908 51782 264920
rect 52472 264908 52500 264948
rect 56502 264936 56508 264948
rect 56560 264936 56566 264988
rect 164234 264936 164240 264988
rect 164292 264976 164298 264988
rect 166258 264976 166264 264988
rect 164292 264948 166264 264976
rect 164292 264936 164298 264948
rect 166258 264936 166264 264948
rect 166316 264936 166322 264988
rect 51776 264880 52500 264908
rect 51776 264868 51782 264880
rect 49694 263576 49700 263628
rect 49752 263616 49758 263628
rect 51810 263616 51816 263628
rect 49752 263588 51816 263616
rect 49752 263576 49758 263588
rect 51810 263576 51816 263588
rect 51868 263576 51874 263628
rect 53282 263576 53288 263628
rect 53340 263616 53346 263628
rect 54570 263616 54576 263628
rect 53340 263588 54576 263616
rect 53340 263576 53346 263588
rect 54570 263576 54576 263588
rect 54628 263576 54634 263628
rect 156598 261944 156604 261996
rect 156656 261984 156662 261996
rect 159358 261984 159364 261996
rect 156656 261956 159364 261984
rect 156656 261944 156662 261956
rect 159358 261944 159364 261956
rect 159416 261944 159422 261996
rect 162118 260040 162124 260092
rect 162176 260080 162182 260092
rect 164234 260080 164240 260092
rect 162176 260052 164240 260080
rect 162176 260040 162182 260052
rect 164234 260040 164240 260052
rect 164292 260040 164298 260092
rect 46934 258952 46940 259004
rect 46992 258992 46998 259004
rect 49694 258992 49700 259004
rect 46992 258964 49700 258992
rect 46992 258952 46998 258964
rect 49694 258952 49700 258964
rect 49752 258952 49758 259004
rect 398282 258068 398288 258120
rect 398340 258108 398346 258120
rect 579982 258108 579988 258120
rect 398340 258080 579988 258108
rect 398340 258068 398346 258080
rect 579982 258068 579988 258080
rect 580040 258068 580046 258120
rect 53282 256748 53288 256760
rect 51092 256720 53288 256748
rect 50430 256640 50436 256692
rect 50488 256680 50494 256692
rect 51092 256680 51120 256720
rect 53282 256708 53288 256720
rect 53340 256708 53346 256760
rect 154022 256708 154028 256760
rect 154080 256748 154086 256760
rect 156598 256748 156604 256760
rect 154080 256720 156604 256748
rect 154080 256708 154086 256720
rect 156598 256708 156604 256720
rect 156656 256708 156662 256760
rect 50488 256652 51120 256680
rect 50488 256640 50494 256652
rect 45554 255280 45560 255332
rect 45612 255320 45618 255332
rect 46934 255320 46940 255332
rect 45612 255292 46940 255320
rect 45612 255280 45618 255292
rect 46934 255280 46940 255292
rect 46992 255280 46998 255332
rect 151078 255280 151084 255332
rect 151136 255320 151142 255332
rect 154022 255320 154028 255332
rect 151136 255292 154028 255320
rect 151136 255280 151142 255292
rect 154022 255280 154028 255292
rect 154080 255280 154086 255332
rect 53190 254028 53196 254040
rect 47044 254000 53196 254028
rect 3142 253920 3148 253972
rect 3200 253960 3206 253972
rect 22738 253960 22744 253972
rect 3200 253932 22744 253960
rect 3200 253920 3206 253932
rect 22738 253920 22744 253932
rect 22796 253920 22802 253972
rect 46198 253852 46204 253904
rect 46256 253892 46262 253904
rect 47044 253892 47072 254000
rect 53190 253988 53196 254000
rect 53248 253988 53254 254040
rect 47578 253920 47584 253972
rect 47636 253960 47642 253972
rect 50430 253960 50436 253972
rect 47636 253932 50436 253960
rect 47636 253920 47642 253932
rect 50430 253920 50436 253932
rect 50488 253920 50494 253972
rect 46256 253864 47072 253892
rect 46256 253852 46262 253864
rect 51810 252560 51816 252612
rect 51868 252600 51874 252612
rect 53098 252600 53104 252612
rect 51868 252572 53104 252600
rect 51868 252560 51874 252572
rect 53098 252560 53104 252572
rect 53156 252560 53162 252612
rect 50338 250792 50344 250844
rect 50396 250832 50402 250844
rect 51810 250832 51816 250844
rect 50396 250804 51816 250832
rect 50396 250792 50402 250804
rect 51810 250792 51816 250804
rect 51868 250792 51874 250844
rect 75178 249704 75184 249756
rect 75236 249744 75242 249756
rect 77938 249744 77944 249756
rect 75236 249716 77944 249744
rect 75236 249704 75242 249716
rect 77938 249704 77944 249716
rect 77996 249704 78002 249756
rect 89162 249704 89168 249756
rect 89220 249744 89226 249756
rect 91738 249744 91744 249756
rect 89220 249716 91744 249744
rect 89220 249704 89226 249716
rect 91738 249704 91744 249716
rect 91796 249704 91802 249756
rect 160094 245896 160100 245948
rect 160152 245936 160158 245948
rect 162118 245936 162124 245948
rect 160152 245908 162124 245936
rect 160152 245896 160158 245908
rect 162118 245896 162124 245908
rect 162176 245896 162182 245948
rect 45830 245624 45836 245676
rect 45888 245664 45894 245676
rect 47578 245664 47584 245676
rect 45888 245636 47584 245664
rect 45888 245624 45894 245636
rect 47578 245624 47584 245636
rect 47636 245624 47642 245676
rect 49694 245624 49700 245676
rect 49752 245664 49758 245676
rect 51718 245664 51724 245676
rect 49752 245636 51724 245664
rect 49752 245624 49758 245636
rect 51718 245624 51724 245636
rect 51776 245624 51782 245676
rect 145190 245624 145196 245676
rect 145248 245664 145254 245676
rect 151078 245664 151084 245676
rect 145248 245636 151084 245664
rect 145248 245624 145254 245636
rect 151078 245624 151084 245636
rect 151136 245624 151142 245676
rect 45186 245556 45192 245608
rect 45244 245596 45250 245608
rect 46198 245596 46204 245608
rect 45244 245568 46204 245596
rect 45244 245556 45250 245568
rect 46198 245556 46204 245568
rect 46256 245556 46262 245608
rect 81434 244876 81440 244928
rect 81492 244916 81498 244928
rect 89162 244916 89168 244928
rect 81492 244888 89168 244916
rect 81492 244876 81498 244888
rect 89162 244876 89168 244888
rect 89220 244876 89226 244928
rect 413278 244264 413284 244316
rect 413336 244304 413342 244316
rect 579982 244304 579988 244316
rect 413336 244276 579988 244304
rect 413336 244264 413342 244276
rect 579982 244264 579988 244276
rect 580040 244264 580046 244316
rect 75086 242972 75092 243024
rect 75144 243012 75150 243024
rect 81434 243012 81440 243024
rect 75144 242984 81440 243012
rect 75144 242972 75150 242984
rect 81434 242972 81440 242984
rect 81492 242972 81498 243024
rect 49694 242944 49700 242956
rect 48332 242916 49700 242944
rect 45738 242836 45744 242888
rect 45796 242876 45802 242888
rect 48332 242876 48360 242916
rect 49694 242904 49700 242916
rect 49752 242904 49758 242956
rect 45796 242848 48360 242876
rect 45796 242836 45802 242848
rect 142982 241816 142988 241868
rect 143040 241856 143046 241868
rect 145190 241856 145196 241868
rect 143040 241828 145196 241856
rect 143040 241816 143046 241828
rect 145190 241816 145196 241828
rect 145248 241816 145254 241868
rect 45094 240932 45100 240984
rect 45152 240972 45158 240984
rect 75086 240972 75092 240984
rect 45152 240944 75092 240972
rect 45152 240932 45158 240944
rect 75086 240932 75092 240944
rect 75144 240932 75150 240984
rect 44910 240864 44916 240916
rect 44968 240904 44974 240916
rect 75178 240904 75184 240916
rect 44968 240876 75184 240904
rect 44968 240864 44974 240876
rect 75178 240864 75184 240876
rect 75236 240864 75242 240916
rect 45370 240796 45376 240848
rect 45428 240836 45434 240848
rect 142982 240836 142988 240848
rect 45428 240808 142988 240836
rect 45428 240796 45434 240808
rect 142982 240796 142988 240808
rect 143040 240796 143046 240848
rect 46842 240728 46848 240780
rect 46900 240768 46906 240780
rect 160094 240768 160100 240780
rect 46900 240740 160100 240768
rect 46900 240728 46906 240740
rect 160094 240728 160100 240740
rect 160152 240728 160158 240780
rect 45646 240388 45652 240440
rect 45704 240428 45710 240440
rect 50338 240428 50344 240440
rect 45704 240400 50344 240428
rect 45704 240388 45710 240400
rect 50338 240388 50344 240400
rect 50396 240388 50402 240440
rect 2774 240184 2780 240236
rect 2832 240224 2838 240236
rect 4982 240224 4988 240236
rect 2832 240196 4988 240224
rect 2832 240184 2838 240196
rect 4982 240184 4988 240196
rect 5040 240184 5046 240236
rect 395338 239980 395344 240032
rect 395396 240020 395402 240032
rect 396626 240020 396632 240032
rect 395396 239992 396632 240020
rect 395396 239980 395402 239992
rect 396626 239980 396632 239992
rect 396684 239980 396690 240032
rect 395430 239776 395436 239828
rect 395488 239816 395494 239828
rect 395488 239788 395936 239816
rect 395488 239776 395494 239788
rect 44818 239708 44824 239760
rect 44876 239748 44882 239760
rect 46842 239748 46848 239760
rect 44876 239720 46848 239748
rect 44876 239708 44882 239720
rect 46842 239708 46848 239720
rect 46900 239708 46906 239760
rect 45462 238756 45468 238808
rect 45520 238796 45526 238808
rect 45830 238796 45836 238808
rect 45520 238768 45836 238796
rect 45520 238756 45526 238768
rect 45830 238756 45836 238768
rect 45888 238756 45894 238808
rect 395908 238728 395936 239788
rect 396534 238728 396540 238740
rect 395908 238700 396540 238728
rect 396534 238688 396540 238700
rect 396592 238688 396598 238740
rect 45738 233044 45744 233096
rect 45796 233084 45802 233096
rect 45796 233056 64874 233084
rect 45796 233044 45802 233056
rect 45646 232976 45652 233028
rect 45704 233016 45710 233028
rect 45704 232988 58940 233016
rect 45704 232976 45710 232988
rect 45462 232908 45468 232960
rect 45520 232948 45526 232960
rect 45830 232948 45836 232960
rect 45520 232920 45836 232948
rect 45520 232908 45526 232920
rect 45830 232908 45836 232920
rect 45888 232908 45894 232960
rect 58912 232812 58940 232988
rect 58912 232784 62804 232812
rect 62776 232416 62804 232784
rect 62758 232364 62764 232416
rect 62816 232364 62822 232416
rect 64846 232404 64874 233056
rect 80698 232404 80704 232416
rect 64846 232376 80704 232404
rect 80698 232364 80704 232376
rect 80756 232364 80762 232416
rect 395430 232364 395436 232416
rect 395488 232404 395494 232416
rect 396534 232404 396540 232416
rect 395488 232376 396540 232404
rect 395488 232364 395494 232376
rect 396534 232364 396540 232376
rect 396592 232364 396598 232416
rect 45370 231956 45376 232008
rect 45428 231996 45434 232008
rect 46566 231996 46572 232008
rect 45428 231968 46572 231996
rect 45428 231956 45434 231968
rect 46566 231956 46572 231968
rect 46624 231956 46630 232008
rect 45094 231888 45100 231940
rect 45152 231928 45158 231940
rect 45152 231900 46980 231928
rect 45152 231888 45158 231900
rect 45278 231820 45284 231872
rect 45336 231860 45342 231872
rect 46842 231860 46848 231872
rect 45336 231832 46848 231860
rect 45336 231820 45342 231832
rect 46842 231820 46848 231832
rect 46900 231820 46906 231872
rect 46952 231792 46980 231900
rect 393958 231820 393964 231872
rect 394016 231860 394022 231872
rect 580074 231860 580080 231872
rect 394016 231832 580080 231860
rect 394016 231820 394022 231832
rect 580074 231820 580080 231832
rect 580132 231820 580138 231872
rect 49142 231792 49148 231804
rect 46952 231764 49148 231792
rect 49142 231752 49148 231764
rect 49200 231752 49206 231804
rect 44818 231684 44824 231736
rect 44876 231724 44882 231736
rect 49786 231724 49792 231736
rect 44876 231696 49792 231724
rect 44876 231684 44882 231696
rect 49786 231684 49792 231696
rect 49844 231684 49850 231736
rect 45830 231140 45836 231192
rect 45888 231180 45894 231192
rect 142154 231180 142160 231192
rect 45888 231152 142160 231180
rect 45888 231140 45894 231152
rect 142154 231140 142160 231152
rect 142212 231140 142218 231192
rect 3326 231072 3332 231124
rect 3384 231112 3390 231124
rect 180794 231112 180800 231124
rect 3384 231084 180800 231112
rect 3384 231072 3390 231084
rect 180794 231072 180800 231084
rect 180852 231072 180858 231124
rect 385678 231072 385684 231124
rect 385736 231112 385742 231124
rect 396626 231112 396632 231124
rect 385736 231084 396632 231112
rect 385736 231072 385742 231084
rect 396626 231072 396632 231084
rect 396684 231072 396690 231124
rect 45186 231004 45192 231056
rect 45244 231044 45250 231056
rect 64874 231044 64880 231056
rect 45244 231016 64880 231044
rect 45244 231004 45250 231016
rect 64874 231004 64880 231016
rect 64932 231004 64938 231056
rect 46566 230460 46572 230512
rect 46624 230500 46630 230512
rect 46624 230472 46980 230500
rect 46624 230460 46630 230472
rect 46952 230432 46980 230472
rect 49694 230432 49700 230444
rect 46952 230404 49700 230432
rect 49694 230392 49700 230404
rect 49752 230392 49758 230444
rect 395338 230392 395344 230444
rect 395396 230432 395402 230444
rect 396442 230432 396448 230444
rect 395396 230404 396448 230432
rect 395396 230392 395402 230404
rect 396442 230392 396448 230404
rect 396500 230392 396506 230444
rect 49786 230120 49792 230172
rect 49844 230160 49850 230172
rect 55122 230160 55128 230172
rect 49844 230132 55128 230160
rect 49844 230120 49850 230132
rect 55122 230120 55128 230132
rect 55180 230120 55186 230172
rect 166258 229712 166264 229764
rect 166316 229752 166322 229764
rect 176654 229752 176660 229764
rect 166316 229724 176660 229752
rect 166316 229712 166322 229724
rect 176654 229712 176660 229724
rect 176712 229712 176718 229764
rect 45002 229032 45008 229084
rect 45060 229072 45066 229084
rect 47026 229072 47032 229084
rect 45060 229044 47032 229072
rect 45060 229032 45066 229044
rect 47026 229032 47032 229044
rect 47084 229032 47090 229084
rect 157978 228420 157984 228472
rect 158036 228460 158042 228472
rect 266538 228460 266544 228472
rect 158036 228432 266544 228460
rect 158036 228420 158042 228432
rect 266538 228420 266544 228432
rect 266596 228420 266602 228472
rect 297358 228420 297364 228472
rect 297416 228460 297422 228472
rect 327074 228460 327080 228472
rect 297416 228432 327080 228460
rect 297416 228420 297422 228432
rect 327074 228420 327080 228432
rect 327132 228420 327138 228472
rect 236638 228352 236644 228404
rect 236696 228392 236702 228404
rect 386506 228392 386512 228404
rect 236696 228364 386512 228392
rect 236696 228352 236702 228364
rect 386506 228352 386512 228364
rect 386564 228352 386570 228404
rect 142154 228284 142160 228336
rect 142212 228324 142218 228336
rect 143534 228324 143540 228336
rect 142212 228296 143540 228324
rect 142212 228284 142218 228296
rect 143534 228284 143540 228296
rect 143592 228284 143598 228336
rect 395430 227780 395436 227792
rect 393286 227752 395436 227780
rect 391198 227672 391204 227724
rect 391256 227712 391262 227724
rect 393286 227712 393314 227752
rect 395430 227740 395436 227752
rect 395488 227740 395494 227792
rect 391256 227684 393314 227712
rect 391256 227672 391262 227684
rect 49694 226312 49700 226364
rect 49752 226352 49758 226364
rect 49752 226324 52500 226352
rect 49752 226312 49758 226324
rect 44910 226244 44916 226296
rect 44968 226284 44974 226296
rect 50430 226284 50436 226296
rect 44968 226256 50436 226284
rect 44968 226244 44974 226256
rect 50430 226244 50436 226256
rect 50488 226244 50494 226296
rect 52472 226284 52500 226324
rect 64874 226312 64880 226364
rect 64932 226352 64938 226364
rect 69566 226352 69572 226364
rect 64932 226324 69572 226352
rect 64932 226312 64938 226324
rect 69566 226312 69572 226324
rect 69624 226312 69630 226364
rect 56226 226284 56232 226296
rect 52472 226256 56232 226284
rect 56226 226244 56232 226256
rect 56284 226244 56290 226296
rect 47026 225700 47032 225752
rect 47084 225740 47090 225752
rect 53834 225740 53840 225752
rect 47084 225712 53840 225740
rect 47084 225700 47090 225712
rect 53834 225700 53840 225712
rect 53892 225700 53898 225752
rect 46934 224952 46940 225004
rect 46992 224992 46998 225004
rect 46992 224964 48360 224992
rect 46992 224952 46998 224964
rect 48332 224924 48360 224964
rect 50338 224924 50344 224936
rect 48332 224896 50344 224924
rect 50338 224884 50344 224896
rect 50396 224884 50402 224936
rect 389818 223048 389824 223100
rect 389876 223088 389882 223100
rect 394326 223088 394332 223100
rect 389876 223060 394332 223088
rect 389876 223048 389882 223060
rect 394326 223048 394332 223060
rect 394384 223048 394390 223100
rect 55214 222912 55220 222964
rect 55272 222952 55278 222964
rect 57330 222952 57336 222964
rect 55272 222924 57336 222952
rect 55272 222912 55278 222924
rect 57330 222912 57336 222924
rect 57388 222912 57394 222964
rect 53834 222844 53840 222896
rect 53892 222884 53898 222896
rect 69658 222884 69664 222896
rect 53892 222856 69664 222884
rect 53892 222844 53898 222856
rect 69658 222844 69664 222856
rect 69716 222844 69722 222896
rect 49142 222164 49148 222216
rect 49200 222204 49206 222216
rect 49200 222176 51120 222204
rect 49200 222164 49206 222176
rect 51092 222136 51120 222176
rect 55122 222136 55128 222148
rect 51092 222108 55128 222136
rect 55122 222096 55128 222108
rect 55180 222096 55186 222148
rect 56226 222096 56232 222148
rect 56284 222136 56290 222148
rect 57238 222136 57244 222148
rect 56284 222108 57244 222136
rect 56284 222096 56290 222108
rect 57238 222096 57244 222108
rect 57296 222096 57302 222148
rect 378042 220804 378048 220856
rect 378100 220844 378106 220856
rect 385678 220844 385684 220856
rect 378100 220816 385684 220844
rect 378100 220804 378106 220816
rect 385678 220804 385684 220816
rect 385736 220804 385742 220856
rect 69658 220056 69664 220108
rect 69716 220096 69722 220108
rect 79318 220096 79324 220108
rect 69716 220068 79324 220096
rect 69716 220056 69722 220068
rect 79318 220056 79324 220068
rect 79376 220056 79382 220108
rect 143534 220056 143540 220108
rect 143592 220096 143598 220108
rect 158622 220096 158628 220108
rect 143592 220068 158628 220096
rect 143592 220056 143598 220068
rect 158622 220056 158628 220068
rect 158680 220056 158686 220108
rect 69658 218628 69664 218680
rect 69716 218668 69722 218680
rect 71866 218668 71872 218680
rect 69716 218640 71872 218668
rect 69716 218628 69722 218640
rect 71866 218628 71872 218640
rect 71924 218628 71930 218680
rect 119430 218016 119436 218068
rect 119488 218056 119494 218068
rect 580074 218056 580080 218068
rect 119488 218028 580080 218056
rect 119488 218016 119494 218028
rect 580074 218016 580080 218028
rect 580132 218016 580138 218068
rect 57330 217268 57336 217320
rect 57388 217308 57394 217320
rect 67542 217308 67548 217320
rect 57388 217280 67548 217308
rect 57388 217268 57394 217280
rect 67542 217268 67548 217280
rect 67600 217268 67606 217320
rect 62758 215908 62764 215960
rect 62816 215948 62822 215960
rect 70394 215948 70400 215960
rect 62816 215920 70400 215948
rect 62816 215908 62822 215920
rect 70394 215908 70400 215920
rect 70452 215908 70458 215960
rect 367738 215908 367744 215960
rect 367796 215948 367802 215960
rect 378042 215948 378048 215960
rect 367796 215920 378048 215948
rect 367796 215908 367802 215920
rect 378042 215908 378048 215920
rect 378100 215908 378106 215960
rect 67542 215568 67548 215620
rect 67600 215608 67606 215620
rect 69014 215608 69020 215620
rect 67600 215580 69020 215608
rect 67600 215568 67606 215580
rect 69014 215568 69020 215580
rect 69072 215568 69078 215620
rect 50430 215092 50436 215144
rect 50488 215132 50494 215144
rect 54478 215132 54484 215144
rect 50488 215104 54484 215132
rect 50488 215092 50494 215104
rect 54478 215092 54484 215104
rect 54536 215092 54542 215144
rect 71866 214548 71872 214600
rect 71924 214588 71930 214600
rect 73982 214588 73988 214600
rect 71924 214560 73988 214588
rect 71924 214548 71930 214560
rect 73982 214548 73988 214560
rect 74040 214548 74046 214600
rect 80698 214548 80704 214600
rect 80756 214588 80762 214600
rect 91738 214588 91744 214600
rect 80756 214560 91744 214588
rect 80756 214548 80762 214560
rect 91738 214548 91744 214560
rect 91796 214548 91802 214600
rect 55214 214072 55220 214124
rect 55272 214112 55278 214124
rect 57330 214112 57336 214124
rect 55272 214084 57336 214112
rect 55272 214072 55278 214084
rect 57330 214072 57336 214084
rect 57388 214072 57394 214124
rect 3326 213936 3332 213988
rect 3384 213976 3390 213988
rect 180978 213976 180984 213988
rect 3384 213948 180984 213976
rect 3384 213936 3390 213948
rect 180978 213936 180984 213948
rect 181036 213936 181042 213988
rect 50338 213868 50344 213920
rect 50396 213908 50402 213920
rect 53098 213908 53104 213920
rect 50396 213880 53104 213908
rect 50396 213868 50402 213880
rect 53098 213868 53104 213880
rect 53156 213868 53162 213920
rect 158714 213868 158720 213920
rect 158772 213908 158778 213920
rect 160094 213908 160100 213920
rect 158772 213880 160100 213908
rect 158772 213868 158778 213880
rect 160094 213868 160100 213880
rect 160152 213868 160158 213920
rect 69014 213528 69020 213580
rect 69072 213568 69078 213580
rect 71038 213568 71044 213580
rect 69072 213540 71044 213568
rect 69072 213528 69078 213540
rect 71038 213528 71044 213540
rect 71096 213528 71102 213580
rect 70394 212984 70400 213036
rect 70452 213024 70458 213036
rect 73798 213024 73804 213036
rect 70452 212996 73804 213024
rect 70452 212984 70458 212996
rect 73798 212984 73804 212996
rect 73856 212984 73862 213036
rect 389910 212168 389916 212220
rect 389968 212208 389974 212220
rect 391198 212208 391204 212220
rect 389968 212180 391204 212208
rect 389968 212168 389974 212180
rect 391198 212168 391204 212180
rect 391256 212168 391262 212220
rect 160094 211148 160100 211200
rect 160152 211188 160158 211200
rect 160152 211160 161474 211188
rect 160152 211148 160158 211160
rect 57238 211080 57244 211132
rect 57296 211120 57302 211132
rect 58618 211120 58624 211132
rect 57296 211092 58624 211120
rect 57296 211080 57302 211092
rect 58618 211080 58624 211092
rect 58676 211080 58682 211132
rect 161446 211120 161474 211160
rect 162854 211120 162860 211132
rect 161446 211092 162860 211120
rect 162854 211080 162860 211092
rect 162912 211080 162918 211132
rect 378778 210400 378784 210452
rect 378836 210440 378842 210452
rect 395338 210440 395344 210452
rect 378836 210412 395344 210440
rect 378836 210400 378842 210412
rect 395338 210400 395344 210412
rect 395396 210400 395402 210452
rect 73982 209720 73988 209772
rect 74040 209760 74046 209772
rect 75454 209760 75460 209772
rect 74040 209732 75460 209760
rect 74040 209720 74046 209732
rect 75454 209720 75460 209732
rect 75512 209720 75518 209772
rect 53098 209448 53104 209500
rect 53156 209488 53162 209500
rect 54570 209488 54576 209500
rect 53156 209460 54576 209488
rect 53156 209448 53162 209460
rect 54570 209448 54576 209460
rect 54628 209448 54634 209500
rect 162854 209108 162860 209160
rect 162912 209148 162918 209160
rect 164234 209148 164240 209160
rect 162912 209120 164240 209148
rect 162912 209108 162918 209120
rect 164234 209108 164240 209120
rect 164292 209108 164298 209160
rect 79318 209040 79324 209092
rect 79376 209080 79382 209092
rect 91094 209080 91100 209092
rect 79376 209052 91100 209080
rect 79376 209040 79382 209052
rect 91094 209040 91100 209052
rect 91152 209040 91158 209092
rect 71038 208904 71044 208956
rect 71096 208944 71102 208956
rect 73890 208944 73896 208956
rect 71096 208916 73896 208944
rect 71096 208904 71102 208916
rect 73890 208904 73896 208916
rect 73948 208904 73954 208956
rect 57330 208360 57336 208412
rect 57388 208400 57394 208412
rect 57388 208372 59400 208400
rect 57388 208360 57394 208372
rect 59372 208332 59400 208372
rect 63494 208332 63500 208344
rect 59372 208304 63500 208332
rect 63494 208292 63500 208304
rect 63552 208292 63558 208344
rect 75454 208292 75460 208344
rect 75512 208332 75518 208344
rect 77570 208332 77576 208344
rect 75512 208304 77576 208332
rect 75512 208292 75518 208304
rect 77570 208292 77576 208304
rect 77628 208292 77634 208344
rect 91738 208292 91744 208344
rect 91796 208332 91802 208344
rect 95142 208332 95148 208344
rect 91796 208304 95148 208332
rect 91796 208292 91802 208304
rect 95142 208292 95148 208304
rect 95200 208292 95206 208344
rect 164234 206660 164240 206712
rect 164292 206700 164298 206712
rect 166350 206700 166356 206712
rect 164292 206672 166356 206700
rect 164292 206660 164298 206672
rect 166350 206660 166356 206672
rect 166408 206660 166414 206712
rect 91094 206252 91100 206304
rect 91152 206292 91158 206304
rect 104710 206292 104716 206304
rect 91152 206264 104716 206292
rect 91152 206252 91158 206264
rect 104710 206252 104716 206264
rect 104768 206252 104774 206304
rect 356698 206252 356704 206304
rect 356756 206292 356762 206304
rect 367738 206292 367744 206304
rect 356756 206264 367744 206292
rect 356756 206252 356762 206264
rect 367738 206252 367744 206264
rect 367796 206252 367802 206304
rect 189718 205640 189724 205692
rect 189776 205680 189782 205692
rect 580074 205680 580080 205692
rect 189776 205652 580080 205680
rect 189776 205640 189782 205652
rect 580074 205640 580080 205652
rect 580132 205640 580138 205692
rect 95142 204892 95148 204944
rect 95200 204932 95206 204944
rect 106642 204932 106648 204944
rect 95200 204904 106648 204932
rect 95200 204892 95206 204904
rect 106642 204892 106648 204904
rect 106700 204892 106706 204944
rect 77570 204824 77576 204876
rect 77628 204864 77634 204876
rect 80054 204864 80060 204876
rect 77628 204836 80060 204864
rect 77628 204824 77634 204836
rect 80054 204824 80060 204836
rect 80112 204824 80118 204876
rect 63494 204212 63500 204264
rect 63552 204252 63558 204264
rect 65518 204252 65524 204264
rect 63552 204224 65524 204252
rect 63552 204212 63558 204224
rect 65518 204212 65524 204224
rect 65576 204212 65582 204264
rect 58618 202784 58624 202836
rect 58676 202824 58682 202836
rect 63494 202824 63500 202836
rect 58676 202796 63500 202824
rect 58676 202784 58682 202796
rect 63494 202784 63500 202796
rect 63552 202784 63558 202836
rect 80054 202784 80060 202836
rect 80112 202824 80118 202836
rect 81802 202824 81808 202836
rect 80112 202796 81808 202824
rect 80112 202784 80118 202796
rect 81802 202784 81808 202796
rect 81860 202784 81866 202836
rect 104710 202784 104716 202836
rect 104768 202824 104774 202836
rect 108666 202824 108672 202836
rect 104768 202796 108672 202824
rect 104768 202784 104774 202796
rect 108666 202784 108672 202796
rect 108724 202784 108730 202836
rect 106642 202716 106648 202768
rect 106700 202756 106706 202768
rect 110230 202756 110236 202768
rect 106700 202728 110236 202756
rect 106700 202716 106706 202728
rect 110230 202716 110236 202728
rect 110288 202716 110294 202768
rect 2958 201492 2964 201544
rect 3016 201532 3022 201544
rect 22830 201532 22836 201544
rect 3016 201504 22836 201532
rect 3016 201492 3022 201504
rect 22830 201492 22836 201504
rect 22888 201492 22894 201544
rect 45554 201424 45560 201476
rect 45612 201464 45618 201476
rect 47578 201464 47584 201476
rect 45612 201436 47584 201464
rect 45612 201424 45618 201436
rect 47578 201424 47584 201436
rect 47636 201424 47642 201476
rect 73798 199384 73804 199436
rect 73856 199424 73862 199436
rect 81434 199424 81440 199436
rect 73856 199396 81440 199424
rect 73856 199384 73862 199396
rect 81434 199384 81440 199396
rect 81492 199384 81498 199436
rect 81802 199384 81808 199436
rect 81860 199424 81866 199436
rect 88978 199424 88984 199436
rect 81860 199396 88984 199424
rect 81860 199384 81866 199396
rect 88978 199384 88984 199396
rect 89036 199384 89042 199436
rect 155954 199384 155960 199436
rect 156012 199424 156018 199436
rect 296714 199424 296720 199436
rect 156012 199396 296720 199424
rect 156012 199384 156018 199396
rect 296714 199384 296720 199396
rect 296772 199384 296778 199436
rect 63494 197956 63500 198008
rect 63552 197996 63558 198008
rect 69566 197996 69572 198008
rect 63552 197968 69572 197996
rect 63552 197956 63558 197968
rect 69566 197956 69572 197968
rect 69624 197956 69630 198008
rect 110230 197956 110236 198008
rect 110288 197996 110294 198008
rect 117314 197996 117320 198008
rect 110288 197968 117320 197996
rect 110288 197956 110294 197968
rect 117314 197956 117320 197968
rect 117372 197956 117378 198008
rect 148962 197956 148968 198008
rect 149020 197996 149026 198008
rect 207014 197996 207020 198008
rect 149020 197968 207020 197996
rect 149020 197956 149026 197968
rect 207014 197956 207020 197968
rect 207072 197956 207078 198008
rect 108666 197480 108672 197532
rect 108724 197520 108730 197532
rect 111058 197520 111064 197532
rect 108724 197492 111064 197520
rect 108724 197480 108730 197492
rect 111058 197480 111064 197492
rect 111116 197480 111122 197532
rect 154482 197412 154488 197464
rect 154540 197452 154546 197464
rect 155954 197452 155960 197464
rect 154540 197424 155960 197452
rect 154540 197412 154546 197424
rect 155954 197412 155960 197424
rect 156012 197412 156018 197464
rect 54570 197276 54576 197328
rect 54628 197316 54634 197328
rect 56502 197316 56508 197328
rect 54628 197288 56508 197316
rect 54628 197276 54634 197288
rect 56502 197276 56508 197288
rect 56560 197276 56566 197328
rect 73890 197276 73896 197328
rect 73948 197316 73954 197328
rect 76282 197316 76288 197328
rect 73948 197288 76288 197316
rect 73948 197276 73954 197288
rect 76282 197276 76288 197288
rect 76340 197276 76346 197328
rect 152734 197276 152740 197328
rect 152792 197316 152798 197328
rect 157978 197316 157984 197328
rect 152792 197288 157984 197316
rect 152792 197276 152798 197288
rect 157978 197276 157984 197288
rect 158036 197276 158042 197328
rect 147950 196732 147956 196784
rect 148008 196772 148014 196784
rect 166258 196772 166264 196784
rect 148008 196744 166264 196772
rect 148008 196732 148014 196744
rect 166258 196732 166264 196744
rect 166316 196732 166322 196784
rect 160830 196664 160836 196716
rect 160888 196704 160894 196716
rect 236638 196704 236644 196716
rect 160888 196676 236644 196704
rect 160888 196664 160894 196676
rect 236638 196664 236644 196676
rect 236696 196664 236702 196716
rect 81434 196596 81440 196648
rect 81492 196636 81498 196648
rect 88334 196636 88340 196648
rect 81492 196608 88340 196636
rect 81492 196596 81498 196608
rect 88334 196596 88340 196608
rect 88392 196596 88398 196648
rect 151170 196596 151176 196648
rect 151228 196636 151234 196648
rect 235994 196636 236000 196648
rect 151228 196608 236000 196636
rect 151228 196596 151234 196608
rect 235994 196596 236000 196608
rect 236052 196596 236058 196648
rect 69566 196120 69572 196172
rect 69624 196160 69630 196172
rect 71774 196160 71780 196172
rect 69624 196132 71780 196160
rect 69624 196120 69630 196132
rect 71774 196120 71780 196132
rect 71832 196120 71838 196172
rect 56594 195916 56600 195968
rect 56652 195956 56658 195968
rect 138106 195956 138112 195968
rect 56652 195928 138112 195956
rect 56652 195916 56658 195928
rect 138106 195916 138112 195928
rect 138164 195916 138170 195968
rect 157518 195916 157524 195968
rect 157576 195956 157582 195968
rect 356054 195956 356060 195968
rect 157576 195928 356060 195956
rect 157576 195916 157582 195928
rect 356054 195916 356060 195928
rect 356112 195916 356118 195968
rect 76282 195848 76288 195900
rect 76340 195888 76346 195900
rect 77938 195888 77944 195900
rect 76340 195860 77944 195888
rect 76340 195848 76346 195860
rect 77938 195848 77944 195860
rect 77996 195848 78002 195900
rect 86954 195848 86960 195900
rect 87012 195888 87018 195900
rect 139394 195888 139400 195900
rect 87012 195860 139400 195888
rect 87012 195848 87018 195860
rect 139394 195848 139400 195860
rect 139452 195848 139458 195900
rect 157426 195848 157432 195900
rect 157484 195888 157490 195900
rect 297358 195888 297364 195900
rect 157484 195860 297364 195888
rect 157484 195848 157490 195860
rect 297358 195848 297364 195860
rect 297416 195848 297422 195900
rect 115934 194556 115940 194608
rect 115992 194596 115998 194608
rect 140774 194596 140780 194608
rect 115992 194568 140780 194596
rect 115992 194556 115998 194568
rect 140774 194556 140780 194568
rect 140832 194556 140838 194608
rect 117314 194352 117320 194404
rect 117372 194392 117378 194404
rect 120718 194392 120724 194404
rect 117372 194364 120724 194392
rect 117372 194352 117378 194364
rect 120718 194352 120724 194364
rect 120776 194352 120782 194404
rect 88334 193536 88340 193588
rect 88392 193576 88398 193588
rect 91738 193576 91744 193588
rect 88392 193548 91744 193576
rect 88392 193536 88398 193548
rect 91738 193536 91744 193548
rect 91796 193536 91802 193588
rect 71774 193128 71780 193180
rect 71832 193168 71838 193180
rect 74258 193168 74264 193180
rect 71832 193140 74264 193168
rect 71832 193128 71838 193140
rect 74258 193128 74264 193140
rect 74316 193128 74322 193180
rect 166350 193128 166356 193180
rect 166408 193168 166414 193180
rect 168466 193168 168472 193180
rect 166408 193140 168472 193168
rect 166408 193128 166414 193140
rect 168466 193128 168472 193140
rect 168524 193128 168530 193180
rect 180058 191836 180064 191888
rect 180116 191876 180122 191888
rect 580074 191876 580080 191888
rect 180116 191848 580080 191876
rect 180116 191836 180122 191848
rect 580074 191836 580080 191848
rect 580132 191836 580138 191888
rect 140958 190992 140964 191004
rect 140792 190964 140964 190992
rect 88978 190612 88984 190664
rect 89036 190652 89042 190664
rect 93854 190652 93860 190664
rect 89036 190624 93860 190652
rect 89036 190612 89042 190624
rect 93854 190612 93860 190624
rect 93912 190612 93918 190664
rect 140792 190528 140820 190964
rect 140958 190952 140964 190964
rect 141016 190952 141022 191004
rect 140774 190476 140780 190528
rect 140832 190476 140838 190528
rect 144454 190476 144460 190528
rect 144512 190516 144518 190528
rect 144512 190488 145052 190516
rect 144512 190476 144518 190488
rect 140774 190340 140780 190392
rect 140832 190340 140838 190392
rect 140792 190244 140820 190340
rect 145024 190324 145052 190488
rect 145006 190272 145012 190324
rect 145064 190272 145070 190324
rect 140866 190244 140872 190256
rect 140792 190216 140872 190244
rect 140866 190204 140872 190216
rect 140924 190204 140930 190256
rect 120718 189252 120724 189304
rect 120776 189292 120782 189304
rect 123662 189292 123668 189304
rect 120776 189264 123668 189292
rect 120776 189252 120782 189264
rect 123662 189252 123668 189264
rect 123720 189252 123726 189304
rect 144638 188912 144644 188964
rect 144696 188952 144702 188964
rect 145006 188952 145012 188964
rect 144696 188924 145012 188952
rect 144696 188912 144702 188924
rect 145006 188912 145012 188924
rect 145064 188912 145070 188964
rect 93854 187892 93860 187944
rect 93912 187932 93918 187944
rect 95878 187932 95884 187944
rect 93912 187904 95884 187932
rect 93912 187892 93918 187904
rect 95878 187892 95884 187904
rect 95936 187892 95942 187944
rect 3326 187688 3332 187740
rect 3384 187728 3390 187740
rect 116578 187728 116584 187740
rect 3384 187700 116584 187728
rect 3384 187688 3390 187700
rect 116578 187688 116584 187700
rect 116636 187688 116642 187740
rect 166166 187620 166172 187672
rect 166224 187660 166230 187672
rect 399478 187660 399484 187672
rect 166224 187632 399484 187660
rect 166224 187620 166230 187632
rect 399478 187620 399484 187632
rect 399536 187620 399542 187672
rect 54478 186940 54484 186992
rect 54536 186980 54542 186992
rect 68278 186980 68284 186992
rect 54536 186952 68284 186980
rect 54536 186940 54542 186952
rect 68278 186940 68284 186952
rect 68336 186940 68342 186992
rect 371234 186940 371240 186992
rect 371292 186980 371298 186992
rect 389818 186980 389824 186992
rect 371292 186952 389824 186980
rect 371292 186940 371298 186952
rect 389818 186940 389824 186952
rect 389876 186940 389882 186992
rect 56594 186396 56600 186448
rect 56652 186436 56658 186448
rect 58618 186436 58624 186448
rect 56652 186408 58624 186436
rect 56652 186396 56658 186408
rect 58618 186396 58624 186408
rect 58676 186396 58682 186448
rect 387794 186328 387800 186380
rect 387852 186368 387858 186380
rect 389910 186368 389916 186380
rect 387852 186340 389916 186368
rect 387852 186328 387858 186340
rect 389910 186328 389916 186340
rect 389968 186328 389974 186380
rect 74258 186260 74264 186312
rect 74316 186300 74322 186312
rect 76558 186300 76564 186312
rect 74316 186272 76564 186300
rect 74316 186260 74322 186272
rect 76558 186260 76564 186272
rect 76616 186260 76622 186312
rect 111058 186260 111064 186312
rect 111116 186300 111122 186312
rect 113818 186300 113824 186312
rect 111116 186272 113824 186300
rect 111116 186260 111122 186272
rect 113818 186260 113824 186272
rect 113876 186260 113882 186312
rect 168466 184832 168472 184884
rect 168524 184872 168530 184884
rect 170398 184872 170404 184884
rect 168524 184844 170404 184872
rect 168524 184832 168530 184844
rect 170398 184832 170404 184844
rect 170456 184832 170462 184884
rect 369118 183880 369124 183932
rect 369176 183920 369182 183932
rect 371234 183920 371240 183932
rect 369176 183892 371240 183920
rect 369176 183880 369182 183892
rect 371234 183880 371240 183892
rect 371292 183880 371298 183932
rect 387794 183580 387800 183592
rect 386432 183552 387800 183580
rect 385034 183472 385040 183524
rect 385092 183512 385098 183524
rect 386432 183512 386460 183552
rect 387794 183540 387800 183552
rect 387852 183540 387858 183592
rect 385092 183484 386460 183512
rect 385092 183472 385098 183484
rect 123662 182112 123668 182164
rect 123720 182152 123726 182164
rect 126514 182152 126520 182164
rect 123720 182124 126520 182152
rect 123720 182112 123726 182124
rect 126514 182112 126520 182124
rect 126572 182112 126578 182164
rect 144638 181500 144644 181552
rect 144696 181540 144702 181552
rect 145190 181540 145196 181552
rect 144696 181512 145196 181540
rect 144696 181500 144702 181512
rect 145190 181500 145196 181512
rect 145248 181500 145254 181552
rect 3234 181432 3240 181484
rect 3292 181472 3298 181484
rect 46198 181472 46204 181484
rect 3292 181444 46204 181472
rect 3292 181432 3298 181444
rect 46198 181432 46204 181444
rect 46256 181432 46262 181484
rect 121454 180072 121460 180124
rect 121512 180112 121518 180124
rect 136358 180112 136364 180124
rect 121512 180084 136364 180112
rect 121512 180072 121518 180084
rect 136358 180072 136364 180084
rect 136416 180072 136422 180124
rect 384298 179392 384304 179444
rect 384356 179432 384362 179444
rect 385034 179432 385040 179444
rect 384356 179404 385040 179432
rect 384356 179392 384362 179404
rect 385034 179392 385040 179404
rect 385092 179392 385098 179444
rect 158806 179324 158812 179376
rect 158864 179364 158870 179376
rect 165154 179364 165160 179376
rect 158864 179336 165160 179364
rect 158864 179324 158870 179336
rect 165154 179324 165160 179336
rect 165212 179364 165218 179376
rect 580810 179364 580816 179376
rect 165212 179336 580816 179364
rect 165212 179324 165218 179336
rect 580810 179324 580816 179336
rect 580868 179324 580874 179376
rect 113818 178916 113824 178968
rect 113876 178956 113882 178968
rect 117958 178956 117964 178968
rect 113876 178928 117964 178956
rect 113876 178916 113882 178928
rect 117958 178916 117964 178928
rect 118016 178916 118022 178968
rect 136358 178780 136364 178832
rect 136416 178820 136422 178832
rect 136726 178820 136732 178832
rect 136416 178792 136732 178820
rect 136416 178780 136422 178792
rect 136726 178780 136732 178792
rect 136784 178780 136790 178832
rect 124858 178712 124864 178764
rect 124916 178752 124922 178764
rect 136450 178752 136456 178764
rect 124916 178724 136456 178752
rect 124916 178712 124922 178724
rect 136450 178712 136456 178724
rect 136508 178712 136514 178764
rect 126514 178644 126520 178696
rect 126572 178684 126578 178696
rect 153930 178684 153936 178696
rect 126572 178656 153936 178684
rect 126572 178644 126578 178656
rect 153930 178644 153936 178656
rect 153988 178644 153994 178696
rect 135990 177760 135996 177812
rect 136048 177800 136054 177812
rect 136634 177800 136640 177812
rect 136048 177772 136640 177800
rect 136048 177760 136054 177772
rect 136634 177760 136640 177772
rect 136692 177760 136698 177812
rect 124214 177284 124220 177336
rect 124272 177324 124278 177336
rect 136450 177324 136456 177336
rect 124272 177296 136456 177324
rect 124272 177284 124278 177296
rect 136450 177284 136456 177296
rect 136508 177284 136514 177336
rect 68278 176604 68284 176656
rect 68336 176644 68342 176656
rect 76650 176644 76656 176656
rect 68336 176616 76656 176644
rect 68336 176604 68342 176616
rect 76650 176604 76656 176616
rect 76708 176604 76714 176656
rect 149238 176644 149244 176656
rect 146266 176616 149244 176644
rect 146266 176440 146294 176616
rect 149238 176604 149244 176616
rect 149296 176604 149302 176656
rect 144886 176412 146294 176440
rect 126974 176060 126980 176112
rect 127032 176100 127038 176112
rect 135990 176100 135996 176112
rect 127032 176072 135996 176100
rect 127032 176060 127038 176072
rect 135990 176060 135996 176072
rect 136048 176060 136054 176112
rect 141786 176060 141792 176112
rect 141844 176100 141850 176112
rect 144886 176100 144914 176412
rect 154390 176400 154396 176452
rect 154448 176440 154454 176452
rect 154448 176412 160508 176440
rect 154448 176400 154454 176412
rect 141844 176072 144914 176100
rect 141844 176060 141850 176072
rect 136358 176032 136364 176044
rect 128326 176004 136364 176032
rect 125594 175924 125600 175976
rect 125652 175964 125658 175976
rect 128326 175964 128354 176004
rect 136358 175992 136364 176004
rect 136416 175992 136422 176044
rect 160480 175976 160508 176412
rect 125652 175936 128354 175964
rect 125652 175924 125658 175936
rect 160462 175924 160468 175976
rect 160520 175924 160526 175976
rect 159174 175856 159180 175908
rect 159232 175896 159238 175908
rect 163590 175896 163596 175908
rect 159232 175868 163596 175896
rect 159232 175856 159238 175868
rect 163590 175856 163596 175868
rect 163648 175856 163654 175908
rect 159082 175788 159088 175840
rect 159140 175828 159146 175840
rect 162486 175828 162492 175840
rect 159140 175800 162492 175828
rect 159140 175788 159146 175800
rect 162486 175788 162492 175800
rect 162544 175788 162550 175840
rect 141602 175652 141608 175704
rect 141660 175692 141666 175704
rect 149330 175692 149336 175704
rect 141660 175664 149336 175692
rect 141660 175652 141666 175664
rect 149330 175652 149336 175664
rect 149388 175652 149394 175704
rect 144454 175516 144460 175568
rect 144512 175556 144518 175568
rect 148686 175556 148692 175568
rect 144512 175528 148692 175556
rect 144512 175516 144518 175528
rect 148686 175516 148692 175528
rect 148744 175516 148750 175568
rect 95878 175244 95884 175296
rect 95936 175284 95942 175296
rect 95936 175256 96660 175284
rect 95936 175244 95942 175256
rect 58618 175176 58624 175228
rect 58676 175216 58682 175228
rect 60642 175216 60648 175228
rect 58676 175188 60648 175216
rect 58676 175176 58682 175188
rect 60642 175176 60648 175188
rect 60700 175176 60706 175228
rect 77938 175176 77944 175228
rect 77996 175216 78002 175228
rect 79410 175216 79416 175228
rect 77996 175188 79416 175216
rect 77996 175176 78002 175188
rect 79410 175176 79416 175188
rect 79468 175176 79474 175228
rect 96632 175216 96660 175256
rect 100018 175216 100024 175228
rect 96632 175188 100024 175216
rect 100018 175176 100024 175188
rect 100076 175176 100082 175228
rect 128354 175176 128360 175228
rect 128412 175216 128418 175228
rect 136450 175216 136456 175228
rect 128412 175188 136456 175216
rect 128412 175176 128418 175188
rect 136450 175176 136456 175188
rect 136508 175176 136514 175228
rect 144086 174904 144092 174956
rect 144144 174944 144150 174956
rect 144144 174916 147674 174944
rect 144144 174904 144150 174916
rect 142062 174836 142068 174888
rect 142120 174836 142126 174888
rect 142080 174332 142108 174836
rect 147646 174536 147674 174916
rect 350534 174564 350540 174616
rect 350592 174604 350598 174616
rect 356698 174604 356704 174616
rect 350592 174576 356704 174604
rect 350592 174564 350598 174576
rect 356698 174564 356704 174576
rect 356756 174564 356762 174616
rect 161474 174536 161480 174548
rect 147646 174508 161480 174536
rect 161474 174496 161480 174508
rect 161532 174496 161538 174548
rect 142080 174304 165476 174332
rect 133874 173884 133880 173936
rect 133932 173924 133938 173936
rect 137278 173924 137284 173936
rect 133932 173896 137284 173924
rect 133932 173884 133938 173896
rect 137278 173884 137284 173896
rect 137336 173884 137342 173936
rect 165448 172984 165476 174304
rect 165430 172932 165436 172984
rect 165488 172932 165494 172984
rect 60642 172524 60648 172576
rect 60700 172564 60706 172576
rect 60700 172536 60872 172564
rect 60700 172524 60706 172536
rect 60844 172496 60872 172536
rect 131114 172524 131120 172576
rect 131172 172564 131178 172576
rect 136634 172564 136640 172576
rect 131172 172536 136640 172564
rect 131172 172524 131178 172536
rect 136634 172524 136640 172536
rect 136692 172524 136698 172576
rect 378778 172564 378784 172576
rect 376772 172536 378784 172564
rect 63494 172496 63500 172508
rect 60844 172468 63500 172496
rect 63494 172456 63500 172468
rect 63552 172456 63558 172508
rect 65518 172456 65524 172508
rect 65576 172496 65582 172508
rect 66254 172496 66260 172508
rect 65576 172468 66260 172496
rect 65576 172456 65582 172468
rect 66254 172456 66260 172468
rect 66312 172456 66318 172508
rect 76558 172456 76564 172508
rect 76616 172496 76622 172508
rect 79318 172496 79324 172508
rect 76616 172468 79324 172496
rect 76616 172456 76622 172468
rect 79318 172456 79324 172468
rect 79376 172456 79382 172508
rect 160462 172456 160468 172508
rect 160520 172496 160526 172508
rect 162118 172496 162124 172508
rect 160520 172468 162124 172496
rect 160520 172456 160526 172468
rect 162118 172456 162124 172468
rect 162176 172456 162182 172508
rect 376110 172456 376116 172508
rect 376168 172496 376174 172508
rect 376772 172496 376800 172536
rect 378778 172524 378784 172536
rect 378836 172524 378842 172576
rect 376168 172468 376800 172496
rect 376168 172456 376174 172468
rect 348418 172320 348424 172372
rect 348476 172360 348482 172372
rect 350534 172360 350540 172372
rect 348476 172332 350540 172360
rect 348476 172320 348482 172332
rect 350534 172320 350540 172332
rect 350592 172320 350598 172372
rect 135254 171912 135260 171964
rect 135312 171952 135318 171964
rect 138658 171952 138664 171964
rect 135312 171924 138664 171952
rect 135312 171912 135318 171924
rect 138658 171912 138664 171924
rect 138716 171912 138722 171964
rect 145466 171844 145472 171896
rect 145524 171884 145530 171896
rect 157978 171884 157984 171896
rect 145524 171856 157984 171884
rect 145524 171844 145530 171856
rect 157978 171844 157984 171856
rect 158036 171844 158042 171896
rect 47578 171776 47584 171828
rect 47636 171816 47642 171828
rect 61654 171816 61660 171828
rect 47636 171788 61660 171816
rect 47636 171776 47642 171788
rect 61654 171776 61660 171788
rect 61712 171776 61718 171828
rect 118694 171776 118700 171828
rect 118752 171816 118758 171828
rect 580166 171816 580172 171828
rect 118752 171788 580172 171816
rect 118752 171776 118758 171788
rect 580166 171776 580172 171788
rect 580224 171776 580230 171828
rect 91738 171164 91744 171216
rect 91796 171204 91802 171216
rect 94498 171204 94504 171216
rect 91796 171176 94504 171204
rect 91796 171164 91802 171176
rect 94498 171164 94504 171176
rect 94556 171164 94562 171216
rect 132494 171096 132500 171148
rect 132552 171136 132558 171148
rect 136726 171136 136732 171148
rect 132552 171108 136732 171136
rect 132552 171096 132558 171108
rect 136726 171096 136732 171108
rect 136784 171096 136790 171148
rect 138014 171096 138020 171148
rect 138072 171136 138078 171148
rect 140774 171136 140780 171148
rect 138072 171108 140780 171136
rect 138072 171096 138078 171108
rect 140774 171096 140780 171108
rect 140832 171096 140838 171148
rect 376018 170348 376024 170400
rect 376076 170388 376082 170400
rect 384298 170388 384304 170400
rect 376076 170360 384304 170388
rect 376076 170348 376082 170360
rect 384298 170348 384304 170360
rect 384356 170348 384362 170400
rect 152366 170280 152372 170332
rect 152424 170320 152430 170332
rect 156506 170320 156512 170332
rect 152424 170292 156512 170320
rect 152424 170280 152430 170292
rect 156506 170280 156512 170292
rect 156564 170280 156570 170332
rect 149330 170008 149336 170060
rect 149388 170048 149394 170060
rect 150434 170048 150440 170060
rect 149388 170020 150440 170048
rect 149388 170008 149394 170020
rect 150434 170008 150440 170020
rect 150492 170008 150498 170060
rect 63494 169532 63500 169584
rect 63552 169572 63558 169584
rect 65610 169572 65616 169584
rect 63552 169544 65616 169572
rect 63552 169532 63558 169544
rect 65610 169532 65616 169544
rect 65668 169532 65674 169584
rect 66254 169532 66260 169584
rect 66312 169572 66318 169584
rect 69658 169572 69664 169584
rect 66312 169544 69664 169572
rect 66312 169532 66318 169544
rect 69658 169532 69664 169544
rect 69716 169532 69722 169584
rect 61654 168716 61660 168768
rect 61712 168756 61718 168768
rect 63494 168756 63500 168768
rect 61712 168728 63500 168756
rect 61712 168716 61718 168728
rect 63494 168716 63500 168728
rect 63552 168716 63558 168768
rect 63494 166268 63500 166320
rect 63552 166308 63558 166320
rect 75178 166308 75184 166320
rect 63552 166280 75184 166308
rect 63552 166268 63558 166280
rect 75178 166268 75184 166280
rect 75236 166268 75242 166320
rect 142430 166268 142436 166320
rect 142488 166308 142494 166320
rect 142614 166308 142620 166320
rect 142488 166280 142620 166308
rect 142488 166268 142494 166280
rect 142614 166268 142620 166280
rect 142672 166268 142678 166320
rect 100018 165588 100024 165640
rect 100076 165628 100082 165640
rect 100076 165600 100800 165628
rect 100076 165588 100082 165600
rect 100772 165560 100800 165600
rect 188338 165588 188344 165640
rect 188396 165628 188402 165640
rect 580166 165628 580172 165640
rect 188396 165600 580172 165628
rect 188396 165588 188402 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 102778 165560 102784 165572
rect 100772 165532 102784 165560
rect 102778 165520 102784 165532
rect 102836 165520 102842 165572
rect 76650 164160 76656 164212
rect 76708 164200 76714 164212
rect 81802 164200 81808 164212
rect 76708 164172 81808 164200
rect 76708 164160 76714 164172
rect 81802 164160 81808 164172
rect 81860 164160 81866 164212
rect 94498 164160 94504 164212
rect 94556 164200 94562 164212
rect 97258 164200 97264 164212
rect 94556 164172 97264 164200
rect 94556 164160 94562 164172
rect 97258 164160 97264 164172
rect 97316 164160 97322 164212
rect 40678 163548 40684 163600
rect 40736 163588 40742 163600
rect 182358 163588 182364 163600
rect 40736 163560 182364 163588
rect 40736 163548 40742 163560
rect 182358 163548 182364 163560
rect 182416 163548 182422 163600
rect 24210 163480 24216 163532
rect 24268 163520 24274 163532
rect 182910 163520 182916 163532
rect 24268 163492 182916 163520
rect 24268 163480 24274 163492
rect 182910 163480 182916 163492
rect 182968 163480 182974 163532
rect 3326 162868 3332 162920
rect 3384 162908 3390 162920
rect 179506 162908 179512 162920
rect 3384 162880 179512 162908
rect 3384 162868 3390 162880
rect 179506 162868 179512 162880
rect 179564 162868 179570 162920
rect 65610 162800 65616 162852
rect 65668 162840 65674 162852
rect 71038 162840 71044 162852
rect 65668 162812 71044 162840
rect 65668 162800 65674 162812
rect 71038 162800 71044 162812
rect 71096 162800 71102 162852
rect 373994 162800 374000 162852
rect 374052 162840 374058 162852
rect 376110 162840 376116 162852
rect 374052 162812 376116 162840
rect 374052 162800 374058 162812
rect 376110 162800 376116 162812
rect 376168 162800 376174 162852
rect 81802 161236 81808 161288
rect 81860 161276 81866 161288
rect 85482 161276 85488 161288
rect 81860 161248 85488 161276
rect 81860 161236 81866 161248
rect 85482 161236 85488 161248
rect 85540 161236 85546 161288
rect 162118 160692 162124 160744
rect 162176 160732 162182 160744
rect 179414 160732 179420 160744
rect 162176 160704 179420 160732
rect 162176 160692 162182 160704
rect 179414 160692 179420 160704
rect 179472 160692 179478 160744
rect 75178 157972 75184 158024
rect 75236 158012 75242 158024
rect 86126 158012 86132 158024
rect 75236 157984 86132 158012
rect 75236 157972 75242 157984
rect 86126 157972 86132 157984
rect 86184 157972 86190 158024
rect 366726 157700 366732 157752
rect 366784 157740 366790 157752
rect 373902 157740 373908 157752
rect 366784 157712 373908 157740
rect 366784 157700 366790 157712
rect 373902 157700 373908 157712
rect 373960 157700 373966 157752
rect 375006 157360 375012 157412
rect 375064 157400 375070 157412
rect 376018 157400 376024 157412
rect 375064 157372 376024 157400
rect 375064 157360 375070 157372
rect 376018 157360 376024 157372
rect 376076 157360 376082 157412
rect 359458 156680 359464 156732
rect 359516 156720 359522 156732
rect 369118 156720 369124 156732
rect 359516 156692 369124 156720
rect 359516 156680 359522 156692
rect 369118 156680 369124 156692
rect 369176 156680 369182 156732
rect 353938 156612 353944 156664
rect 353996 156652 354002 156664
rect 366726 156652 366732 156664
rect 353996 156624 366732 156652
rect 353996 156612 354002 156624
rect 366726 156612 366732 156624
rect 366784 156612 366790 156664
rect 85482 155864 85488 155916
rect 85540 155904 85546 155916
rect 90358 155904 90364 155916
rect 85540 155876 90364 155904
rect 85540 155864 85546 155876
rect 90358 155864 90364 155876
rect 90416 155864 90422 155916
rect 86126 154504 86132 154556
rect 86184 154544 86190 154556
rect 91738 154544 91744 154556
rect 86184 154516 91744 154544
rect 86184 154504 86190 154516
rect 91738 154504 91744 154516
rect 91796 154504 91802 154556
rect 170398 153892 170404 153944
rect 170456 153932 170462 153944
rect 172514 153932 172520 153944
rect 170456 153904 172520 153932
rect 170456 153892 170462 153904
rect 172514 153892 172520 153904
rect 172572 153892 172578 153944
rect 71038 153824 71044 153876
rect 71096 153864 71102 153876
rect 100018 153864 100024 153876
rect 71096 153836 100024 153864
rect 71096 153824 71102 153836
rect 100018 153824 100024 153836
rect 100076 153824 100082 153876
rect 373350 153212 373356 153264
rect 373408 153252 373414 153264
rect 375006 153252 375012 153264
rect 373408 153224 375012 153252
rect 373408 153212 373414 153224
rect 375006 153212 375012 153224
rect 375064 153212 375070 153264
rect 154482 152464 154488 152516
rect 154540 152504 154546 152516
rect 169754 152504 169760 152516
rect 154540 152476 169760 152504
rect 154540 152464 154546 152476
rect 169754 152464 169760 152476
rect 169812 152464 169818 152516
rect 97258 152260 97264 152312
rect 97316 152300 97322 152312
rect 103606 152300 103612 152312
rect 97316 152272 103612 152300
rect 97316 152260 97322 152272
rect 103606 152260 103612 152272
rect 103664 152260 103670 152312
rect 180150 151784 180156 151836
rect 180208 151824 180214 151836
rect 580166 151824 580172 151836
rect 180208 151796 580172 151824
rect 180208 151784 180214 151796
rect 580166 151784 580172 151796
rect 580224 151784 580230 151836
rect 102778 151376 102784 151428
rect 102836 151416 102842 151428
rect 104526 151416 104532 151428
rect 102836 151388 104532 151416
rect 102836 151376 102842 151388
rect 104526 151376 104532 151388
rect 104584 151376 104590 151428
rect 172514 150492 172520 150544
rect 172572 150532 172578 150544
rect 176562 150532 176568 150544
rect 172572 150504 176568 150532
rect 172572 150492 172578 150504
rect 176562 150492 176568 150504
rect 176620 150492 176626 150544
rect 103606 149540 103612 149592
rect 103664 149580 103670 149592
rect 109678 149580 109684 149592
rect 103664 149552 109684 149580
rect 103664 149540 103670 149552
rect 109678 149540 109684 149552
rect 109736 149540 109742 149592
rect 3326 149064 3332 149116
rect 3384 149104 3390 149116
rect 24210 149104 24216 149116
rect 3384 149076 24216 149104
rect 3384 149064 3390 149076
rect 24210 149064 24216 149076
rect 24268 149064 24274 149116
rect 104526 148860 104532 148912
rect 104584 148900 104590 148912
rect 106274 148900 106280 148912
rect 104584 148872 106280 148900
rect 104584 148860 104590 148872
rect 106274 148860 106280 148872
rect 106332 148860 106338 148912
rect 339862 146956 339868 147008
rect 339920 146996 339926 147008
rect 353938 146996 353944 147008
rect 339920 146968 353944 146996
rect 339920 146956 339926 146968
rect 353938 146956 353944 146968
rect 353996 146956 354002 147008
rect 118786 146888 118792 146940
rect 118844 146928 118850 146940
rect 580074 146928 580080 146940
rect 118844 146900 580080 146928
rect 118844 146888 118850 146900
rect 580074 146888 580080 146900
rect 580132 146888 580138 146940
rect 176654 146208 176660 146260
rect 176712 146248 176718 146260
rect 178678 146248 178684 146260
rect 176712 146220 178684 146248
rect 176712 146208 176718 146220
rect 178678 146208 178684 146220
rect 178736 146208 178742 146260
rect 371878 146208 371884 146260
rect 371936 146248 371942 146260
rect 373350 146248 373356 146260
rect 371936 146220 373356 146248
rect 371936 146208 371942 146220
rect 373350 146208 373356 146220
rect 373408 146208 373414 146260
rect 157978 145596 157984 145648
rect 158036 145636 158042 145648
rect 164970 145636 164976 145648
rect 158036 145608 164976 145636
rect 158036 145596 158042 145608
rect 164970 145596 164976 145608
rect 165028 145596 165034 145648
rect 119062 145528 119068 145580
rect 119120 145568 119126 145580
rect 477494 145568 477500 145580
rect 119120 145540 477500 145568
rect 119120 145528 119126 145540
rect 477494 145528 477500 145540
rect 477552 145528 477558 145580
rect 69658 144848 69664 144900
rect 69716 144888 69722 144900
rect 71038 144888 71044 144900
rect 69716 144860 71044 144888
rect 69716 144848 69722 144860
rect 71038 144848 71044 144860
rect 71096 144848 71102 144900
rect 335998 144304 336004 144356
rect 336056 144344 336062 144356
rect 339862 144344 339868 144356
rect 336056 144316 339868 144344
rect 336056 144304 336062 144316
rect 339862 144304 339868 144316
rect 339920 144304 339926 144356
rect 343634 144236 343640 144288
rect 343692 144276 343698 144288
rect 348418 144276 348424 144288
rect 343692 144248 348424 144276
rect 343692 144236 343698 144248
rect 348418 144236 348424 144248
rect 348476 144236 348482 144288
rect 118970 144168 118976 144220
rect 119028 144208 119034 144220
rect 580258 144208 580264 144220
rect 119028 144180 580264 144208
rect 119028 144168 119034 144180
rect 580258 144168 580264 144180
rect 580316 144168 580322 144220
rect 79410 143488 79416 143540
rect 79468 143528 79474 143540
rect 80698 143528 80704 143540
rect 79468 143500 80704 143528
rect 79468 143488 79474 143500
rect 80698 143488 80704 143500
rect 80756 143488 80762 143540
rect 164970 143488 164976 143540
rect 165028 143528 165034 143540
rect 168374 143528 168380 143540
rect 165028 143500 168380 143528
rect 165028 143488 165034 143500
rect 168374 143488 168380 143500
rect 168432 143488 168438 143540
rect 24118 143012 24124 143064
rect 24176 143052 24182 143064
rect 182726 143052 182732 143064
rect 24176 143024 182732 143052
rect 24176 143012 24182 143024
rect 182726 143012 182732 143024
rect 182784 143012 182790 143064
rect 20070 142944 20076 142996
rect 20128 142984 20134 142996
rect 182818 142984 182824 142996
rect 20128 142956 182824 142984
rect 20128 142944 20134 142956
rect 182818 142944 182824 142956
rect 182876 142944 182882 142996
rect 6270 142876 6276 142928
rect 6328 142916 6334 142928
rect 182266 142916 182272 142928
rect 6328 142888 182272 142916
rect 6328 142876 6334 142888
rect 182266 142876 182272 142888
rect 182324 142876 182330 142928
rect 118326 142808 118332 142860
rect 118384 142848 118390 142860
rect 398098 142848 398104 142860
rect 118384 142820 398104 142848
rect 118384 142808 118390 142820
rect 398098 142808 398104 142820
rect 398156 142808 398162 142860
rect 106274 142128 106280 142180
rect 106332 142168 106338 142180
rect 106332 142140 107700 142168
rect 106332 142128 106338 142140
rect 107672 142100 107700 142140
rect 330938 142128 330944 142180
rect 330996 142168 331002 142180
rect 335998 142168 336004 142180
rect 330996 142140 336004 142168
rect 330996 142128 331002 142140
rect 335998 142128 336004 142140
rect 336056 142128 336062 142180
rect 109770 142100 109776 142112
rect 107672 142072 109776 142100
rect 109770 142060 109776 142072
rect 109828 142060 109834 142112
rect 40034 141652 40040 141704
rect 40092 141692 40098 141704
rect 181070 141692 181076 141704
rect 40092 141664 181076 141692
rect 40092 141652 40098 141664
rect 181070 141652 181076 141664
rect 181128 141652 181134 141704
rect 19978 141584 19984 141636
rect 20036 141624 20042 141636
rect 182634 141624 182640 141636
rect 20036 141596 182640 141624
rect 20036 141584 20042 141596
rect 182634 141584 182640 141596
rect 182692 141584 182698 141636
rect 326338 141584 326344 141636
rect 326396 141624 326402 141636
rect 343634 141624 343640 141636
rect 326396 141596 343640 141624
rect 326396 141584 326402 141596
rect 343634 141584 343640 141596
rect 343692 141584 343698 141636
rect 118510 141516 118516 141568
rect 118568 141556 118574 141568
rect 398282 141556 398288 141568
rect 118568 141528 398288 141556
rect 118568 141516 118574 141528
rect 398282 141516 398288 141528
rect 398340 141516 398346 141568
rect 118418 141448 118424 141500
rect 118476 141488 118482 141500
rect 398190 141488 398196 141500
rect 118476 141460 398196 141488
rect 118476 141448 118482 141460
rect 398190 141448 398196 141460
rect 398248 141448 398254 141500
rect 119154 141380 119160 141432
rect 119212 141420 119218 141432
rect 580442 141420 580448 141432
rect 119212 141392 580448 141420
rect 119212 141380 119218 141392
rect 580442 141380 580448 141392
rect 580500 141380 580506 141432
rect 369854 140768 369860 140820
rect 369912 140808 369918 140820
rect 371878 140808 371884 140820
rect 369912 140780 371884 140808
rect 369912 140768 369918 140780
rect 371878 140768 371884 140780
rect 371936 140768 371942 140820
rect 140682 140700 140688 140752
rect 140740 140740 140746 140752
rect 142246 140740 142252 140752
rect 140740 140712 142252 140740
rect 140740 140700 140746 140712
rect 142246 140700 142252 140712
rect 142304 140700 142310 140752
rect 90358 140564 90364 140616
rect 90416 140604 90422 140616
rect 94498 140604 94504 140616
rect 90416 140576 94504 140604
rect 90416 140564 90422 140576
rect 94498 140564 94504 140576
rect 94556 140564 94562 140616
rect 150526 140496 150532 140548
rect 150584 140536 150590 140548
rect 154574 140536 154580 140548
rect 150584 140508 154580 140536
rect 150584 140496 150590 140508
rect 154574 140496 154580 140508
rect 154632 140496 154638 140548
rect 163682 140428 163688 140480
rect 163740 140468 163746 140480
rect 174630 140468 174636 140480
rect 163740 140440 174636 140468
rect 163740 140428 163746 140440
rect 174630 140428 174636 140440
rect 174688 140428 174694 140480
rect 164510 140360 164516 140412
rect 164568 140400 164574 140412
rect 176194 140400 176200 140412
rect 164568 140372 176200 140400
rect 164568 140360 164574 140372
rect 176194 140360 176200 140372
rect 176252 140360 176258 140412
rect 144454 140292 144460 140344
rect 144512 140332 144518 140344
rect 160554 140332 160560 140344
rect 144512 140304 160560 140332
rect 144512 140292 144518 140304
rect 160554 140292 160560 140304
rect 160612 140292 160618 140344
rect 163498 140292 163504 140344
rect 163556 140332 163562 140344
rect 178034 140332 178040 140344
rect 163556 140304 178040 140332
rect 163556 140292 163562 140304
rect 178034 140292 178040 140304
rect 178092 140292 178098 140344
rect 142522 140224 142528 140276
rect 142580 140264 142586 140276
rect 173066 140264 173072 140276
rect 142580 140236 173072 140264
rect 142580 140224 142586 140236
rect 173066 140224 173072 140236
rect 173124 140224 173130 140276
rect 119338 140156 119344 140208
rect 119396 140196 119402 140208
rect 412634 140196 412640 140208
rect 119396 140168 412640 140196
rect 119396 140156 119402 140168
rect 412634 140156 412640 140168
rect 412692 140156 412698 140208
rect 120718 140088 120724 140140
rect 120776 140128 120782 140140
rect 542354 140128 542360 140140
rect 120776 140100 542360 140128
rect 120776 140088 120782 140100
rect 542354 140088 542360 140100
rect 542412 140088 542418 140140
rect 118878 140020 118884 140072
rect 118936 140060 118942 140072
rect 580902 140060 580908 140072
rect 118936 140032 580908 140060
rect 118936 140020 118942 140032
rect 580902 140020 580908 140032
rect 580960 140020 580966 140072
rect 178678 139952 178684 140004
rect 178736 139992 178742 140004
rect 179690 139992 179696 140004
rect 178736 139964 179696 139992
rect 178736 139952 178742 139964
rect 179690 139952 179696 139964
rect 179748 139952 179754 140004
rect 123662 139748 123668 139800
rect 123720 139788 123726 139800
rect 124858 139788 124864 139800
rect 123720 139760 124864 139788
rect 123720 139748 123726 139760
rect 124858 139748 124864 139760
rect 124916 139748 124922 139800
rect 146478 139748 146484 139800
rect 146536 139788 146542 139800
rect 148042 139788 148048 139800
rect 146536 139760 148048 139788
rect 146536 139748 146542 139760
rect 148042 139748 148048 139760
rect 148100 139748 148106 139800
rect 153470 139748 153476 139800
rect 153528 139788 153534 139800
rect 158990 139788 158996 139800
rect 153528 139760 158996 139788
rect 153528 139748 153534 139760
rect 158990 139748 158996 139760
rect 159048 139748 159054 139800
rect 137738 139680 137744 139732
rect 137796 139720 137802 139732
rect 139578 139720 139584 139732
rect 137796 139692 139584 139720
rect 137796 139680 137802 139692
rect 139578 139680 139584 139692
rect 139636 139680 139642 139732
rect 147490 139680 147496 139732
rect 147548 139720 147554 139732
rect 149606 139720 149612 139732
rect 147548 139692 149612 139720
rect 147548 139680 147554 139692
rect 149606 139680 149612 139692
rect 149664 139680 149670 139732
rect 152458 139680 152464 139732
rect 152516 139720 152522 139732
rect 157426 139720 157432 139732
rect 152516 139692 157432 139720
rect 152516 139680 152522 139692
rect 157426 139680 157432 139692
rect 157484 139680 157490 139732
rect 149514 139612 149520 139664
rect 149572 139652 149578 139664
rect 152734 139652 152740 139664
rect 149572 139624 152740 139652
rect 149572 139612 149578 139624
rect 152734 139612 152740 139624
rect 152792 139612 152798 139664
rect 120626 138932 120632 138984
rect 120684 138972 120690 138984
rect 158438 138972 158444 138984
rect 120684 138944 158444 138972
rect 120684 138932 120690 138944
rect 158438 138932 158444 138944
rect 158496 138932 158502 138984
rect 100018 138864 100024 138916
rect 100076 138904 100082 138916
rect 182450 138904 182456 138916
rect 100076 138876 182456 138904
rect 100076 138864 100082 138876
rect 182450 138864 182456 138876
rect 182508 138864 182514 138916
rect 3602 138796 3608 138848
rect 3660 138836 3666 138848
rect 179598 138836 179604 138848
rect 3660 138808 179604 138836
rect 3660 138796 3666 138808
rect 179598 138796 179604 138808
rect 179656 138796 179662 138848
rect 3418 138728 3424 138780
rect 3476 138768 3482 138780
rect 182542 138768 182548 138780
rect 3476 138740 182548 138768
rect 3476 138728 3482 138740
rect 182542 138728 182548 138740
rect 182600 138728 182606 138780
rect 320174 138728 320180 138780
rect 320232 138768 320238 138780
rect 330938 138768 330944 138780
rect 320232 138740 330944 138768
rect 320232 138728 320238 138740
rect 330938 138728 330944 138740
rect 330996 138728 331002 138780
rect 119246 138660 119252 138712
rect 119304 138700 119310 138712
rect 580626 138700 580632 138712
rect 119304 138672 580632 138700
rect 119304 138660 119310 138672
rect 580626 138660 580632 138672
rect 580684 138660 580690 138712
rect 117866 137980 117872 138032
rect 117924 138020 117930 138032
rect 580166 138020 580172 138032
rect 117924 137992 580172 138020
rect 117924 137980 117930 137992
rect 580166 137980 580172 137992
rect 580224 137980 580230 138032
rect 179690 137912 179696 137964
rect 179748 137952 179754 137964
rect 181162 137952 181168 137964
rect 179748 137924 181168 137952
rect 179748 137912 179754 137924
rect 181162 137912 181168 137924
rect 181220 137912 181226 137964
rect 366358 137300 366364 137352
rect 366416 137340 366422 137352
rect 369854 137340 369860 137352
rect 366416 137312 369860 137340
rect 366416 137300 366422 137312
rect 369854 137300 369860 137312
rect 369912 137300 369918 137352
rect 46198 137232 46204 137284
rect 46256 137272 46262 137284
rect 117314 137272 117320 137284
rect 46256 137244 117320 137272
rect 46256 137232 46262 137244
rect 117314 137232 117320 137244
rect 117372 137232 117378 137284
rect 119522 137232 119528 137284
rect 119580 137272 119586 137284
rect 359458 137272 359464 137284
rect 119580 137244 359464 137272
rect 119580 137232 119586 137244
rect 359458 137232 359464 137244
rect 359516 137232 359522 137284
rect 318242 136960 318248 137012
rect 318300 137000 318306 137012
rect 320174 137000 320180 137012
rect 318300 136972 320180 137000
rect 318300 136960 318306 136972
rect 320174 136960 320180 136972
rect 320232 136960 320238 137012
rect 3418 136688 3424 136740
rect 3476 136728 3482 136740
rect 116670 136728 116676 136740
rect 3476 136700 116676 136728
rect 3476 136688 3482 136700
rect 116670 136688 116676 136700
rect 116728 136688 116734 136740
rect 19978 136620 19984 136672
rect 20036 136660 20042 136672
rect 182174 136660 182180 136672
rect 20036 136632 182180 136660
rect 20036 136620 20042 136632
rect 182174 136620 182180 136632
rect 182232 136620 182238 136672
rect 94498 136484 94504 136536
rect 94556 136524 94562 136536
rect 100110 136524 100116 136536
rect 94556 136496 100116 136524
rect 94556 136484 94562 136496
rect 100110 136484 100116 136496
rect 100168 136484 100174 136536
rect 306742 135872 306748 135924
rect 306800 135912 306806 135924
rect 318242 135912 318248 135924
rect 306800 135884 318248 135912
rect 306800 135872 306806 135884
rect 318242 135872 318248 135884
rect 318300 135872 318306 135924
rect 91738 134580 91744 134632
rect 91796 134620 91802 134632
rect 94222 134620 94228 134632
rect 91796 134592 94228 134620
rect 91796 134580 91802 134592
rect 94222 134580 94228 134592
rect 94280 134580 94286 134632
rect 3418 133900 3424 133952
rect 3476 133940 3482 133952
rect 117314 133940 117320 133952
rect 3476 133912 117320 133940
rect 3476 133900 3482 133912
rect 117314 133900 117320 133912
rect 117372 133900 117378 133952
rect 304994 133900 305000 133952
rect 305052 133940 305058 133952
rect 306742 133940 306748 133952
rect 305052 133912 306748 133940
rect 305052 133900 305058 133912
rect 306742 133900 306748 133912
rect 306800 133900 306806 133952
rect 3602 132472 3608 132524
rect 3660 132512 3666 132524
rect 117314 132512 117320 132524
rect 3660 132484 117320 132512
rect 3660 132472 3666 132484
rect 117314 132472 117320 132484
rect 117372 132472 117378 132524
rect 71038 131996 71044 132048
rect 71096 132036 71102 132048
rect 72510 132036 72516 132048
rect 71096 132008 72516 132036
rect 71096 131996 71102 132008
rect 72510 131996 72516 132008
rect 72568 131996 72574 132048
rect 100110 131928 100116 131980
rect 100168 131968 100174 131980
rect 105538 131968 105544 131980
rect 100168 131940 105544 131968
rect 100168 131928 100174 131940
rect 105538 131928 105544 131940
rect 105596 131928 105602 131980
rect 94222 131180 94228 131232
rect 94280 131220 94286 131232
rect 99374 131220 99380 131232
rect 94280 131192 99380 131220
rect 94280 131180 94286 131192
rect 99374 131180 99380 131192
rect 99432 131180 99438 131232
rect 3326 131112 3332 131164
rect 3384 131152 3390 131164
rect 117314 131152 117320 131164
rect 3384 131124 117320 131152
rect 3384 131112 3390 131124
rect 117314 131112 117320 131124
rect 117372 131112 117378 131164
rect 361942 129888 361948 129940
rect 362000 129928 362006 129940
rect 366358 129928 366364 129940
rect 362000 129900 366364 129928
rect 362000 129888 362006 129900
rect 366358 129888 366364 129900
rect 366416 129888 366422 129940
rect 24210 129684 24216 129736
rect 24268 129724 24274 129736
rect 117314 129724 117320 129736
rect 24268 129696 117320 129724
rect 24268 129684 24274 129696
rect 117314 129684 117320 129696
rect 117372 129684 117378 129736
rect 300762 128324 300768 128376
rect 300820 128364 300826 128376
rect 304994 128364 305000 128376
rect 300820 128336 305000 128364
rect 300820 128324 300826 128336
rect 304994 128324 305000 128336
rect 305052 128324 305058 128376
rect 22830 128256 22836 128308
rect 22888 128296 22894 128308
rect 117314 128296 117320 128308
rect 22888 128268 117320 128296
rect 22888 128256 22894 128268
rect 117314 128256 117320 128268
rect 117372 128256 117378 128308
rect 22738 126896 22744 126948
rect 22796 126936 22802 126948
rect 117314 126936 117320 126948
rect 22796 126908 117320 126936
rect 22796 126896 22802 126908
rect 117314 126896 117320 126908
rect 117372 126896 117378 126948
rect 99374 126828 99380 126880
rect 99432 126868 99438 126880
rect 106182 126868 106188 126880
rect 99432 126840 106188 126868
rect 99432 126828 99438 126840
rect 106182 126828 106188 126840
rect 106240 126828 106246 126880
rect 314654 126216 314660 126268
rect 314712 126256 314718 126268
rect 326338 126256 326344 126268
rect 314712 126228 326344 126256
rect 314712 126216 314718 126228
rect 326338 126216 326344 126228
rect 326396 126216 326402 126268
rect 184198 125604 184204 125656
rect 184256 125644 184262 125656
rect 580074 125644 580080 125656
rect 184256 125616 580080 125644
rect 184256 125604 184262 125616
rect 580074 125604 580080 125616
rect 580132 125604 580138 125656
rect 72510 125536 72516 125588
rect 72568 125576 72574 125588
rect 73890 125576 73896 125588
rect 72568 125548 73896 125576
rect 72568 125536 72574 125548
rect 73890 125536 73896 125548
rect 73948 125536 73954 125588
rect 6362 124108 6368 124160
rect 6420 124148 6426 124160
rect 117314 124148 117320 124160
rect 6420 124120 117320 124148
rect 6420 124108 6426 124120
rect 117314 124108 117320 124120
rect 117372 124108 117378 124160
rect 118602 124108 118608 124160
rect 118660 124148 118666 124160
rect 119522 124148 119528 124160
rect 118660 124120 119528 124148
rect 118660 124108 118666 124120
rect 119522 124108 119528 124120
rect 119580 124108 119586 124160
rect 312170 123904 312176 123956
rect 312228 123944 312234 123956
rect 314654 123944 314660 123956
rect 312228 123916 314660 123944
rect 312228 123904 312234 123916
rect 314654 123904 314660 123916
rect 314712 123904 314718 123956
rect 360930 123632 360936 123684
rect 360988 123672 360994 123684
rect 361942 123672 361948 123684
rect 360988 123644 361948 123672
rect 360988 123632 360994 123644
rect 361942 123632 361948 123644
rect 362000 123632 362006 123684
rect 106182 123428 106188 123480
rect 106240 123468 106246 123480
rect 115290 123468 115296 123480
rect 106240 123440 115296 123468
rect 106240 123428 106246 123440
rect 115290 123428 115296 123440
rect 115348 123428 115354 123480
rect 295242 123428 295248 123480
rect 295300 123468 295306 123480
rect 300762 123468 300768 123480
rect 295300 123440 300768 123468
rect 295300 123428 295306 123440
rect 300762 123428 300768 123440
rect 300820 123428 300826 123480
rect 10318 122748 10324 122800
rect 10376 122788 10382 122800
rect 117314 122788 117320 122800
rect 10376 122760 117320 122788
rect 10376 122748 10382 122760
rect 117314 122748 117320 122760
rect 117372 122748 117378 122800
rect 73890 122680 73896 122732
rect 73948 122720 73954 122732
rect 75454 122720 75460 122732
rect 73948 122692 75460 122720
rect 73948 122680 73954 122692
rect 75454 122680 75460 122692
rect 75512 122680 75518 122732
rect 109770 121932 109776 121984
rect 109828 121972 109834 121984
rect 111794 121972 111800 121984
rect 109828 121944 111800 121972
rect 109828 121932 109834 121944
rect 111794 121932 111800 121944
rect 111852 121932 111858 121984
rect 8938 121388 8944 121440
rect 8996 121428 9002 121440
rect 117314 121428 117320 121440
rect 8996 121400 117320 121428
rect 8996 121388 9002 121400
rect 117314 121388 117320 121400
rect 117372 121388 117378 121440
rect 80698 120640 80704 120692
rect 80756 120680 80762 120692
rect 82814 120680 82820 120692
rect 80756 120652 82820 120680
rect 80756 120640 80762 120652
rect 82814 120640 82820 120652
rect 82872 120640 82878 120692
rect 4798 120028 4804 120080
rect 4856 120068 4862 120080
rect 117314 120068 117320 120080
rect 4856 120040 117320 120068
rect 4856 120028 4862 120040
rect 117314 120028 117320 120040
rect 117372 120028 117378 120080
rect 105538 119076 105544 119128
rect 105596 119116 105602 119128
rect 109770 119116 109776 119128
rect 105596 119088 109776 119116
rect 105596 119076 105602 119088
rect 109770 119076 109776 119088
rect 109828 119076 109834 119128
rect 43438 118600 43444 118652
rect 43496 118640 43502 118652
rect 117314 118640 117320 118652
rect 43496 118612 117320 118640
rect 43496 118600 43502 118612
rect 117314 118600 117320 118612
rect 117372 118600 117378 118652
rect 82814 118532 82820 118584
rect 82872 118572 82878 118584
rect 86218 118572 86224 118584
rect 82872 118544 86224 118572
rect 82872 118532 82878 118544
rect 86218 118532 86224 118544
rect 86276 118532 86282 118584
rect 79318 118260 79324 118312
rect 79376 118300 79382 118312
rect 81066 118300 81072 118312
rect 79376 118272 81072 118300
rect 79376 118260 79382 118272
rect 81066 118260 81072 118272
rect 81124 118260 81130 118312
rect 307018 117512 307024 117564
rect 307076 117552 307082 117564
rect 312170 117552 312176 117564
rect 307076 117524 312176 117552
rect 307076 117512 307082 117524
rect 312170 117512 312176 117524
rect 312228 117512 312234 117564
rect 358814 117512 358820 117564
rect 358872 117552 358878 117564
rect 360930 117552 360936 117564
rect 358872 117524 360936 117552
rect 358872 117512 358878 117524
rect 360930 117512 360936 117524
rect 360988 117512 360994 117564
rect 292574 117376 292580 117428
rect 292632 117416 292638 117428
rect 295242 117416 295248 117428
rect 292632 117388 295248 117416
rect 292632 117376 292638 117388
rect 295242 117376 295248 117388
rect 295300 117376 295306 117428
rect 15838 117240 15844 117292
rect 15896 117280 15902 117292
rect 117314 117280 117320 117292
rect 15896 117252 117320 117280
rect 15896 117240 15902 117252
rect 117314 117240 117320 117252
rect 117372 117240 117378 117292
rect 111794 117172 111800 117224
rect 111852 117212 111858 117224
rect 115198 117212 115204 117224
rect 111852 117184 115204 117212
rect 111852 117172 111858 117184
rect 115198 117172 115204 117184
rect 115256 117172 115262 117224
rect 6178 115880 6184 115932
rect 6236 115920 6242 115932
rect 117314 115920 117320 115932
rect 6236 115892 117320 115920
rect 6236 115880 6242 115892
rect 117314 115880 117320 115892
rect 117372 115880 117378 115932
rect 354674 115880 354680 115932
rect 354732 115920 354738 115932
rect 358814 115920 358820 115932
rect 354732 115892 358820 115920
rect 354732 115880 354738 115892
rect 358814 115880 358820 115892
rect 358872 115880 358878 115932
rect 81066 115812 81072 115864
rect 81124 115852 81130 115864
rect 82722 115852 82728 115864
rect 81124 115824 82728 115852
rect 81124 115812 81130 115824
rect 82722 115812 82728 115824
rect 82780 115812 82786 115864
rect 118142 114792 118148 114844
rect 118200 114832 118206 114844
rect 119430 114832 119436 114844
rect 118200 114804 119436 114832
rect 118200 114792 118206 114804
rect 119430 114792 119436 114804
rect 119488 114792 119494 114844
rect 75454 114520 75460 114572
rect 75512 114560 75518 114572
rect 75512 114532 75960 114560
rect 75512 114520 75518 114532
rect 75932 114492 75960 114532
rect 81342 114492 81348 114504
rect 75932 114464 81348 114492
rect 81342 114452 81348 114464
rect 81400 114452 81406 114504
rect 291102 114248 291108 114300
rect 291160 114288 291166 114300
rect 292574 114288 292580 114300
rect 291160 114260 292580 114288
rect 291160 114248 291166 114260
rect 292574 114248 292580 114260
rect 292632 114248 292638 114300
rect 33778 113092 33784 113144
rect 33836 113132 33842 113144
rect 117314 113132 117320 113144
rect 33836 113104 117320 113132
rect 33836 113092 33842 113104
rect 117314 113092 117320 113104
rect 117372 113092 117378 113144
rect 86218 112412 86224 112464
rect 86276 112452 86282 112464
rect 87414 112452 87420 112464
rect 86276 112424 87420 112452
rect 86276 112412 86282 112424
rect 87414 112412 87420 112424
rect 87472 112412 87478 112464
rect 180242 111800 180248 111852
rect 180300 111840 180306 111852
rect 580166 111840 580172 111852
rect 180300 111812 580172 111840
rect 180300 111800 180306 111812
rect 580166 111800 580172 111812
rect 580224 111800 580230 111852
rect 3234 111732 3240 111784
rect 3292 111772 3298 111784
rect 19978 111772 19984 111784
rect 3292 111744 19984 111772
rect 3292 111732 3298 111744
rect 19978 111732 19984 111744
rect 20036 111732 20042 111784
rect 115290 111732 115296 111784
rect 115348 111772 115354 111784
rect 117314 111772 117320 111784
rect 115348 111744 117320 111772
rect 115348 111732 115354 111744
rect 117314 111732 117320 111744
rect 117372 111732 117378 111784
rect 303614 111052 303620 111104
rect 303672 111092 303678 111104
rect 307018 111092 307024 111104
rect 303672 111064 307024 111092
rect 303672 111052 303678 111064
rect 307018 111052 307024 111064
rect 307076 111052 307082 111104
rect 81342 110440 81348 110492
rect 81400 110480 81406 110492
rect 81400 110452 84194 110480
rect 81400 110440 81406 110452
rect 84166 110412 84194 110452
rect 117314 110412 117320 110424
rect 84166 110384 117320 110412
rect 117314 110372 117320 110384
rect 117372 110372 117378 110424
rect 87414 109692 87420 109744
rect 87472 109732 87478 109744
rect 97902 109732 97908 109744
rect 87472 109704 97908 109732
rect 87472 109692 87478 109704
rect 97902 109692 97908 109704
rect 97960 109692 97966 109744
rect 97902 108944 97908 108996
rect 97960 108984 97966 108996
rect 117314 108984 117320 108996
rect 97960 108956 117320 108984
rect 97960 108944 97966 108956
rect 117314 108944 117320 108956
rect 117372 108944 117378 108996
rect 183462 108944 183468 108996
rect 183520 108984 183526 108996
rect 354582 108984 354588 108996
rect 183520 108956 354588 108984
rect 183520 108944 183526 108956
rect 354582 108944 354588 108956
rect 354640 108944 354646 108996
rect 291102 107692 291108 107704
rect 289096 107664 291108 107692
rect 82814 107584 82820 107636
rect 82872 107624 82878 107636
rect 117314 107624 117320 107636
rect 82872 107596 117320 107624
rect 82872 107584 82878 107596
rect 117314 107584 117320 107596
rect 117372 107584 117378 107636
rect 183462 107584 183468 107636
rect 183520 107624 183526 107636
rect 289096 107624 289124 107664
rect 291102 107652 291108 107664
rect 291160 107652 291166 107704
rect 183520 107596 289124 107624
rect 183520 107584 183526 107596
rect 109678 107516 109684 107568
rect 109736 107556 109742 107568
rect 112438 107556 112444 107568
rect 109736 107528 112444 107556
rect 109736 107516 109742 107528
rect 112438 107516 112444 107528
rect 112496 107516 112502 107568
rect 183462 106224 183468 106276
rect 183520 106264 183526 106276
rect 410518 106264 410524 106276
rect 183520 106236 410524 106264
rect 183520 106224 183526 106236
rect 410518 106224 410524 106236
rect 410576 106224 410582 106276
rect 291838 105544 291844 105596
rect 291896 105584 291902 105596
rect 303614 105584 303620 105596
rect 291896 105556 303620 105584
rect 291896 105544 291902 105556
rect 303614 105544 303620 105556
rect 303672 105544 303678 105596
rect 183462 104796 183468 104848
rect 183520 104836 183526 104848
rect 409138 104836 409144 104848
rect 183520 104808 409144 104836
rect 183520 104796 183526 104808
rect 409138 104796 409144 104808
rect 409196 104796 409202 104848
rect 183462 103436 183468 103488
rect 183520 103476 183526 103488
rect 407758 103476 407764 103488
rect 183520 103448 407764 103476
rect 183520 103436 183526 103448
rect 407758 103436 407764 103448
rect 407816 103436 407822 103488
rect 183462 102076 183468 102128
rect 183520 102116 183526 102128
rect 544378 102116 544384 102128
rect 183520 102088 544384 102116
rect 183520 102076 183526 102088
rect 544378 102076 544384 102088
rect 544436 102076 544442 102128
rect 109770 102008 109776 102060
rect 109828 102048 109834 102060
rect 115842 102048 115848 102060
rect 109828 102020 115848 102048
rect 109828 102008 109834 102020
rect 115842 102008 115848 102020
rect 115900 102008 115906 102060
rect 182818 100648 182824 100700
rect 182876 100688 182882 100700
rect 406378 100688 406384 100700
rect 182876 100660 406384 100688
rect 182876 100648 182882 100660
rect 406378 100648 406384 100660
rect 406436 100648 406442 100700
rect 180334 99356 180340 99408
rect 180392 99396 180398 99408
rect 580166 99396 580172 99408
rect 180392 99368 580172 99396
rect 180392 99356 180398 99368
rect 580166 99356 580172 99368
rect 580224 99356 580230 99408
rect 182818 99288 182824 99340
rect 182876 99328 182882 99340
rect 404998 99328 405004 99340
rect 182876 99300 405004 99328
rect 182876 99288 182882 99300
rect 404998 99288 405004 99300
rect 405056 99288 405062 99340
rect 117958 98676 117964 98728
rect 118016 98716 118022 98728
rect 120902 98716 120908 98728
rect 118016 98688 120908 98716
rect 118016 98676 118022 98688
rect 120902 98676 120908 98688
rect 120960 98676 120966 98728
rect 115198 97928 115204 97980
rect 115256 97968 115262 97980
rect 116762 97968 116768 97980
rect 115256 97940 116768 97968
rect 115256 97928 115262 97940
rect 116762 97928 116768 97940
rect 116820 97928 116826 97980
rect 183462 97928 183468 97980
rect 183520 97968 183526 97980
rect 403618 97968 403624 97980
rect 183520 97940 403624 97968
rect 183520 97928 183526 97940
rect 403618 97928 403624 97940
rect 403676 97928 403682 97980
rect 115842 95140 115848 95192
rect 115900 95180 115906 95192
rect 120810 95180 120816 95192
rect 115900 95152 120816 95180
rect 115900 95140 115906 95152
rect 120810 95140 120816 95152
rect 120868 95140 120874 95192
rect 183462 95140 183468 95192
rect 183520 95180 183526 95192
rect 400858 95180 400864 95192
rect 183520 95152 400864 95180
rect 183520 95140 183526 95152
rect 400858 95140 400864 95152
rect 400916 95140 400922 95192
rect 183462 93780 183468 93832
rect 183520 93820 183526 93832
rect 418798 93820 418804 93832
rect 183520 93792 418804 93820
rect 183520 93780 183526 93792
rect 418798 93780 418804 93792
rect 418856 93780 418862 93832
rect 183462 92420 183468 92472
rect 183520 92460 183526 92472
rect 417418 92460 417424 92472
rect 183520 92432 417424 92460
rect 183520 92420 183526 92432
rect 417418 92420 417424 92432
rect 417476 92420 417482 92472
rect 183462 90992 183468 91044
rect 183520 91032 183526 91044
rect 414658 91032 414664 91044
rect 183520 91004 414664 91032
rect 183520 90992 183526 91004
rect 414658 90992 414664 91004
rect 414716 90992 414722 91044
rect 182266 89632 182272 89684
rect 182324 89672 182330 89684
rect 413278 89672 413284 89684
rect 182324 89644 413284 89672
rect 182324 89632 182330 89644
rect 413278 89632 413284 89644
rect 413336 89632 413342 89684
rect 116762 88952 116768 89004
rect 116820 88992 116826 89004
rect 117958 88992 117964 89004
rect 116820 88964 117964 88992
rect 116820 88952 116826 88964
rect 117958 88952 117964 88964
rect 118016 88952 118022 89004
rect 183462 88136 183468 88188
rect 183520 88176 183526 88188
rect 189718 88176 189724 88188
rect 183520 88148 189724 88176
rect 183520 88136 183526 88148
rect 189718 88136 189724 88148
rect 189776 88136 189782 88188
rect 284938 87592 284944 87644
rect 284996 87632 285002 87644
rect 291838 87632 291844 87644
rect 284996 87604 291844 87632
rect 284996 87592 285002 87604
rect 291838 87592 291844 87604
rect 291896 87592 291902 87644
rect 183462 86844 183468 86896
rect 183520 86884 183526 86896
rect 188338 86884 188344 86896
rect 183520 86856 188344 86884
rect 183520 86844 183526 86856
rect 188338 86844 188344 86856
rect 188396 86844 188402 86896
rect 182266 85552 182272 85604
rect 182324 85592 182330 85604
rect 580166 85592 580172 85604
rect 182324 85564 580172 85592
rect 182324 85552 182330 85564
rect 580166 85552 580172 85564
rect 580224 85552 580230 85604
rect 182174 85484 182180 85536
rect 182232 85524 182238 85536
rect 184198 85524 184204 85536
rect 182232 85496 184204 85524
rect 182232 85484 182238 85496
rect 184198 85484 184204 85496
rect 184256 85484 184262 85536
rect 120902 85008 120908 85060
rect 120960 85008 120966 85060
rect 120920 84856 120948 85008
rect 120902 84804 120908 84856
rect 120960 84804 120966 84856
rect 3142 84192 3148 84244
rect 3200 84232 3206 84244
rect 120718 84232 120724 84244
rect 3200 84204 120724 84232
rect 3200 84192 3206 84204
rect 120718 84192 120724 84204
rect 120776 84192 120782 84244
rect 117958 81404 117964 81456
rect 118016 81444 118022 81456
rect 118016 81416 118694 81444
rect 118016 81404 118022 81416
rect 118666 81376 118694 81416
rect 120810 81376 120816 81388
rect 118666 81348 120816 81376
rect 120810 81336 120816 81348
rect 120868 81336 120874 81388
rect 183462 80044 183468 80096
rect 183520 80084 183526 80096
rect 555418 80084 555424 80096
rect 183520 80056 555424 80084
rect 183520 80044 183526 80056
rect 555418 80044 555424 80056
rect 555476 80044 555482 80096
rect 178954 79296 178960 79348
rect 179012 79336 179018 79348
rect 580534 79336 580540 79348
rect 179012 79308 580540 79336
rect 179012 79296 179018 79308
rect 580534 79296 580540 79308
rect 580592 79296 580598 79348
rect 180334 78724 180340 78736
rect 154546 78696 166994 78724
rect 120626 78616 120632 78668
rect 120684 78656 120690 78668
rect 124766 78656 124772 78668
rect 120684 78628 124772 78656
rect 120684 78616 120690 78628
rect 124766 78616 124772 78628
rect 124824 78616 124830 78668
rect 133846 78628 144822 78656
rect 124950 78548 124956 78600
rect 125008 78588 125014 78600
rect 133846 78588 133874 78628
rect 125008 78560 133874 78588
rect 125008 78548 125014 78560
rect 4890 78480 4896 78532
rect 4948 78520 4954 78532
rect 4948 78492 144730 78520
rect 4948 78480 4954 78492
rect 133846 78424 144638 78452
rect 4062 78344 4068 78396
rect 4120 78384 4126 78396
rect 133846 78384 133874 78424
rect 4120 78356 124214 78384
rect 4120 78344 4126 78356
rect 124186 78316 124214 78356
rect 126210 78356 133874 78384
rect 134030 78356 143626 78384
rect 126210 78316 126238 78356
rect 134030 78316 134058 78356
rect 124186 78288 126238 78316
rect 130488 78288 134058 78316
rect 3878 78208 3884 78260
rect 3936 78248 3942 78260
rect 118786 78248 118792 78260
rect 3936 78220 118792 78248
rect 3936 78208 3942 78220
rect 118786 78208 118792 78220
rect 118844 78208 118850 78260
rect 122098 78072 122104 78124
rect 122156 78112 122162 78124
rect 122156 78084 127434 78112
rect 122156 78072 122162 78084
rect 124858 78004 124864 78056
rect 124916 78044 124922 78056
rect 124916 78016 127066 78044
rect 124916 78004 124922 78016
rect 112438 77936 112444 77988
rect 112496 77976 112502 77988
rect 124766 77976 124772 77988
rect 112496 77948 124772 77976
rect 112496 77936 112502 77948
rect 124766 77936 124772 77948
rect 124824 77936 124830 77988
rect 127038 77920 127066 78016
rect 125318 77868 125324 77920
rect 125376 77908 125382 77920
rect 125824 77908 125830 77920
rect 125376 77880 125830 77908
rect 125376 77868 125382 77880
rect 125824 77868 125830 77880
rect 125882 77868 125888 77920
rect 126928 77908 126934 77920
rect 126854 77880 126934 77908
rect 121638 77800 121644 77852
rect 121696 77840 121702 77852
rect 126100 77840 126106 77852
rect 121696 77812 126106 77840
rect 121696 77800 121702 77812
rect 126100 77800 126106 77812
rect 126158 77800 126164 77852
rect 126192 77800 126198 77852
rect 126250 77800 126256 77852
rect 126376 77840 126382 77852
rect 126348 77800 126382 77840
rect 126434 77800 126440 77852
rect 126210 77716 126238 77800
rect 126348 77716 126376 77800
rect 126146 77664 126152 77716
rect 126204 77676 126238 77716
rect 126204 77664 126210 77676
rect 126330 77664 126336 77716
rect 126388 77664 126394 77716
rect 126652 77664 126658 77716
rect 126710 77664 126716 77716
rect 119798 77596 119804 77648
rect 119856 77636 119862 77648
rect 119856 77608 122834 77636
rect 119856 77596 119862 77608
rect 122806 77364 122834 77608
rect 125042 77460 125048 77512
rect 125100 77500 125106 77512
rect 126670 77500 126698 77664
rect 125100 77472 126698 77500
rect 125100 77460 125106 77472
rect 125870 77392 125876 77444
rect 125928 77432 125934 77444
rect 126854 77432 126882 77880
rect 126928 77868 126934 77880
rect 126986 77868 126992 77920
rect 127020 77868 127026 77920
rect 127078 77868 127084 77920
rect 127112 77868 127118 77920
rect 127170 77868 127176 77920
rect 127204 77868 127210 77920
rect 127262 77868 127268 77920
rect 127130 77784 127158 77868
rect 127066 77732 127072 77784
rect 127124 77744 127158 77784
rect 127124 77732 127130 77744
rect 126974 77664 126980 77716
rect 127032 77704 127038 77716
rect 127222 77704 127250 77868
rect 127406 77852 127434 78084
rect 128418 77948 129458 77976
rect 127480 77868 127486 77920
rect 127538 77868 127544 77920
rect 127664 77868 127670 77920
rect 127722 77868 127728 77920
rect 127756 77868 127762 77920
rect 127814 77868 127820 77920
rect 127848 77868 127854 77920
rect 127906 77868 127912 77920
rect 127940 77868 127946 77920
rect 127998 77908 128004 77920
rect 127998 77868 128032 77908
rect 128124 77868 128130 77920
rect 128182 77868 128188 77920
rect 128216 77868 128222 77920
rect 128274 77868 128280 77920
rect 128308 77868 128314 77920
rect 128366 77868 128372 77920
rect 127296 77800 127302 77852
rect 127354 77800 127360 77852
rect 127388 77800 127394 77852
rect 127446 77800 127452 77852
rect 127032 77676 127250 77704
rect 127032 77664 127038 77676
rect 127314 77648 127342 77800
rect 127498 77648 127526 77868
rect 127682 77716 127710 77868
rect 127774 77784 127802 77868
rect 127866 77840 127894 77868
rect 127866 77812 127940 77840
rect 127912 77784 127940 77812
rect 127774 77744 127808 77784
rect 127802 77732 127808 77744
rect 127860 77732 127866 77784
rect 127894 77732 127900 77784
rect 127952 77732 127958 77784
rect 128004 77716 128032 77868
rect 128142 77716 128170 77868
rect 127618 77664 127624 77716
rect 127676 77676 127710 77716
rect 127676 77664 127682 77676
rect 127986 77664 127992 77716
rect 128044 77664 128050 77716
rect 128078 77664 128084 77716
rect 128136 77676 128170 77716
rect 128136 77664 128142 77676
rect 127250 77596 127256 77648
rect 127308 77608 127342 77648
rect 127308 77596 127314 77608
rect 127434 77596 127440 77648
rect 127492 77608 127526 77648
rect 127492 77596 127498 77608
rect 128234 77568 128262 77868
rect 128326 77716 128354 77868
rect 128308 77664 128314 77716
rect 128366 77664 128372 77716
rect 127498 77540 128262 77568
rect 125928 77404 126882 77432
rect 125928 77392 125934 77404
rect 127342 77392 127348 77444
rect 127400 77432 127406 77444
rect 127498 77432 127526 77540
rect 127710 77460 127716 77512
rect 127768 77500 127774 77512
rect 128418 77500 128446 77948
rect 129430 77920 129458 77948
rect 128492 77868 128498 77920
rect 128550 77868 128556 77920
rect 128584 77868 128590 77920
rect 128642 77868 128648 77920
rect 128676 77868 128682 77920
rect 128734 77868 128740 77920
rect 129136 77868 129142 77920
rect 129194 77868 129200 77920
rect 129320 77868 129326 77920
rect 129378 77868 129384 77920
rect 129412 77868 129418 77920
rect 129470 77868 129476 77920
rect 129504 77868 129510 77920
rect 129562 77868 129568 77920
rect 129596 77868 129602 77920
rect 129654 77868 129660 77920
rect 129964 77908 129970 77920
rect 129752 77880 129970 77908
rect 128510 77580 128538 77868
rect 128602 77636 128630 77868
rect 128694 77704 128722 77868
rect 129154 77772 129182 77868
rect 129228 77800 129234 77852
rect 129286 77800 129292 77852
rect 129016 77744 129182 77772
rect 128694 77676 128860 77704
rect 128602 77608 128676 77636
rect 128648 77580 128676 77608
rect 128510 77540 128544 77580
rect 128538 77528 128544 77540
rect 128596 77528 128602 77580
rect 128630 77528 128636 77580
rect 128688 77528 128694 77580
rect 128832 77512 128860 77676
rect 129016 77636 129044 77744
rect 129090 77664 129096 77716
rect 129148 77704 129154 77716
rect 129246 77704 129274 77800
rect 129148 77676 129274 77704
rect 129338 77716 129366 77868
rect 129522 77784 129550 77868
rect 129458 77732 129464 77784
rect 129516 77744 129550 77784
rect 129516 77732 129522 77744
rect 129614 77716 129642 77868
rect 129338 77676 129372 77716
rect 129148 77664 129154 77676
rect 129366 77664 129372 77676
rect 129424 77664 129430 77716
rect 129550 77664 129556 77716
rect 129608 77676 129642 77716
rect 129608 77664 129614 77676
rect 129182 77636 129188 77648
rect 129016 77608 129188 77636
rect 129182 77596 129188 77608
rect 129240 77596 129246 77648
rect 129752 77568 129780 77880
rect 129964 77868 129970 77880
rect 130022 77868 130028 77920
rect 130148 77868 130154 77920
rect 130206 77868 130212 77920
rect 130240 77868 130246 77920
rect 130298 77868 130304 77920
rect 129918 77732 129924 77784
rect 129976 77772 129982 77784
rect 130166 77772 130194 77868
rect 129976 77744 130194 77772
rect 129976 77732 129982 77744
rect 130258 77716 130286 77868
rect 130194 77664 130200 77716
rect 130252 77676 130286 77716
rect 130252 77664 130258 77676
rect 130010 77568 130016 77580
rect 129752 77540 130016 77568
rect 130010 77528 130016 77540
rect 130068 77528 130074 77580
rect 127768 77472 128446 77500
rect 127768 77460 127774 77472
rect 128814 77460 128820 77512
rect 128872 77460 128878 77512
rect 127400 77404 127526 77432
rect 127400 77392 127406 77404
rect 129274 77392 129280 77444
rect 129332 77432 129338 77444
rect 130488 77432 130516 78288
rect 143598 78180 143626 78356
rect 143598 78152 143764 78180
rect 142080 78016 142522 78044
rect 136376 77948 136634 77976
rect 130608 77908 130614 77920
rect 130580 77868 130614 77908
rect 130666 77868 130672 77920
rect 130700 77868 130706 77920
rect 130758 77868 130764 77920
rect 130792 77868 130798 77920
rect 130850 77868 130856 77920
rect 130976 77868 130982 77920
rect 131034 77868 131040 77920
rect 131160 77868 131166 77920
rect 131218 77868 131224 77920
rect 131252 77868 131258 77920
rect 131310 77868 131316 77920
rect 131436 77868 131442 77920
rect 131494 77868 131500 77920
rect 131528 77868 131534 77920
rect 131586 77868 131592 77920
rect 131804 77868 131810 77920
rect 131862 77868 131868 77920
rect 131896 77868 131902 77920
rect 131954 77908 131960 77920
rect 132172 77908 132178 77920
rect 131954 77880 132080 77908
rect 131954 77868 131960 77880
rect 130580 77636 130608 77868
rect 130718 77840 130746 77868
rect 130672 77812 130746 77840
rect 130672 77784 130700 77812
rect 130810 77784 130838 77868
rect 130654 77732 130660 77784
rect 130712 77732 130718 77784
rect 130746 77732 130752 77784
rect 130804 77744 130838 77784
rect 130804 77732 130810 77744
rect 130994 77648 131022 77868
rect 131178 77840 131206 77868
rect 131132 77812 131206 77840
rect 131132 77648 131160 77812
rect 131270 77784 131298 77868
rect 131206 77732 131212 77784
rect 131264 77744 131298 77784
rect 131264 77732 131270 77744
rect 130838 77636 130844 77648
rect 130580 77608 130844 77636
rect 130838 77596 130844 77608
rect 130896 77596 130902 77648
rect 130930 77596 130936 77648
rect 130988 77608 131022 77648
rect 130988 77596 130994 77608
rect 131114 77596 131120 77648
rect 131172 77596 131178 77648
rect 129332 77404 130516 77432
rect 131454 77432 131482 77868
rect 131546 77648 131574 77868
rect 131822 77840 131850 77868
rect 131822 77812 131988 77840
rect 131546 77608 131580 77648
rect 131574 77596 131580 77608
rect 131632 77596 131638 77648
rect 131666 77528 131672 77580
rect 131724 77568 131730 77580
rect 131960 77568 131988 77812
rect 131724 77540 131988 77568
rect 131724 77528 131730 77540
rect 131758 77460 131764 77512
rect 131816 77500 131822 77512
rect 132052 77500 132080 77880
rect 132144 77868 132178 77908
rect 132230 77868 132236 77920
rect 132264 77868 132270 77920
rect 132322 77868 132328 77920
rect 132448 77868 132454 77920
rect 132506 77868 132512 77920
rect 132632 77908 132638 77920
rect 132604 77868 132638 77908
rect 132690 77868 132696 77920
rect 132724 77868 132730 77920
rect 132782 77868 132788 77920
rect 133092 77868 133098 77920
rect 133150 77868 133156 77920
rect 133368 77868 133374 77920
rect 133426 77868 133432 77920
rect 133460 77868 133466 77920
rect 133518 77868 133524 77920
rect 133552 77868 133558 77920
rect 133610 77868 133616 77920
rect 133736 77868 133742 77920
rect 133794 77868 133800 77920
rect 133920 77868 133926 77920
rect 133978 77868 133984 77920
rect 134012 77868 134018 77920
rect 134070 77868 134076 77920
rect 134104 77868 134110 77920
rect 134162 77868 134168 77920
rect 134196 77868 134202 77920
rect 134254 77868 134260 77920
rect 134472 77868 134478 77920
rect 134530 77868 134536 77920
rect 134564 77868 134570 77920
rect 134622 77908 134628 77920
rect 134622 77880 134748 77908
rect 134622 77868 134628 77880
rect 132144 77568 132172 77868
rect 132282 77840 132310 77868
rect 132236 77812 132310 77840
rect 132236 77648 132264 77812
rect 132310 77664 132316 77716
rect 132368 77704 132374 77716
rect 132466 77704 132494 77868
rect 132604 77784 132632 77868
rect 132742 77840 132770 77868
rect 132696 77812 132770 77840
rect 132586 77732 132592 77784
rect 132644 77732 132650 77784
rect 132368 77676 132494 77704
rect 132368 77664 132374 77676
rect 132696 77648 132724 77812
rect 132816 77772 132822 77784
rect 132788 77732 132822 77772
rect 132874 77732 132880 77784
rect 132218 77596 132224 77648
rect 132276 77596 132282 77648
rect 132678 77596 132684 77648
rect 132736 77596 132742 77648
rect 132402 77568 132408 77580
rect 132144 77540 132408 77568
rect 132402 77528 132408 77540
rect 132460 77528 132466 77580
rect 132788 77568 132816 77732
rect 133110 77636 133138 77868
rect 133230 77636 133236 77648
rect 133110 77608 133236 77636
rect 133230 77596 133236 77608
rect 133288 77596 133294 77648
rect 133046 77568 133052 77580
rect 132788 77540 133052 77568
rect 133046 77528 133052 77540
rect 133104 77528 133110 77580
rect 133138 77528 133144 77580
rect 133196 77568 133202 77580
rect 133386 77568 133414 77868
rect 133196 77540 133414 77568
rect 133196 77528 133202 77540
rect 133478 77512 133506 77868
rect 131816 77472 132080 77500
rect 131816 77460 131822 77472
rect 133414 77460 133420 77512
rect 133472 77472 133506 77512
rect 133472 77460 133478 77472
rect 133570 77444 133598 77868
rect 133754 77580 133782 77868
rect 133938 77784 133966 77868
rect 133874 77732 133880 77784
rect 133932 77744 133966 77784
rect 133932 77732 133938 77744
rect 134030 77704 134058 77868
rect 133690 77528 133696 77580
rect 133748 77540 133782 77580
rect 133984 77676 134058 77704
rect 133984 77568 134012 77676
rect 134122 77648 134150 77868
rect 134058 77596 134064 77648
rect 134116 77608 134150 77648
rect 134214 77636 134242 77868
rect 134490 77784 134518 77868
rect 134426 77732 134432 77784
rect 134484 77744 134518 77784
rect 134484 77732 134490 77744
rect 134214 77608 134472 77636
rect 134116 77596 134122 77608
rect 134334 77568 134340 77580
rect 133984 77540 134340 77568
rect 133748 77528 133754 77540
rect 134334 77528 134340 77540
rect 134392 77528 134398 77580
rect 133966 77460 133972 77512
rect 134024 77500 134030 77512
rect 134444 77500 134472 77608
rect 134720 77580 134748 77880
rect 134840 77868 134846 77920
rect 134898 77868 134904 77920
rect 134932 77868 134938 77920
rect 134990 77868 134996 77920
rect 135024 77868 135030 77920
rect 135082 77868 135088 77920
rect 135208 77868 135214 77920
rect 135266 77868 135272 77920
rect 135300 77868 135306 77920
rect 135358 77868 135364 77920
rect 135484 77868 135490 77920
rect 135542 77868 135548 77920
rect 135576 77868 135582 77920
rect 135634 77868 135640 77920
rect 135668 77868 135674 77920
rect 135726 77868 135732 77920
rect 135852 77868 135858 77920
rect 135910 77868 135916 77920
rect 135944 77868 135950 77920
rect 136002 77868 136008 77920
rect 134858 77840 134886 77868
rect 134812 77812 134886 77840
rect 134812 77716 134840 77812
rect 134950 77772 134978 77868
rect 134904 77744 134978 77772
rect 134904 77716 134932 77744
rect 135042 77716 135070 77868
rect 134794 77664 134800 77716
rect 134852 77664 134858 77716
rect 134886 77664 134892 77716
rect 134944 77664 134950 77716
rect 134978 77664 134984 77716
rect 135036 77676 135070 77716
rect 135226 77716 135254 77868
rect 135318 77772 135346 77868
rect 135502 77840 135530 77868
rect 135456 77812 135530 77840
rect 135318 77744 135392 77772
rect 135226 77676 135260 77716
rect 135036 77664 135042 77676
rect 135254 77664 135260 77676
rect 135312 77664 135318 77716
rect 135364 77648 135392 77744
rect 135456 77648 135484 77812
rect 135594 77772 135622 77868
rect 135548 77744 135622 77772
rect 135346 77596 135352 77648
rect 135404 77596 135410 77648
rect 135438 77596 135444 77648
rect 135496 77596 135502 77648
rect 134702 77528 134708 77580
rect 134760 77528 134766 77580
rect 135548 77512 135576 77744
rect 135686 77716 135714 77868
rect 135622 77664 135628 77716
rect 135680 77676 135714 77716
rect 135680 77664 135686 77676
rect 135870 77648 135898 77868
rect 135962 77704 135990 77868
rect 136128 77800 136134 77852
rect 136186 77840 136192 77852
rect 136186 77812 136312 77840
rect 136186 77800 136192 77812
rect 136082 77704 136088 77716
rect 135962 77676 136088 77704
rect 136082 77664 136088 77676
rect 136140 77664 136146 77716
rect 136284 77648 136312 77812
rect 135870 77608 135904 77648
rect 135898 77596 135904 77608
rect 135956 77596 135962 77648
rect 136266 77596 136272 77648
rect 136324 77596 136330 77648
rect 135990 77528 135996 77580
rect 136048 77568 136054 77580
rect 136376 77568 136404 77948
rect 136496 77868 136502 77920
rect 136554 77868 136560 77920
rect 136048 77540 136404 77568
rect 136514 77580 136542 77868
rect 136606 77852 136634 77948
rect 137710 77948 138014 77976
rect 136772 77868 136778 77920
rect 136830 77868 136836 77920
rect 137324 77908 137330 77920
rect 136928 77880 137330 77908
rect 136588 77800 136594 77852
rect 136646 77800 136652 77852
rect 136790 77716 136818 77868
rect 136726 77664 136732 77716
rect 136784 77676 136818 77716
rect 136784 77664 136790 77676
rect 136634 77596 136640 77648
rect 136692 77636 136698 77648
rect 136928 77636 136956 77880
rect 137324 77868 137330 77880
rect 137382 77868 137388 77920
rect 137508 77868 137514 77920
rect 137566 77868 137572 77920
rect 137600 77868 137606 77920
rect 137658 77868 137664 77920
rect 137048 77800 137054 77852
rect 137106 77800 137112 77852
rect 136692 77608 136956 77636
rect 136692 77596 136698 77608
rect 136514 77540 136548 77580
rect 136048 77528 136054 77540
rect 136542 77528 136548 77540
rect 136600 77528 136606 77580
rect 136910 77528 136916 77580
rect 136968 77568 136974 77580
rect 137066 77568 137094 77800
rect 137526 77716 137554 77868
rect 137462 77664 137468 77716
rect 137520 77676 137554 77716
rect 137520 77664 137526 77676
rect 136968 77540 137094 77568
rect 137618 77580 137646 77868
rect 137710 77704 137738 77948
rect 137986 77920 138014 77948
rect 138538 77948 139118 77976
rect 138538 77920 138566 77948
rect 137784 77868 137790 77920
rect 137842 77868 137848 77920
rect 137876 77868 137882 77920
rect 137934 77868 137940 77920
rect 137968 77868 137974 77920
rect 138026 77868 138032 77920
rect 138152 77868 138158 77920
rect 138210 77868 138216 77920
rect 138244 77868 138250 77920
rect 138302 77868 138308 77920
rect 138336 77868 138342 77920
rect 138394 77908 138400 77920
rect 138394 77868 138428 77908
rect 138520 77868 138526 77920
rect 138578 77868 138584 77920
rect 138612 77868 138618 77920
rect 138670 77868 138676 77920
rect 138796 77868 138802 77920
rect 138854 77868 138860 77920
rect 138980 77868 138986 77920
rect 139038 77868 139044 77920
rect 137802 77784 137830 77868
rect 137894 77840 137922 77868
rect 137894 77812 138060 77840
rect 137802 77744 137836 77784
rect 137830 77732 137836 77744
rect 137888 77732 137894 77784
rect 137922 77704 137928 77716
rect 137710 77676 137928 77704
rect 137922 77664 137928 77676
rect 137980 77664 137986 77716
rect 137618 77540 137652 77580
rect 136968 77528 136974 77540
rect 137646 77528 137652 77540
rect 137704 77528 137710 77580
rect 138032 77568 138060 77812
rect 138170 77716 138198 77868
rect 138262 77784 138290 77868
rect 138262 77744 138296 77784
rect 138290 77732 138296 77744
rect 138348 77732 138354 77784
rect 138170 77676 138204 77716
rect 138198 77664 138204 77676
rect 138256 77664 138262 77716
rect 138106 77568 138112 77580
rect 138032 77540 138112 77568
rect 138106 77528 138112 77540
rect 138164 77528 138170 77580
rect 138400 77568 138428 77868
rect 138630 77704 138658 77868
rect 138630 77676 138704 77704
rect 138262 77540 138428 77568
rect 134024 77472 134472 77500
rect 134024 77460 134030 77472
rect 135530 77460 135536 77512
rect 135588 77460 135594 77512
rect 131850 77432 131856 77444
rect 131454 77404 131856 77432
rect 129332 77392 129338 77404
rect 131850 77392 131856 77404
rect 131908 77392 131914 77444
rect 133506 77392 133512 77444
rect 133564 77404 133598 77444
rect 138262 77432 138290 77540
rect 138676 77444 138704 77676
rect 138814 77648 138842 77868
rect 138998 77704 139026 77868
rect 138952 77676 139026 77704
rect 138952 77648 138980 77676
rect 138814 77608 138848 77648
rect 138842 77596 138848 77608
rect 138900 77596 138906 77648
rect 138934 77596 138940 77648
rect 138992 77596 138998 77648
rect 138750 77528 138756 77580
rect 138808 77568 138814 77580
rect 139090 77568 139118 77948
rect 140930 77948 141142 77976
rect 139164 77868 139170 77920
rect 139222 77868 139228 77920
rect 139348 77908 139354 77920
rect 139320 77868 139354 77908
rect 139406 77868 139412 77920
rect 139440 77868 139446 77920
rect 139498 77868 139504 77920
rect 139532 77868 139538 77920
rect 139590 77868 139596 77920
rect 139624 77868 139630 77920
rect 139682 77868 139688 77920
rect 139716 77868 139722 77920
rect 139774 77868 139780 77920
rect 140176 77868 140182 77920
rect 140234 77868 140240 77920
rect 140360 77868 140366 77920
rect 140418 77868 140424 77920
rect 140728 77908 140734 77920
rect 140700 77868 140734 77908
rect 140786 77868 140792 77920
rect 140820 77868 140826 77920
rect 140878 77868 140884 77920
rect 138808 77540 139118 77568
rect 138808 77528 138814 77540
rect 139026 77460 139032 77512
rect 139084 77500 139090 77512
rect 139182 77500 139210 77868
rect 139320 77648 139348 77868
rect 139458 77840 139486 77868
rect 139412 77812 139486 77840
rect 139412 77648 139440 77812
rect 139550 77716 139578 77868
rect 139486 77664 139492 77716
rect 139544 77676 139578 77716
rect 139544 77664 139550 77676
rect 139302 77596 139308 77648
rect 139360 77596 139366 77648
rect 139394 77596 139400 77648
rect 139452 77596 139458 77648
rect 139084 77472 139210 77500
rect 139642 77500 139670 77868
rect 139734 77568 139762 77868
rect 140194 77648 140222 77868
rect 140378 77648 140406 77868
rect 140544 77800 140550 77852
rect 140602 77800 140608 77852
rect 140194 77608 140228 77648
rect 140222 77596 140228 77608
rect 140280 77596 140286 77648
rect 140378 77608 140412 77648
rect 140406 77596 140412 77608
rect 140464 77596 140470 77648
rect 139946 77568 139952 77580
rect 139734 77540 139952 77568
rect 139946 77528 139952 77540
rect 140004 77528 140010 77580
rect 139762 77500 139768 77512
rect 139642 77472 139768 77500
rect 139084 77460 139090 77472
rect 139762 77460 139768 77472
rect 139820 77460 139826 77512
rect 139854 77460 139860 77512
rect 139912 77500 139918 77512
rect 140562 77500 140590 77800
rect 140700 77648 140728 77868
rect 140838 77840 140866 77868
rect 140792 77812 140866 77840
rect 140792 77716 140820 77812
rect 140774 77664 140780 77716
rect 140832 77664 140838 77716
rect 140682 77596 140688 77648
rect 140740 77596 140746 77648
rect 139912 77472 140590 77500
rect 139912 77460 139918 77472
rect 138032 77404 138290 77432
rect 133564 77392 133570 77404
rect 126698 77364 126704 77376
rect 122806 77336 126704 77364
rect 126698 77324 126704 77336
rect 126756 77324 126762 77376
rect 128372 77336 129228 77364
rect 118786 77188 118792 77240
rect 118844 77228 118850 77240
rect 128372 77228 128400 77336
rect 129200 77296 129228 77336
rect 130562 77324 130568 77376
rect 130620 77364 130626 77376
rect 130746 77364 130752 77376
rect 130620 77336 130752 77364
rect 130620 77324 130626 77336
rect 130746 77324 130752 77336
rect 130804 77324 130810 77376
rect 134150 77296 134156 77308
rect 129200 77268 134156 77296
rect 134150 77256 134156 77268
rect 134208 77256 134214 77308
rect 118844 77200 128400 77228
rect 138032 77228 138060 77404
rect 138658 77392 138664 77444
rect 138716 77392 138722 77444
rect 138566 77324 138572 77376
rect 138624 77364 138630 77376
rect 139578 77364 139584 77376
rect 138624 77336 139584 77364
rect 138624 77324 138630 77336
rect 139578 77324 139584 77336
rect 139636 77324 139642 77376
rect 140930 77364 140958 77948
rect 141114 77920 141142 77948
rect 141004 77868 141010 77920
rect 141062 77868 141068 77920
rect 141096 77868 141102 77920
rect 141154 77868 141160 77920
rect 141188 77868 141194 77920
rect 141246 77868 141252 77920
rect 141280 77868 141286 77920
rect 141338 77868 141344 77920
rect 141556 77908 141562 77920
rect 141528 77868 141562 77908
rect 141614 77868 141620 77920
rect 141648 77868 141654 77920
rect 141706 77868 141712 77920
rect 141832 77868 141838 77920
rect 141890 77868 141896 77920
rect 141924 77868 141930 77920
rect 141982 77868 141988 77920
rect 141022 77432 141050 77868
rect 141206 77648 141234 77868
rect 141142 77596 141148 77648
rect 141200 77608 141234 77648
rect 141200 77596 141206 77608
rect 141298 77512 141326 77868
rect 141298 77472 141332 77512
rect 141326 77460 141332 77472
rect 141384 77460 141390 77512
rect 141234 77432 141240 77444
rect 141022 77404 141240 77432
rect 141234 77392 141240 77404
rect 141292 77392 141298 77444
rect 141142 77364 141148 77376
rect 140930 77336 141148 77364
rect 141142 77324 141148 77336
rect 141200 77324 141206 77376
rect 138566 77228 138572 77240
rect 138032 77200 138572 77228
rect 118844 77188 118850 77200
rect 138566 77188 138572 77200
rect 138624 77188 138630 77240
rect 140958 77188 140964 77240
rect 141016 77228 141022 77240
rect 141528 77228 141556 77868
rect 141666 77784 141694 77868
rect 141850 77840 141878 77868
rect 141602 77732 141608 77784
rect 141660 77744 141694 77784
rect 141804 77812 141878 77840
rect 141660 77732 141666 77744
rect 141804 77648 141832 77812
rect 141942 77716 141970 77868
rect 141878 77664 141884 77716
rect 141936 77676 141970 77716
rect 141936 77664 141942 77676
rect 141786 77596 141792 77648
rect 141844 77596 141850 77648
rect 142080 77432 142108 78016
rect 142494 77920 142522 78016
rect 142200 77868 142206 77920
rect 142258 77868 142264 77920
rect 142292 77868 142298 77920
rect 142350 77868 142356 77920
rect 142476 77868 142482 77920
rect 142534 77868 142540 77920
rect 142568 77868 142574 77920
rect 142626 77868 142632 77920
rect 142660 77868 142666 77920
rect 142718 77868 142724 77920
rect 142752 77868 142758 77920
rect 142810 77908 142816 77920
rect 142810 77880 143166 77908
rect 142810 77868 142816 77880
rect 142218 77716 142246 77868
rect 142310 77840 142338 77868
rect 142310 77812 142476 77840
rect 142218 77676 142252 77716
rect 142246 77664 142252 77676
rect 142304 77664 142310 77716
rect 142448 77648 142476 77812
rect 142586 77772 142614 77868
rect 142540 77744 142614 77772
rect 142430 77596 142436 77648
rect 142488 77596 142494 77648
rect 142540 77636 142568 77744
rect 142678 77716 142706 77868
rect 143028 77800 143034 77852
rect 143086 77800 143092 77852
rect 142614 77664 142620 77716
rect 142672 77676 142706 77716
rect 142672 77664 142678 77676
rect 142706 77636 142712 77648
rect 142540 77608 142712 77636
rect 142706 77596 142712 77608
rect 142764 77596 142770 77648
rect 142338 77528 142344 77580
rect 142396 77568 142402 77580
rect 142890 77568 142896 77580
rect 142396 77540 142896 77568
rect 142396 77528 142402 77540
rect 142890 77528 142896 77540
rect 142948 77528 142954 77580
rect 142154 77460 142160 77512
rect 142212 77500 142218 77512
rect 143046 77500 143074 77800
rect 142212 77472 143074 77500
rect 142212 77460 142218 77472
rect 142338 77432 142344 77444
rect 142080 77404 142344 77432
rect 142338 77392 142344 77404
rect 142396 77392 142402 77444
rect 142614 77324 142620 77376
rect 142672 77364 142678 77376
rect 143138 77364 143166 77880
rect 143304 77868 143310 77920
rect 143362 77868 143368 77920
rect 143322 77444 143350 77868
rect 143488 77800 143494 77852
rect 143546 77800 143552 77852
rect 143506 77444 143534 77800
rect 143736 77772 143764 78152
rect 143856 77868 143862 77920
rect 143914 77868 143920 77920
rect 143948 77868 143954 77920
rect 144006 77868 144012 77920
rect 144040 77868 144046 77920
rect 144098 77868 144104 77920
rect 144408 77868 144414 77920
rect 144466 77868 144472 77920
rect 144500 77868 144506 77920
rect 144558 77868 144564 77920
rect 143644 77744 143764 77772
rect 143644 77580 143672 77744
rect 143626 77528 143632 77580
rect 143684 77528 143690 77580
rect 143874 77500 143902 77868
rect 143966 77568 143994 77868
rect 144058 77716 144086 77868
rect 144132 77800 144138 77852
rect 144190 77840 144196 77852
rect 144190 77800 144224 77840
rect 144058 77676 144092 77716
rect 144086 77664 144092 77676
rect 144144 77664 144150 77716
rect 144196 77580 144224 77800
rect 144426 77772 144454 77868
rect 144288 77744 144454 77772
rect 143966 77540 144132 77568
rect 143994 77500 144000 77512
rect 143874 77472 144000 77500
rect 143994 77460 144000 77472
rect 144052 77460 144058 77512
rect 143258 77392 143264 77444
rect 143316 77404 143350 77444
rect 143316 77392 143322 77404
rect 143442 77392 143448 77444
rect 143500 77404 143534 77444
rect 143500 77392 143506 77404
rect 143902 77392 143908 77444
rect 143960 77432 143966 77444
rect 144104 77432 144132 77540
rect 144178 77528 144184 77580
rect 144236 77528 144242 77580
rect 143960 77404 144132 77432
rect 143960 77392 143966 77404
rect 142672 77336 143166 77364
rect 142672 77324 142678 77336
rect 143534 77256 143540 77308
rect 143592 77296 143598 77308
rect 144288 77296 144316 77744
rect 144518 77716 144546 77868
rect 144454 77664 144460 77716
rect 144512 77676 144546 77716
rect 144512 77664 144518 77676
rect 144610 77648 144638 78424
rect 144546 77596 144552 77648
rect 144604 77608 144638 77648
rect 144604 77596 144610 77608
rect 143592 77268 144316 77296
rect 143592 77256 143598 77268
rect 141016 77200 141556 77228
rect 144702 77228 144730 78492
rect 144794 77432 144822 78628
rect 154546 78520 154574 78696
rect 166966 78656 166994 78696
rect 168346 78696 180340 78724
rect 168346 78656 168374 78696
rect 180334 78684 180340 78696
rect 180392 78684 180398 78736
rect 174538 78656 174544 78668
rect 146956 78492 154574 78520
rect 162826 78628 164234 78656
rect 166966 78628 168374 78656
rect 171106 78628 174544 78656
rect 146956 78248 146984 78492
rect 145024 78220 146984 78248
rect 154546 78424 155954 78452
rect 145024 77500 145052 78220
rect 154546 78180 154574 78424
rect 145898 78152 154574 78180
rect 155926 78180 155954 78424
rect 162826 78180 162854 78628
rect 164206 78588 164234 78628
rect 171106 78588 171134 78628
rect 174538 78616 174544 78628
rect 174596 78616 174602 78668
rect 164206 78560 171134 78588
rect 165586 78492 166994 78520
rect 165586 78452 165614 78492
rect 155926 78152 158484 78180
rect 145346 78016 145834 78044
rect 145144 77840 145150 77852
rect 144886 77472 145052 77500
rect 145116 77800 145150 77840
rect 145202 77800 145208 77852
rect 145236 77800 145242 77852
rect 145294 77800 145300 77852
rect 145346 77840 145374 78016
rect 145438 77948 145742 77976
rect 145438 77920 145466 77948
rect 145420 77868 145426 77920
rect 145478 77868 145484 77920
rect 145512 77868 145518 77920
rect 145570 77868 145576 77920
rect 145604 77868 145610 77920
rect 145662 77868 145668 77920
rect 145346 77812 145466 77840
rect 145116 77500 145144 77800
rect 145254 77580 145282 77800
rect 145328 77732 145334 77784
rect 145386 77732 145392 77784
rect 145190 77528 145196 77580
rect 145248 77540 145282 77580
rect 145346 77580 145374 77732
rect 145438 77716 145466 77812
rect 145420 77664 145426 77716
rect 145478 77664 145484 77716
rect 145346 77540 145380 77580
rect 145248 77528 145254 77540
rect 145374 77528 145380 77540
rect 145432 77528 145438 77580
rect 145530 77500 145558 77868
rect 145622 77784 145650 77868
rect 145604 77732 145610 77784
rect 145662 77732 145668 77784
rect 145714 77568 145742 77948
rect 145806 77920 145834 78016
rect 145788 77868 145794 77920
rect 145846 77868 145852 77920
rect 145898 77580 145926 78152
rect 153166 78084 156046 78112
rect 153166 78044 153194 78084
rect 152338 78016 153194 78044
rect 154500 78016 155172 78044
rect 146174 77948 146754 77976
rect 146064 77868 146070 77920
rect 146122 77868 146128 77920
rect 145714 77540 145788 77568
rect 145650 77500 145656 77512
rect 145116 77472 145282 77500
rect 145530 77472 145656 77500
rect 144886 77432 144914 77472
rect 144794 77404 144914 77432
rect 145254 77444 145282 77472
rect 145650 77460 145656 77472
rect 145708 77460 145714 77512
rect 145254 77404 145288 77444
rect 145282 77392 145288 77404
rect 145340 77392 145346 77444
rect 145466 77392 145472 77444
rect 145524 77392 145530 77444
rect 145484 77364 145512 77392
rect 145116 77336 145512 77364
rect 144914 77256 144920 77308
rect 144972 77296 144978 77308
rect 145116 77296 145144 77336
rect 144972 77268 145144 77296
rect 144972 77256 144978 77268
rect 145466 77256 145472 77308
rect 145524 77296 145530 77308
rect 145760 77296 145788 77540
rect 145834 77528 145840 77580
rect 145892 77540 145926 77580
rect 145892 77528 145898 77540
rect 145834 77392 145840 77444
rect 145892 77432 145898 77444
rect 146082 77432 146110 77868
rect 145892 77404 146110 77432
rect 146174 77432 146202 77948
rect 146726 77920 146754 77948
rect 147738 77948 150940 77976
rect 147738 77920 147766 77948
rect 146266 77880 146478 77908
rect 146266 77500 146294 77880
rect 146450 77852 146478 77880
rect 146708 77868 146714 77920
rect 146766 77868 146772 77920
rect 147168 77908 147174 77920
rect 147140 77868 147174 77908
rect 147226 77868 147232 77920
rect 147260 77868 147266 77920
rect 147318 77868 147324 77920
rect 147352 77868 147358 77920
rect 147410 77868 147416 77920
rect 147444 77868 147450 77920
rect 147502 77868 147508 77920
rect 147536 77868 147542 77920
rect 147594 77868 147600 77920
rect 147628 77868 147634 77920
rect 147686 77868 147692 77920
rect 147720 77868 147726 77920
rect 147778 77868 147784 77920
rect 147996 77868 148002 77920
rect 148054 77868 148060 77920
rect 148272 77868 148278 77920
rect 148330 77868 148336 77920
rect 148364 77868 148370 77920
rect 148422 77868 148428 77920
rect 148456 77868 148462 77920
rect 148514 77868 148520 77920
rect 148548 77868 148554 77920
rect 148606 77868 148612 77920
rect 148732 77908 148738 77920
rect 148704 77868 148738 77908
rect 148790 77868 148796 77920
rect 148824 77868 148830 77920
rect 148882 77868 148888 77920
rect 148916 77868 148922 77920
rect 148974 77868 148980 77920
rect 149008 77868 149014 77920
rect 149066 77868 149072 77920
rect 149192 77908 149198 77920
rect 149164 77868 149198 77908
rect 149250 77868 149256 77920
rect 149284 77868 149290 77920
rect 149342 77868 149348 77920
rect 149376 77868 149382 77920
rect 149434 77868 149440 77920
rect 149468 77868 149474 77920
rect 149526 77868 149532 77920
rect 149744 77908 149750 77920
rect 149578 77880 149750 77908
rect 146340 77800 146346 77852
rect 146398 77800 146404 77852
rect 146432 77800 146438 77852
rect 146490 77800 146496 77852
rect 146358 77568 146386 77800
rect 146984 77732 146990 77784
rect 147042 77732 147048 77784
rect 146846 77596 146852 77648
rect 146904 77636 146910 77648
rect 147002 77636 147030 77732
rect 146904 77608 147030 77636
rect 146904 77596 146910 77608
rect 146938 77568 146944 77580
rect 146358 77540 146944 77568
rect 146938 77528 146944 77540
rect 146996 77528 147002 77580
rect 146386 77500 146392 77512
rect 146266 77472 146392 77500
rect 146386 77460 146392 77472
rect 146444 77460 146450 77512
rect 146662 77460 146668 77512
rect 146720 77500 146726 77512
rect 147140 77500 147168 77868
rect 147278 77840 147306 77868
rect 147232 77812 147306 77840
rect 147232 77784 147260 77812
rect 147214 77732 147220 77784
rect 147272 77732 147278 77784
rect 147370 77772 147398 77868
rect 147324 77744 147398 77772
rect 147324 77716 147352 77744
rect 147462 77716 147490 77868
rect 147306 77664 147312 77716
rect 147364 77664 147370 77716
rect 147398 77664 147404 77716
rect 147456 77676 147490 77716
rect 147456 77664 147462 77676
rect 147554 77648 147582 77868
rect 147646 77784 147674 77868
rect 147646 77744 147680 77784
rect 147674 77732 147680 77744
rect 147732 77732 147738 77784
rect 147490 77596 147496 77648
rect 147548 77608 147582 77648
rect 147548 77596 147554 77608
rect 148014 77580 148042 77868
rect 148290 77840 148318 77868
rect 148244 77812 148318 77840
rect 148244 77636 148272 77812
rect 148382 77784 148410 77868
rect 148318 77732 148324 77784
rect 148376 77744 148410 77784
rect 148376 77732 148382 77744
rect 148318 77636 148324 77648
rect 148244 77608 148324 77636
rect 148318 77596 148324 77608
rect 148376 77596 148382 77648
rect 147950 77528 147956 77580
rect 148008 77540 148042 77580
rect 148008 77528 148014 77540
rect 146720 77472 147168 77500
rect 146720 77460 146726 77472
rect 146294 77432 146300 77444
rect 146174 77404 146300 77432
rect 145892 77392 145898 77404
rect 146294 77392 146300 77404
rect 146352 77392 146358 77444
rect 148226 77392 148232 77444
rect 148284 77432 148290 77444
rect 148474 77432 148502 77868
rect 148284 77404 148502 77432
rect 148284 77392 148290 77404
rect 148566 77376 148594 77868
rect 148704 77580 148732 77868
rect 148842 77840 148870 77868
rect 148796 77812 148870 77840
rect 148796 77716 148824 77812
rect 148934 77772 148962 77868
rect 148888 77744 148962 77772
rect 148888 77716 148916 77744
rect 149026 77716 149054 77868
rect 148778 77664 148784 77716
rect 148836 77664 148842 77716
rect 148870 77664 148876 77716
rect 148928 77664 148934 77716
rect 148962 77664 148968 77716
rect 149020 77676 149054 77716
rect 149020 77664 149026 77676
rect 148686 77528 148692 77580
rect 148744 77528 148750 77580
rect 148502 77324 148508 77376
rect 148560 77336 148594 77376
rect 149164 77364 149192 77868
rect 149302 77840 149330 77868
rect 149256 77812 149330 77840
rect 149256 77784 149284 77812
rect 149238 77732 149244 77784
rect 149296 77732 149302 77784
rect 149394 77772 149422 77868
rect 149348 77744 149422 77772
rect 149348 77716 149376 77744
rect 149486 77716 149514 77868
rect 149330 77664 149336 77716
rect 149388 77664 149394 77716
rect 149422 77664 149428 77716
rect 149480 77676 149514 77716
rect 149480 77664 149486 77676
rect 149578 77512 149606 77880
rect 149744 77868 149750 77880
rect 149802 77868 149808 77920
rect 149836 77868 149842 77920
rect 149894 77868 149900 77920
rect 149928 77868 149934 77920
rect 149986 77868 149992 77920
rect 150112 77868 150118 77920
rect 150170 77868 150176 77920
rect 150296 77908 150302 77920
rect 150268 77868 150302 77908
rect 150354 77868 150360 77920
rect 150388 77868 150394 77920
rect 150446 77868 150452 77920
rect 150480 77868 150486 77920
rect 150538 77868 150544 77920
rect 150572 77868 150578 77920
rect 150630 77868 150636 77920
rect 149854 77840 149882 77868
rect 149808 77812 149882 77840
rect 149808 77784 149836 77812
rect 149946 77784 149974 77868
rect 149652 77732 149658 77784
rect 149710 77772 149716 77784
rect 149710 77732 149744 77772
rect 149790 77732 149796 77784
rect 149848 77732 149854 77784
rect 149882 77732 149888 77784
rect 149940 77744 149974 77784
rect 149940 77732 149946 77744
rect 149716 77648 149744 77732
rect 150130 77648 150158 77868
rect 149698 77596 149704 77648
rect 149756 77596 149762 77648
rect 150130 77608 150164 77648
rect 150158 77596 150164 77608
rect 150216 77596 150222 77648
rect 149974 77528 149980 77580
rect 150032 77568 150038 77580
rect 150268 77568 150296 77868
rect 150406 77840 150434 77868
rect 150360 77812 150434 77840
rect 150360 77784 150388 77812
rect 150342 77732 150348 77784
rect 150400 77732 150406 77784
rect 150498 77772 150526 77868
rect 150452 77744 150526 77772
rect 150032 77540 150296 77568
rect 150032 77528 150038 77540
rect 149578 77472 149612 77512
rect 149606 77460 149612 77472
rect 149664 77460 149670 77512
rect 149330 77364 149336 77376
rect 149164 77336 149336 77364
rect 148560 77324 148566 77336
rect 149330 77324 149336 77336
rect 149388 77324 149394 77376
rect 150452 77364 150480 77744
rect 150590 77716 150618 77868
rect 150526 77664 150532 77716
rect 150584 77676 150618 77716
rect 150584 77664 150590 77676
rect 150912 77432 150940 77948
rect 151032 77868 151038 77920
rect 151090 77868 151096 77920
rect 151124 77868 151130 77920
rect 151182 77868 151188 77920
rect 151308 77868 151314 77920
rect 151366 77868 151372 77920
rect 151492 77868 151498 77920
rect 151550 77868 151556 77920
rect 151768 77868 151774 77920
rect 151826 77868 151832 77920
rect 151860 77868 151866 77920
rect 151918 77908 151924 77920
rect 152136 77908 152142 77920
rect 151918 77868 151952 77908
rect 151050 77716 151078 77868
rect 150986 77664 150992 77716
rect 151044 77676 151078 77716
rect 151044 77664 151050 77676
rect 151142 77648 151170 77868
rect 151142 77608 151176 77648
rect 151170 77596 151176 77608
rect 151228 77596 151234 77648
rect 151326 77580 151354 77868
rect 151510 77704 151538 77868
rect 151786 77784 151814 77868
rect 151722 77732 151728 77784
rect 151780 77744 151814 77784
rect 151780 77732 151786 77744
rect 151814 77704 151820 77716
rect 151510 77676 151820 77704
rect 151814 77664 151820 77676
rect 151872 77664 151878 77716
rect 151326 77540 151360 77580
rect 151354 77528 151360 77540
rect 151412 77528 151418 77580
rect 151924 77568 151952 77868
rect 152016 77880 152142 77908
rect 152016 77636 152044 77880
rect 152136 77868 152142 77880
rect 152194 77868 152200 77920
rect 152338 77772 152366 78016
rect 153258 77948 154022 77976
rect 153258 77920 153286 77948
rect 152412 77868 152418 77920
rect 152470 77868 152476 77920
rect 152504 77868 152510 77920
rect 152562 77908 152568 77920
rect 152562 77868 152596 77908
rect 152688 77868 152694 77920
rect 152746 77868 152752 77920
rect 152872 77868 152878 77920
rect 152930 77868 152936 77920
rect 152964 77868 152970 77920
rect 153022 77868 153028 77920
rect 153056 77868 153062 77920
rect 153114 77868 153120 77920
rect 153240 77868 153246 77920
rect 153298 77868 153304 77920
rect 153884 77908 153890 77920
rect 153396 77880 153890 77908
rect 152430 77840 152458 77868
rect 152430 77812 152504 77840
rect 152338 77744 152412 77772
rect 152182 77636 152188 77648
rect 152016 77608 152188 77636
rect 152182 77596 152188 77608
rect 152240 77596 152246 77648
rect 152274 77568 152280 77580
rect 151924 77540 152280 77568
rect 152274 77528 152280 77540
rect 152332 77528 152338 77580
rect 151998 77460 152004 77512
rect 152056 77500 152062 77512
rect 152384 77500 152412 77744
rect 152476 77716 152504 77812
rect 152458 77664 152464 77716
rect 152516 77664 152522 77716
rect 152568 77648 152596 77868
rect 152550 77596 152556 77648
rect 152608 77596 152614 77648
rect 152706 77580 152734 77868
rect 152890 77840 152918 77868
rect 152844 77812 152918 77840
rect 152844 77716 152872 77812
rect 152982 77716 153010 77868
rect 152826 77664 152832 77716
rect 152884 77664 152890 77716
rect 152918 77664 152924 77716
rect 152976 77676 153010 77716
rect 153074 77704 153102 77868
rect 153074 77676 153240 77704
rect 152976 77664 152982 77676
rect 153212 77580 153240 77676
rect 152642 77528 152648 77580
rect 152700 77540 152734 77580
rect 152700 77528 152706 77540
rect 153194 77528 153200 77580
rect 153252 77528 153258 77580
rect 153396 77512 153424 77880
rect 153884 77868 153890 77880
rect 153942 77868 153948 77920
rect 153792 77840 153798 77852
rect 153764 77800 153798 77840
rect 153850 77800 153856 77852
rect 153764 77716 153792 77800
rect 153746 77664 153752 77716
rect 153804 77664 153810 77716
rect 153994 77648 154022 77948
rect 154160 77800 154166 77852
rect 154218 77800 154224 77852
rect 154252 77800 154258 77852
rect 154310 77800 154316 77852
rect 154178 77716 154206 77800
rect 154114 77664 154120 77716
rect 154172 77676 154206 77716
rect 154172 77664 154178 77676
rect 153930 77596 153936 77648
rect 153988 77608 154022 77648
rect 153988 77596 153994 77608
rect 152056 77472 152412 77500
rect 152056 77460 152062 77472
rect 153378 77460 153384 77512
rect 153436 77460 153442 77512
rect 154270 77500 154298 77800
rect 154390 77500 154396 77512
rect 154270 77472 154396 77500
rect 154390 77460 154396 77472
rect 154448 77460 154454 77512
rect 154500 77432 154528 78016
rect 154804 77868 154810 77920
rect 154862 77868 154868 77920
rect 154822 77772 154850 77868
rect 154776 77744 154850 77772
rect 154776 77636 154804 77744
rect 154942 77636 154948 77648
rect 154776 77608 154948 77636
rect 154942 77596 154948 77608
rect 155000 77596 155006 77648
rect 150912 77404 154528 77432
rect 150452 77336 152964 77364
rect 145524 77268 145788 77296
rect 145524 77256 145530 77268
rect 149054 77256 149060 77308
rect 149112 77296 149118 77308
rect 152366 77296 152372 77308
rect 149112 77268 152372 77296
rect 149112 77256 149118 77268
rect 152366 77256 152372 77268
rect 152424 77256 152430 77308
rect 152936 77296 152964 77336
rect 154666 77324 154672 77376
rect 154724 77364 154730 77376
rect 154850 77364 154856 77376
rect 154724 77336 154856 77364
rect 154724 77324 154730 77336
rect 154850 77324 154856 77336
rect 154908 77324 154914 77376
rect 155144 77364 155172 78016
rect 155264 77908 155270 77920
rect 155236 77868 155270 77908
rect 155322 77868 155328 77920
rect 155356 77868 155362 77920
rect 155414 77868 155420 77920
rect 155448 77868 155454 77920
rect 155506 77868 155512 77920
rect 155724 77868 155730 77920
rect 155782 77868 155788 77920
rect 155816 77868 155822 77920
rect 155874 77868 155880 77920
rect 155236 77580 155264 77868
rect 155374 77840 155402 77868
rect 155328 77812 155402 77840
rect 155218 77528 155224 77580
rect 155276 77528 155282 77580
rect 155328 77432 155356 77812
rect 155466 77716 155494 77868
rect 155742 77840 155770 77868
rect 155402 77664 155408 77716
rect 155460 77676 155494 77716
rect 155604 77812 155770 77840
rect 155460 77664 155466 77676
rect 155604 77648 155632 77812
rect 155834 77784 155862 77868
rect 155834 77744 155868 77784
rect 155862 77732 155868 77744
rect 155920 77732 155926 77784
rect 155586 77596 155592 77648
rect 155644 77596 155650 77648
rect 156018 77500 156046 78084
rect 156478 77948 156690 77976
rect 156478 77920 156506 77948
rect 156092 77868 156098 77920
rect 156150 77868 156156 77920
rect 156368 77868 156374 77920
rect 156426 77868 156432 77920
rect 156460 77868 156466 77920
rect 156518 77868 156524 77920
rect 156552 77868 156558 77920
rect 156610 77868 156616 77920
rect 156110 77636 156138 77868
rect 156386 77784 156414 77868
rect 156386 77744 156420 77784
rect 156414 77732 156420 77744
rect 156472 77732 156478 77784
rect 156570 77648 156598 77868
rect 156230 77636 156236 77648
rect 156110 77608 156236 77636
rect 156230 77596 156236 77608
rect 156288 77596 156294 77648
rect 156506 77596 156512 77648
rect 156564 77608 156598 77648
rect 156564 77596 156570 77608
rect 156662 77580 156690 77948
rect 156736 77868 156742 77920
rect 156794 77868 156800 77920
rect 156828 77868 156834 77920
rect 156886 77868 156892 77920
rect 157288 77868 157294 77920
rect 157346 77908 157352 77920
rect 157472 77908 157478 77920
rect 157346 77868 157380 77908
rect 156754 77784 156782 77868
rect 156846 77840 156874 77868
rect 156846 77812 156920 77840
rect 156754 77744 156788 77784
rect 156782 77732 156788 77744
rect 156840 77732 156846 77784
rect 156892 77580 156920 77812
rect 157352 77716 157380 77868
rect 157444 77868 157478 77908
rect 157530 77868 157536 77920
rect 157564 77868 157570 77920
rect 157622 77868 157628 77920
rect 157656 77868 157662 77920
rect 157714 77868 157720 77920
rect 157840 77868 157846 77920
rect 157898 77868 157904 77920
rect 157932 77868 157938 77920
rect 157990 77868 157996 77920
rect 158208 77908 158214 77920
rect 158180 77868 158214 77908
rect 158266 77868 158272 77920
rect 158300 77868 158306 77920
rect 158358 77868 158364 77920
rect 157334 77664 157340 77716
rect 157392 77664 157398 77716
rect 157150 77596 157156 77648
rect 157208 77636 157214 77648
rect 157444 77636 157472 77868
rect 157582 77784 157610 77868
rect 157518 77732 157524 77784
rect 157576 77744 157610 77784
rect 157674 77784 157702 77868
rect 157674 77744 157708 77784
rect 157576 77732 157582 77744
rect 157702 77732 157708 77744
rect 157760 77732 157766 77784
rect 157858 77704 157886 77868
rect 157720 77676 157886 77704
rect 157720 77648 157748 77676
rect 157208 77608 157472 77636
rect 157208 77596 157214 77608
rect 157702 77596 157708 77648
rect 157760 77596 157766 77648
rect 157794 77596 157800 77648
rect 157852 77636 157858 77648
rect 157950 77636 157978 77868
rect 157852 77608 157978 77636
rect 158180 77636 158208 77868
rect 158318 77716 158346 77868
rect 158254 77664 158260 77716
rect 158312 77676 158346 77716
rect 158312 77664 158318 77676
rect 158180 77608 158300 77636
rect 157852 77596 157858 77608
rect 156598 77528 156604 77580
rect 156656 77540 156690 77580
rect 156656 77528 156662 77540
rect 156874 77528 156880 77580
rect 156932 77528 156938 77580
rect 156966 77528 156972 77580
rect 157024 77568 157030 77580
rect 157242 77568 157248 77580
rect 157024 77540 157248 77568
rect 157024 77528 157030 77540
rect 157242 77528 157248 77540
rect 157300 77528 157306 77580
rect 156018 77472 157104 77500
rect 156966 77432 156972 77444
rect 155328 77404 156972 77432
rect 156966 77392 156972 77404
rect 157024 77392 157030 77444
rect 157076 77432 157104 77472
rect 158070 77460 158076 77512
rect 158128 77500 158134 77512
rect 158272 77500 158300 77608
rect 158456 77512 158484 78152
rect 158548 78152 162854 78180
rect 164206 78424 165614 78452
rect 166966 78452 166994 78492
rect 168346 78492 171134 78520
rect 168346 78452 168374 78492
rect 166966 78424 168374 78452
rect 171106 78452 171134 78492
rect 175918 78452 175924 78464
rect 171106 78424 175924 78452
rect 158128 77472 158300 77500
rect 158128 77460 158134 77472
rect 158438 77460 158444 77512
rect 158496 77460 158502 77512
rect 158548 77432 158576 78152
rect 160526 78084 163222 78112
rect 158640 78016 160278 78044
rect 158640 77500 158668 78016
rect 158732 77948 160094 77976
rect 158732 77568 158760 77948
rect 160066 77920 160094 77948
rect 158852 77908 158858 77920
rect 158824 77868 158858 77908
rect 158910 77868 158916 77920
rect 158944 77868 158950 77920
rect 159002 77868 159008 77920
rect 159036 77868 159042 77920
rect 159094 77868 159100 77920
rect 159128 77868 159134 77920
rect 159186 77868 159192 77920
rect 159588 77868 159594 77920
rect 159646 77868 159652 77920
rect 159772 77868 159778 77920
rect 159830 77868 159836 77920
rect 159864 77868 159870 77920
rect 159922 77868 159928 77920
rect 159956 77868 159962 77920
rect 160014 77868 160020 77920
rect 160048 77868 160054 77920
rect 160106 77868 160112 77920
rect 160140 77868 160146 77920
rect 160198 77868 160204 77920
rect 158824 77648 158852 77868
rect 158962 77648 158990 77868
rect 159054 77704 159082 77868
rect 159146 77772 159174 77868
rect 159312 77800 159318 77852
rect 159370 77800 159376 77852
rect 159404 77800 159410 77852
rect 159462 77800 159468 77852
rect 159146 77744 159220 77772
rect 159054 77676 159128 77704
rect 159100 77648 159128 77676
rect 158806 77596 158812 77648
rect 158864 77596 158870 77648
rect 158962 77608 158996 77648
rect 158990 77596 158996 77608
rect 159048 77596 159054 77648
rect 159082 77596 159088 77648
rect 159140 77596 159146 77648
rect 159192 77580 159220 77744
rect 158898 77568 158904 77580
rect 158732 77540 158904 77568
rect 158898 77528 158904 77540
rect 158956 77528 158962 77580
rect 159174 77528 159180 77580
rect 159232 77528 159238 77580
rect 159330 77512 159358 77800
rect 158640 77472 158852 77500
rect 157076 77404 158576 77432
rect 158824 77364 158852 77472
rect 159266 77460 159272 77512
rect 159324 77472 159358 77512
rect 159324 77460 159330 77472
rect 159422 77376 159450 77800
rect 159606 77704 159634 77868
rect 159560 77676 159634 77704
rect 159560 77568 159588 77676
rect 159634 77596 159640 77648
rect 159692 77636 159698 77648
rect 159790 77636 159818 77868
rect 159692 77608 159818 77636
rect 159882 77648 159910 77868
rect 159974 77840 160002 77868
rect 159974 77812 160048 77840
rect 160020 77648 160048 77812
rect 160158 77704 160186 77868
rect 160112 77676 160186 77704
rect 160112 77648 160140 77676
rect 159882 77608 159916 77648
rect 159692 77596 159698 77608
rect 159910 77596 159916 77608
rect 159968 77596 159974 77648
rect 160002 77596 160008 77648
rect 160060 77596 160066 77648
rect 160094 77596 160100 77648
rect 160152 77596 160158 77648
rect 160250 77636 160278 78016
rect 160526 77976 160554 78084
rect 160434 77948 160554 77976
rect 160756 78016 161290 78044
rect 160324 77868 160330 77920
rect 160382 77868 160388 77920
rect 160204 77608 160278 77636
rect 159560 77540 160048 77568
rect 155144 77336 158852 77364
rect 159358 77324 159364 77376
rect 159416 77336 159450 77376
rect 159416 77324 159422 77336
rect 156690 77296 156696 77308
rect 152936 77268 156696 77296
rect 156690 77256 156696 77268
rect 156748 77256 156754 77308
rect 158438 77256 158444 77308
rect 158496 77296 158502 77308
rect 160020 77296 160048 77540
rect 160204 77432 160232 77608
rect 160342 77580 160370 77868
rect 160278 77528 160284 77580
rect 160336 77540 160370 77580
rect 160336 77528 160342 77540
rect 160434 77500 160462 77948
rect 160508 77868 160514 77920
rect 160566 77868 160572 77920
rect 160526 77648 160554 77868
rect 160600 77800 160606 77852
rect 160658 77840 160664 77852
rect 160658 77800 160692 77840
rect 160526 77608 160560 77648
rect 160554 77596 160560 77608
rect 160612 77596 160618 77648
rect 160664 77580 160692 77800
rect 160756 77648 160784 78016
rect 160986 77948 161198 77976
rect 160986 77920 161014 77948
rect 160876 77868 160882 77920
rect 160934 77868 160940 77920
rect 160968 77868 160974 77920
rect 161026 77868 161032 77920
rect 160894 77716 160922 77868
rect 160894 77676 160928 77716
rect 160922 77664 160928 77676
rect 160980 77664 160986 77716
rect 160738 77596 160744 77648
rect 160796 77596 160802 77648
rect 160646 77528 160652 77580
rect 160704 77528 160710 77580
rect 161014 77528 161020 77580
rect 161072 77568 161078 77580
rect 161170 77568 161198 77948
rect 161262 77852 161290 78016
rect 161630 77948 161934 77976
rect 161630 77920 161658 77948
rect 161612 77868 161618 77920
rect 161670 77868 161676 77920
rect 161704 77868 161710 77920
rect 161762 77868 161768 77920
rect 161796 77868 161802 77920
rect 161854 77868 161860 77920
rect 161244 77800 161250 77852
rect 161302 77800 161308 77852
rect 161336 77800 161342 77852
rect 161394 77800 161400 77852
rect 161428 77800 161434 77852
rect 161486 77800 161492 77852
rect 161354 77772 161382 77800
rect 161308 77744 161382 77772
rect 161308 77716 161336 77744
rect 161446 77716 161474 77800
rect 161290 77664 161296 77716
rect 161348 77664 161354 77716
rect 161382 77664 161388 77716
rect 161440 77676 161474 77716
rect 161440 77664 161446 77676
rect 161072 77540 161198 77568
rect 161722 77580 161750 77868
rect 161814 77636 161842 77868
rect 161906 77772 161934 77948
rect 161998 77948 162348 77976
rect 161998 77920 162026 77948
rect 161980 77868 161986 77920
rect 162038 77868 162044 77920
rect 162164 77868 162170 77920
rect 162222 77868 162228 77920
rect 162072 77840 162078 77852
rect 162044 77800 162078 77840
rect 162130 77800 162136 77852
rect 161906 77744 161980 77772
rect 161814 77608 161888 77636
rect 161722 77540 161756 77580
rect 161072 77528 161078 77540
rect 161750 77528 161756 77540
rect 161808 77528 161814 77580
rect 161198 77500 161204 77512
rect 160434 77472 161204 77500
rect 161198 77460 161204 77472
rect 161256 77460 161262 77512
rect 161658 77460 161664 77512
rect 161716 77500 161722 77512
rect 161860 77500 161888 77608
rect 161952 77580 161980 77744
rect 162044 77716 162072 77800
rect 162182 77716 162210 77868
rect 162026 77664 162032 77716
rect 162084 77664 162090 77716
rect 162118 77664 162124 77716
rect 162176 77676 162210 77716
rect 162176 77664 162182 77676
rect 162320 77648 162348 77948
rect 162734 77948 162854 77976
rect 162440 77868 162446 77920
rect 162498 77868 162504 77920
rect 162624 77868 162630 77920
rect 162682 77868 162688 77920
rect 162458 77840 162486 77868
rect 162412 77812 162486 77840
rect 162302 77596 162308 77648
rect 162360 77596 162366 77648
rect 161934 77528 161940 77580
rect 161992 77528 161998 77580
rect 161716 77472 161888 77500
rect 161716 77460 161722 77472
rect 162210 77432 162216 77444
rect 160204 77404 162216 77432
rect 162210 77392 162216 77404
rect 162268 77392 162274 77444
rect 162412 77432 162440 77812
rect 162642 77772 162670 77868
rect 162504 77744 162670 77772
rect 162504 77512 162532 77744
rect 162734 77704 162762 77948
rect 162826 77920 162854 77948
rect 162918 77948 163130 77976
rect 162918 77920 162946 77948
rect 162808 77868 162814 77920
rect 162866 77868 162872 77920
rect 162900 77868 162906 77920
rect 162958 77868 162964 77920
rect 162992 77868 162998 77920
rect 163050 77868 163056 77920
rect 162688 77676 162762 77704
rect 162486 77460 162492 77512
rect 162544 77460 162550 77512
rect 162578 77432 162584 77444
rect 162412 77404 162584 77432
rect 162578 77392 162584 77404
rect 162636 77392 162642 77444
rect 162688 77364 162716 77676
rect 162854 77596 162860 77648
rect 162912 77636 162918 77648
rect 163010 77636 163038 77868
rect 162912 77608 163038 77636
rect 162912 77596 162918 77608
rect 162762 77528 162768 77580
rect 162820 77568 162826 77580
rect 163102 77568 163130 77948
rect 162820 77540 163130 77568
rect 163194 77568 163222 78084
rect 163360 77868 163366 77920
rect 163418 77908 163424 77920
rect 163544 77908 163550 77920
rect 163418 77868 163452 77908
rect 163424 77784 163452 77868
rect 163516 77868 163550 77908
rect 163602 77868 163608 77920
rect 163636 77868 163642 77920
rect 163694 77868 163700 77920
rect 163728 77868 163734 77920
rect 163786 77868 163792 77920
rect 163820 77868 163826 77920
rect 163878 77868 163884 77920
rect 163912 77868 163918 77920
rect 163970 77868 163976 77920
rect 163406 77732 163412 77784
rect 163464 77732 163470 77784
rect 163516 77648 163544 77868
rect 163654 77840 163682 77868
rect 163608 77812 163682 77840
rect 163498 77596 163504 77648
rect 163556 77596 163562 77648
rect 163608 77636 163636 77812
rect 163746 77772 163774 77868
rect 163700 77744 163774 77772
rect 163700 77716 163728 77744
rect 163838 77716 163866 77868
rect 163930 77784 163958 77868
rect 163930 77744 163964 77784
rect 163958 77732 163964 77744
rect 164016 77732 164022 77784
rect 163682 77664 163688 77716
rect 163740 77664 163746 77716
rect 163774 77664 163780 77716
rect 163832 77676 163866 77716
rect 164206 77704 164234 78424
rect 175918 78412 175924 78424
rect 175976 78412 175982 78464
rect 174630 78316 174636 78328
rect 170278 78288 174636 78316
rect 165034 77948 165706 77976
rect 165034 77920 165062 77948
rect 164280 77868 164286 77920
rect 164338 77868 164344 77920
rect 164464 77868 164470 77920
rect 164522 77868 164528 77920
rect 164556 77868 164562 77920
rect 164614 77868 164620 77920
rect 164924 77868 164930 77920
rect 164982 77868 164988 77920
rect 165016 77868 165022 77920
rect 165074 77868 165080 77920
rect 165108 77868 165114 77920
rect 165166 77868 165172 77920
rect 165200 77868 165206 77920
rect 165258 77868 165264 77920
rect 163976 77676 164234 77704
rect 163832 77664 163838 77676
rect 163866 77636 163872 77648
rect 163608 77608 163872 77636
rect 163866 77596 163872 77608
rect 163924 77596 163930 77648
rect 163590 77568 163596 77580
rect 163194 77540 163596 77568
rect 162820 77528 162826 77540
rect 163590 77528 163596 77540
rect 163648 77528 163654 77580
rect 162946 77460 162952 77512
rect 163004 77500 163010 77512
rect 163976 77500 164004 77676
rect 164298 77648 164326 77868
rect 164482 77772 164510 77868
rect 164436 77744 164510 77772
rect 164298 77608 164332 77648
rect 164326 77596 164332 77608
rect 164384 77596 164390 77648
rect 164142 77528 164148 77580
rect 164200 77568 164206 77580
rect 164436 77568 164464 77744
rect 164574 77716 164602 77868
rect 164510 77664 164516 77716
rect 164568 77676 164602 77716
rect 164568 77664 164574 77676
rect 164942 77636 164970 77868
rect 165126 77772 165154 77868
rect 165080 77744 165154 77772
rect 165080 77716 165108 77744
rect 165218 77716 165246 77868
rect 165568 77800 165574 77852
rect 165626 77800 165632 77852
rect 165062 77664 165068 77716
rect 165120 77664 165126 77716
rect 165154 77664 165160 77716
rect 165212 77676 165246 77716
rect 165212 77664 165218 77676
rect 164200 77540 164464 77568
rect 164528 77608 164970 77636
rect 164200 77528 164206 77540
rect 163004 77472 164004 77500
rect 163004 77460 163010 77472
rect 164418 77460 164424 77512
rect 164476 77500 164482 77512
rect 164528 77500 164556 77608
rect 165246 77596 165252 77648
rect 165304 77636 165310 77648
rect 165586 77636 165614 77800
rect 165304 77608 165614 77636
rect 165304 77596 165310 77608
rect 164878 77528 164884 77580
rect 164936 77528 164942 77580
rect 164970 77528 164976 77580
rect 165028 77568 165034 77580
rect 165678 77568 165706 77948
rect 165862 77948 166166 77976
rect 165862 77784 165890 77948
rect 166138 77920 166166 77948
rect 165936 77868 165942 77920
rect 165994 77908 166000 77920
rect 165994 77880 166074 77908
rect 165994 77868 166000 77880
rect 165862 77744 165896 77784
rect 165890 77732 165896 77744
rect 165948 77732 165954 77784
rect 166046 77648 166074 77880
rect 166120 77868 166126 77920
rect 166178 77868 166184 77920
rect 166212 77868 166218 77920
rect 166270 77868 166276 77920
rect 166488 77868 166494 77920
rect 166546 77868 166552 77920
rect 166580 77868 166586 77920
rect 166638 77868 166644 77920
rect 166672 77868 166678 77920
rect 166730 77868 166736 77920
rect 167684 77908 167690 77920
rect 167564 77880 167690 77908
rect 166046 77608 166080 77648
rect 166074 77596 166080 77608
rect 166132 77596 166138 77648
rect 165028 77540 165706 77568
rect 165028 77528 165034 77540
rect 164476 77472 164556 77500
rect 164476 77460 164482 77472
rect 164694 77460 164700 77512
rect 164752 77500 164758 77512
rect 164896 77500 164924 77528
rect 164752 77472 164924 77500
rect 166230 77500 166258 77868
rect 166506 77840 166534 77868
rect 166460 77812 166534 77840
rect 166460 77636 166488 77812
rect 166598 77772 166626 77868
rect 166552 77744 166626 77772
rect 166552 77716 166580 77744
rect 166690 77716 166718 77868
rect 166534 77664 166540 77716
rect 166592 77664 166598 77716
rect 166626 77664 166632 77716
rect 166684 77676 166718 77716
rect 166684 77664 166690 77676
rect 166810 77636 166816 77648
rect 166460 77608 166816 77636
rect 166810 77596 166816 77608
rect 166868 77596 166874 77648
rect 166350 77500 166356 77512
rect 166230 77472 166356 77500
rect 164752 77460 164758 77472
rect 166350 77460 166356 77472
rect 166408 77460 166414 77512
rect 166902 77460 166908 77512
rect 166960 77500 166966 77512
rect 167564 77500 167592 77880
rect 167684 77868 167690 77880
rect 167742 77868 167748 77920
rect 167776 77868 167782 77920
rect 167834 77868 167840 77920
rect 168144 77908 168150 77920
rect 167932 77880 168150 77908
rect 167794 77716 167822 77868
rect 167932 77772 167960 77880
rect 168144 77868 168150 77880
rect 168202 77868 168208 77920
rect 168328 77868 168334 77920
rect 168386 77868 168392 77920
rect 168420 77868 168426 77920
rect 168478 77868 168484 77920
rect 168972 77868 168978 77920
rect 169030 77908 169036 77920
rect 169030 77880 169524 77908
rect 169030 77868 169036 77880
rect 168098 77772 168104 77784
rect 167932 77744 168104 77772
rect 168098 77732 168104 77744
rect 168156 77732 168162 77784
rect 167730 77664 167736 77716
rect 167788 77676 167822 77716
rect 167788 77664 167794 77676
rect 168346 77648 168374 77868
rect 168282 77596 168288 77648
rect 168340 77608 168374 77648
rect 168340 77596 168346 77608
rect 166960 77472 167592 77500
rect 168438 77500 168466 77868
rect 168880 77800 168886 77852
rect 168938 77840 168944 77852
rect 168938 77800 168972 77840
rect 168944 77648 168972 77800
rect 168926 77596 168932 77648
rect 168984 77596 168990 77648
rect 169496 77636 169524 77880
rect 169616 77868 169622 77920
rect 169674 77868 169680 77920
rect 169984 77868 169990 77920
rect 170042 77868 170048 77920
rect 169634 77772 169662 77868
rect 169708 77800 169714 77852
rect 169766 77800 169772 77852
rect 169588 77744 169662 77772
rect 169588 77716 169616 77744
rect 169726 77716 169754 77800
rect 170002 77716 170030 77868
rect 170278 77784 170306 78288
rect 174630 78276 174636 78288
rect 174688 78276 174694 78328
rect 174722 78248 174728 78260
rect 171106 78220 174728 78248
rect 170352 77868 170358 77920
rect 170410 77868 170416 77920
rect 170720 77868 170726 77920
rect 170778 77908 170784 77920
rect 171106 77908 171134 78220
rect 174722 78208 174728 78220
rect 174780 78208 174786 78260
rect 174814 78180 174820 78192
rect 171198 78152 174820 78180
rect 171198 77920 171226 78152
rect 174814 78140 174820 78152
rect 174872 78140 174878 78192
rect 180058 78112 180064 78124
rect 171290 78084 180064 78112
rect 171290 77920 171318 78084
rect 180058 78072 180064 78084
rect 180116 78072 180122 78124
rect 183526 78084 186314 78112
rect 183526 78044 183554 78084
rect 171382 78016 183554 78044
rect 186286 78044 186314 78084
rect 393958 78044 393964 78056
rect 186286 78016 393964 78044
rect 171382 77920 171410 78016
rect 393958 78004 393964 78016
rect 394016 78004 394022 78056
rect 174630 77976 174636 77988
rect 172026 77948 173618 77976
rect 172026 77920 172054 77948
rect 170778 77880 171134 77908
rect 170778 77868 170784 77880
rect 171180 77868 171186 77920
rect 171238 77868 171244 77920
rect 171272 77868 171278 77920
rect 171330 77868 171336 77920
rect 171364 77868 171370 77920
rect 171422 77868 171428 77920
rect 171732 77868 171738 77920
rect 171790 77908 171796 77920
rect 171916 77908 171922 77920
rect 171790 77868 171824 77908
rect 170370 77840 170398 77868
rect 170370 77812 170720 77840
rect 170692 77784 170720 77812
rect 171088 77800 171094 77852
rect 171146 77800 171152 77852
rect 170278 77744 170312 77784
rect 170306 77732 170312 77744
rect 170364 77732 170370 77784
rect 170674 77732 170680 77784
rect 170732 77732 170738 77784
rect 171106 77772 171134 77800
rect 171106 77744 171732 77772
rect 169570 77664 169576 77716
rect 169628 77664 169634 77716
rect 169662 77664 169668 77716
rect 169720 77676 169754 77716
rect 169720 77664 169726 77676
rect 169984 77664 169990 77716
rect 170042 77664 170048 77716
rect 171704 77648 171732 77744
rect 171796 77648 171824 77868
rect 171888 77868 171922 77908
rect 171974 77868 171980 77920
rect 172008 77868 172014 77920
rect 172066 77868 172072 77920
rect 173020 77868 173026 77920
rect 173078 77868 173084 77920
rect 170398 77636 170404 77648
rect 169496 77608 170404 77636
rect 170398 77596 170404 77608
rect 170456 77596 170462 77648
rect 171686 77596 171692 77648
rect 171744 77596 171750 77648
rect 171778 77596 171784 77648
rect 171836 77596 171842 77648
rect 171502 77528 171508 77580
rect 171560 77568 171566 77580
rect 171888 77568 171916 77868
rect 173038 77772 173066 77868
rect 173590 77840 173618 77948
rect 173682 77948 174636 77976
rect 173682 77920 173710 77948
rect 174630 77936 174636 77948
rect 174688 77936 174694 77988
rect 580350 77976 580356 77988
rect 176028 77948 580356 77976
rect 173664 77868 173670 77920
rect 173722 77868 173728 77920
rect 173756 77868 173762 77920
rect 173814 77908 173820 77920
rect 174538 77908 174544 77920
rect 173814 77880 174544 77908
rect 173814 77868 173820 77880
rect 174538 77868 174544 77880
rect 174596 77868 174602 77920
rect 176028 77840 176056 77948
rect 580350 77936 580356 77948
rect 580408 77936 580414 77988
rect 173590 77812 176056 77840
rect 176102 77800 176108 77852
rect 176160 77840 176166 77852
rect 396902 77840 396908 77852
rect 176160 77812 396908 77840
rect 176160 77800 176166 77812
rect 396902 77800 396908 77812
rect 396960 77800 396966 77852
rect 171980 77744 173066 77772
rect 171980 77716 172008 77744
rect 171962 77664 171968 77716
rect 172020 77664 172026 77716
rect 172100 77664 172106 77716
rect 172158 77704 172164 77716
rect 175826 77704 175832 77716
rect 172158 77676 175832 77704
rect 172158 77664 172164 77676
rect 175826 77664 175832 77676
rect 175884 77664 175890 77716
rect 175918 77664 175924 77716
rect 175976 77704 175982 77716
rect 231854 77704 231860 77716
rect 175976 77676 231860 77704
rect 175976 77664 175982 77676
rect 231854 77664 231860 77676
rect 231912 77664 231918 77716
rect 172238 77596 172244 77648
rect 172296 77636 172302 77648
rect 172296 77608 173480 77636
rect 172296 77596 172302 77608
rect 171560 77540 171916 77568
rect 171560 77528 171566 77540
rect 172054 77528 172060 77580
rect 172112 77568 172118 77580
rect 173452 77568 173480 77608
rect 173618 77596 173624 77648
rect 173676 77636 173682 77648
rect 200114 77636 200120 77648
rect 173676 77608 200120 77636
rect 173676 77596 173682 77608
rect 200114 77596 200120 77608
rect 200172 77596 200178 77648
rect 175826 77568 175832 77580
rect 172112 77540 172284 77568
rect 173452 77540 175832 77568
rect 172112 77528 172118 77540
rect 168558 77500 168564 77512
rect 168438 77472 168564 77500
rect 166960 77460 166966 77472
rect 168558 77460 168564 77472
rect 168616 77460 168622 77512
rect 172256 77500 172284 77540
rect 175826 77528 175832 77540
rect 175884 77528 175890 77580
rect 175918 77528 175924 77580
rect 175976 77568 175982 77580
rect 284294 77568 284300 77580
rect 175976 77540 284300 77568
rect 175976 77528 175982 77540
rect 284294 77528 284300 77540
rect 284352 77528 284358 77580
rect 252554 77500 252560 77512
rect 172256 77472 252560 77500
rect 252554 77460 252560 77472
rect 252612 77460 252618 77512
rect 167546 77392 167552 77444
rect 167604 77432 167610 77444
rect 172054 77432 172060 77444
rect 167604 77404 172060 77432
rect 167604 77392 167610 77404
rect 172054 77392 172060 77404
rect 172112 77392 172118 77444
rect 172238 77392 172244 77444
rect 172296 77432 172302 77444
rect 302234 77432 302240 77444
rect 172296 77404 302240 77432
rect 172296 77392 172302 77404
rect 302234 77392 302240 77404
rect 302292 77392 302298 77444
rect 165430 77364 165436 77376
rect 162688 77336 165436 77364
rect 165430 77324 165436 77336
rect 165488 77324 165494 77376
rect 165798 77324 165804 77376
rect 165856 77364 165862 77376
rect 320174 77364 320180 77376
rect 165856 77336 320180 77364
rect 165856 77324 165862 77336
rect 320174 77324 320180 77336
rect 320232 77324 320238 77376
rect 158496 77268 160048 77296
rect 158496 77256 158502 77268
rect 161566 77256 161572 77308
rect 161624 77296 161630 77308
rect 462406 77296 462412 77308
rect 161624 77268 462412 77296
rect 161624 77256 161630 77268
rect 462406 77256 462412 77268
rect 462464 77256 462470 77308
rect 147582 77228 147588 77240
rect 144702 77200 147588 77228
rect 141016 77188 141022 77200
rect 147582 77188 147588 77200
rect 147640 77188 147646 77240
rect 149146 77188 149152 77240
rect 149204 77228 149210 77240
rect 162946 77228 162952 77240
rect 149204 77200 162952 77228
rect 149204 77188 149210 77200
rect 162946 77188 162952 77200
rect 163004 77188 163010 77240
rect 163590 77188 163596 77240
rect 163648 77228 163654 77240
rect 170306 77228 170312 77240
rect 163648 77200 170312 77228
rect 163648 77188 163654 77200
rect 170306 77188 170312 77200
rect 170364 77188 170370 77240
rect 171686 77188 171692 77240
rect 171744 77228 171750 77240
rect 171744 77200 179414 77228
rect 171744 77188 171750 77200
rect 116578 77120 116584 77172
rect 116636 77160 116642 77172
rect 171962 77160 171968 77172
rect 116636 77132 171968 77160
rect 116636 77120 116642 77132
rect 171962 77120 171968 77132
rect 172020 77120 172026 77172
rect 179386 77160 179414 77200
rect 180242 77160 180248 77172
rect 179386 77132 180248 77160
rect 180242 77120 180248 77132
rect 180300 77120 180306 77172
rect 116670 77052 116676 77104
rect 116728 77092 116734 77104
rect 173986 77092 173992 77104
rect 116728 77064 173992 77092
rect 116728 77052 116734 77064
rect 173986 77052 173992 77064
rect 174044 77052 174050 77104
rect 120718 76984 120724 77036
rect 120776 77024 120782 77036
rect 174170 77024 174176 77036
rect 120776 76996 174176 77024
rect 120776 76984 120782 76996
rect 174170 76984 174176 76996
rect 174228 76984 174234 77036
rect 142246 76916 142252 76968
rect 142304 76956 142310 76968
rect 213914 76956 213920 76968
rect 142304 76928 213920 76956
rect 142304 76916 142310 76928
rect 213914 76916 213920 76928
rect 213972 76916 213978 76968
rect 144270 76848 144276 76900
rect 144328 76888 144334 76900
rect 144546 76888 144552 76900
rect 144328 76860 144552 76888
rect 144328 76848 144334 76860
rect 144546 76848 144552 76860
rect 144604 76848 144610 76900
rect 146938 76848 146944 76900
rect 146996 76888 147002 76900
rect 267734 76888 267740 76900
rect 146996 76860 162946 76888
rect 146996 76848 147002 76860
rect 118666 76792 138014 76820
rect 4982 76576 4988 76628
rect 5040 76616 5046 76628
rect 118666 76616 118694 76792
rect 124766 76712 124772 76764
rect 124824 76752 124830 76764
rect 130930 76752 130936 76764
rect 124824 76724 130936 76752
rect 124824 76712 124830 76724
rect 130930 76712 130936 76724
rect 130988 76712 130994 76764
rect 5040 76588 118694 76616
rect 137986 76616 138014 76792
rect 147582 76780 147588 76832
rect 147640 76820 147646 76832
rect 151998 76820 152004 76832
rect 147640 76792 152004 76820
rect 147640 76780 147646 76792
rect 151998 76780 152004 76792
rect 152056 76780 152062 76832
rect 155310 76780 155316 76832
rect 155368 76820 155374 76832
rect 162670 76820 162676 76832
rect 155368 76792 162676 76820
rect 155368 76780 155374 76792
rect 162670 76780 162676 76792
rect 162728 76780 162734 76832
rect 162918 76820 162946 76860
rect 163378 76860 267740 76888
rect 162918 76792 163084 76820
rect 158622 76712 158628 76764
rect 158680 76752 158686 76764
rect 163056 76752 163084 76792
rect 163378 76752 163406 76860
rect 267734 76848 267740 76860
rect 267792 76848 267798 76900
rect 165522 76780 165528 76832
rect 165580 76820 165586 76832
rect 306374 76820 306380 76832
rect 165580 76792 306380 76820
rect 165580 76780 165586 76792
rect 306374 76780 306380 76792
rect 306432 76780 306438 76832
rect 166994 76752 167000 76764
rect 158680 76724 161474 76752
rect 163056 76724 163406 76752
rect 163470 76724 167000 76752
rect 158680 76712 158686 76724
rect 154666 76644 154672 76696
rect 154724 76684 154730 76696
rect 155310 76684 155316 76696
rect 154724 76656 155316 76684
rect 154724 76644 154730 76656
rect 155310 76644 155316 76656
rect 155368 76644 155374 76696
rect 155678 76644 155684 76696
rect 155736 76684 155742 76696
rect 156138 76684 156144 76696
rect 155736 76656 156144 76684
rect 155736 76644 155742 76656
rect 156138 76644 156144 76656
rect 156196 76644 156202 76696
rect 157518 76644 157524 76696
rect 157576 76684 157582 76696
rect 158714 76684 158720 76696
rect 157576 76656 158720 76684
rect 157576 76644 157582 76656
rect 158714 76644 158720 76656
rect 158772 76644 158778 76696
rect 137986 76588 150434 76616
rect 5040 76576 5046 76588
rect 121362 76440 121368 76492
rect 121420 76480 121426 76492
rect 126974 76480 126980 76492
rect 121420 76452 126980 76480
rect 121420 76440 121426 76452
rect 126974 76440 126980 76452
rect 127032 76440 127038 76492
rect 146294 76480 146300 76492
rect 146220 76452 146300 76480
rect 125778 76304 125784 76356
rect 125836 76344 125842 76356
rect 126146 76344 126152 76356
rect 125836 76316 126152 76344
rect 125836 76304 125842 76316
rect 126146 76304 126152 76316
rect 126204 76304 126210 76356
rect 127250 76304 127256 76356
rect 127308 76344 127314 76356
rect 127618 76344 127624 76356
rect 127308 76316 127624 76344
rect 127308 76304 127314 76316
rect 127618 76304 127624 76316
rect 127676 76304 127682 76356
rect 129826 76304 129832 76356
rect 129884 76344 129890 76356
rect 130102 76344 130108 76356
rect 129884 76316 130108 76344
rect 129884 76304 129890 76316
rect 130102 76304 130108 76316
rect 130160 76304 130166 76356
rect 130286 76304 130292 76356
rect 130344 76344 130350 76356
rect 130746 76344 130752 76356
rect 130344 76316 130752 76344
rect 130344 76304 130350 76316
rect 130746 76304 130752 76316
rect 130804 76304 130810 76356
rect 130010 76236 130016 76288
rect 130068 76276 130074 76288
rect 130470 76276 130476 76288
rect 130068 76248 130476 76276
rect 130068 76236 130074 76248
rect 130470 76236 130476 76248
rect 130528 76236 130534 76288
rect 127618 76168 127624 76220
rect 127676 76208 127682 76220
rect 129090 76208 129096 76220
rect 127676 76180 129096 76208
rect 127676 76168 127682 76180
rect 129090 76168 129096 76180
rect 129148 76168 129154 76220
rect 126054 76100 126060 76152
rect 126112 76140 126118 76152
rect 126238 76140 126244 76152
rect 126112 76112 126244 76140
rect 126112 76100 126118 76112
rect 126238 76100 126244 76112
rect 126296 76100 126302 76152
rect 146220 76072 146248 76452
rect 146294 76440 146300 76452
rect 146352 76440 146358 76492
rect 150406 76480 150434 76588
rect 152366 76576 152372 76628
rect 152424 76616 152430 76628
rect 161198 76616 161204 76628
rect 152424 76588 161204 76616
rect 152424 76576 152430 76588
rect 161198 76576 161204 76588
rect 161256 76576 161262 76628
rect 161446 76616 161474 76724
rect 162210 76644 162216 76696
rect 162268 76684 162274 76696
rect 163470 76684 163498 76724
rect 166994 76712 167000 76724
rect 167052 76712 167058 76764
rect 168650 76712 168656 76764
rect 168708 76752 168714 76764
rect 170766 76752 170772 76764
rect 168708 76724 170772 76752
rect 168708 76712 168714 76724
rect 170766 76712 170772 76724
rect 170824 76712 170830 76764
rect 171134 76712 171140 76764
rect 171192 76752 171198 76764
rect 175918 76752 175924 76764
rect 171192 76724 175924 76752
rect 171192 76712 171198 76724
rect 175918 76712 175924 76724
rect 175976 76712 175982 76764
rect 178402 76712 178408 76764
rect 178460 76752 178466 76764
rect 431954 76752 431960 76764
rect 178460 76724 431960 76752
rect 178460 76712 178466 76724
rect 431954 76712 431960 76724
rect 432012 76712 432018 76764
rect 426434 76684 426440 76696
rect 162268 76656 163498 76684
rect 164160 76656 426440 76684
rect 162268 76644 162274 76656
rect 164160 76616 164188 76656
rect 426434 76644 426440 76656
rect 426492 76644 426498 76696
rect 171042 76616 171048 76628
rect 161446 76588 164188 76616
rect 164252 76588 171048 76616
rect 156138 76508 156144 76560
rect 156196 76548 156202 76560
rect 156782 76548 156788 76560
rect 156196 76520 156788 76548
rect 156196 76508 156202 76520
rect 156782 76508 156788 76520
rect 156840 76508 156846 76560
rect 160094 76508 160100 76560
rect 160152 76548 160158 76560
rect 164252 76548 164280 76588
rect 171042 76576 171048 76588
rect 171100 76576 171106 76628
rect 171318 76576 171324 76628
rect 171376 76616 171382 76628
rect 176102 76616 176108 76628
rect 171376 76588 176108 76616
rect 171376 76576 171382 76588
rect 176102 76576 176108 76588
rect 176160 76576 176166 76628
rect 176194 76576 176200 76628
rect 176252 76616 176258 76628
rect 462314 76616 462320 76628
rect 176252 76588 462320 76616
rect 176252 76576 176258 76588
rect 462314 76576 462320 76588
rect 462372 76576 462378 76628
rect 160152 76520 164280 76548
rect 160152 76508 160158 76520
rect 164326 76508 164332 76560
rect 164384 76548 164390 76560
rect 168742 76548 168748 76560
rect 164384 76520 168748 76548
rect 164384 76508 164390 76520
rect 168742 76508 168748 76520
rect 168800 76508 168806 76560
rect 170398 76508 170404 76560
rect 170456 76548 170462 76560
rect 557534 76548 557540 76560
rect 170456 76520 557540 76548
rect 170456 76508 170462 76520
rect 557534 76508 557540 76520
rect 557592 76508 557598 76560
rect 150406 76452 162854 76480
rect 156414 76372 156420 76424
rect 156472 76412 156478 76424
rect 156782 76412 156788 76424
rect 156472 76384 156788 76412
rect 156472 76372 156478 76384
rect 156782 76372 156788 76384
rect 156840 76372 156846 76424
rect 146294 76304 146300 76356
rect 146352 76344 146358 76356
rect 146846 76344 146852 76356
rect 146352 76316 146852 76344
rect 146352 76304 146358 76316
rect 146846 76304 146852 76316
rect 146904 76304 146910 76356
rect 161566 76304 161572 76356
rect 161624 76344 161630 76356
rect 161934 76344 161940 76356
rect 161624 76316 161940 76344
rect 161624 76304 161630 76316
rect 161934 76304 161940 76316
rect 161992 76304 161998 76356
rect 156046 76236 156052 76288
rect 156104 76276 156110 76288
rect 156414 76276 156420 76288
rect 156104 76248 156420 76276
rect 156104 76236 156110 76248
rect 156414 76236 156420 76248
rect 156472 76236 156478 76288
rect 162826 76276 162854 76452
rect 164234 76440 164240 76492
rect 164292 76480 164298 76492
rect 165338 76480 165344 76492
rect 164292 76452 165344 76480
rect 164292 76440 164298 76452
rect 165338 76440 165344 76452
rect 165396 76440 165402 76492
rect 167270 76440 167276 76492
rect 167328 76480 167334 76492
rect 168098 76480 168104 76492
rect 167328 76452 168104 76480
rect 167328 76440 167334 76452
rect 168098 76440 168104 76452
rect 168156 76440 168162 76492
rect 168650 76440 168656 76492
rect 168708 76480 168714 76492
rect 169386 76480 169392 76492
rect 168708 76452 169392 76480
rect 168708 76440 168714 76452
rect 169386 76440 169392 76452
rect 169444 76440 169450 76492
rect 171962 76440 171968 76492
rect 172020 76480 172026 76492
rect 173894 76480 173900 76492
rect 172020 76452 173900 76480
rect 172020 76440 172026 76452
rect 173894 76440 173900 76452
rect 173952 76440 173958 76492
rect 163038 76372 163044 76424
rect 163096 76412 163102 76424
rect 172054 76412 172060 76424
rect 163096 76384 172060 76412
rect 163096 76372 163102 76384
rect 172054 76372 172060 76384
rect 172112 76372 172118 76424
rect 172330 76372 172336 76424
rect 172388 76412 172394 76424
rect 175826 76412 175832 76424
rect 172388 76384 175832 76412
rect 172388 76372 172394 76384
rect 175826 76372 175832 76384
rect 175884 76372 175890 76424
rect 162946 76304 162952 76356
rect 163004 76344 163010 76356
rect 172238 76344 172244 76356
rect 163004 76316 172244 76344
rect 163004 76304 163010 76316
rect 172238 76304 172244 76316
rect 172296 76304 172302 76356
rect 174354 76276 174360 76288
rect 162826 76248 174360 76276
rect 174354 76236 174360 76248
rect 174412 76236 174418 76288
rect 146570 76168 146576 76220
rect 146628 76208 146634 76220
rect 147306 76208 147312 76220
rect 146628 76180 147312 76208
rect 146628 76168 146634 76180
rect 147306 76168 147312 76180
rect 147364 76168 147370 76220
rect 159542 76168 159548 76220
rect 159600 76208 159606 76220
rect 159910 76208 159916 76220
rect 159600 76180 159916 76208
rect 159600 76168 159606 76180
rect 159910 76168 159916 76180
rect 159968 76168 159974 76220
rect 161934 76168 161940 76220
rect 161992 76208 161998 76220
rect 165798 76208 165804 76220
rect 161992 76180 165804 76208
rect 161992 76168 161998 76180
rect 165798 76168 165804 76180
rect 165856 76168 165862 76220
rect 171134 76168 171140 76220
rect 171192 76208 171198 76220
rect 172698 76208 172704 76220
rect 171192 76180 172704 76208
rect 171192 76168 171198 76180
rect 172698 76168 172704 76180
rect 172756 76168 172762 76220
rect 146386 76100 146392 76152
rect 146444 76140 146450 76152
rect 146754 76140 146760 76152
rect 146444 76112 146760 76140
rect 146444 76100 146450 76112
rect 146754 76100 146760 76112
rect 146812 76100 146818 76152
rect 147674 76100 147680 76152
rect 147732 76140 147738 76152
rect 150158 76140 150164 76152
rect 147732 76112 150164 76140
rect 147732 76100 147738 76112
rect 150158 76100 150164 76112
rect 150216 76100 150222 76152
rect 153102 76100 153108 76152
rect 153160 76140 153166 76152
rect 158530 76140 158536 76152
rect 153160 76112 158536 76140
rect 153160 76100 153166 76112
rect 158530 76100 158536 76112
rect 158588 76100 158594 76152
rect 160462 76100 160468 76152
rect 160520 76140 160526 76152
rect 167546 76140 167552 76152
rect 160520 76112 167552 76140
rect 160520 76100 160526 76112
rect 167546 76100 167552 76112
rect 167604 76100 167610 76152
rect 168006 76100 168012 76152
rect 168064 76140 168070 76152
rect 169386 76140 169392 76152
rect 168064 76112 169392 76140
rect 168064 76100 168070 76112
rect 169386 76100 169392 76112
rect 169444 76100 169450 76152
rect 146570 76072 146576 76084
rect 146220 76044 146576 76072
rect 146570 76032 146576 76044
rect 146628 76032 146634 76084
rect 159174 76032 159180 76084
rect 159232 76072 159238 76084
rect 159910 76072 159916 76084
rect 159232 76044 159916 76072
rect 159232 76032 159238 76044
rect 159910 76032 159916 76044
rect 159968 76032 159974 76084
rect 160094 76032 160100 76084
rect 160152 76072 160158 76084
rect 195974 76072 195980 76084
rect 160152 76044 195980 76072
rect 160152 76032 160158 76044
rect 195974 76032 195980 76044
rect 196032 76032 196038 76084
rect 148594 75964 148600 76016
rect 148652 76004 148658 76016
rect 155586 76004 155592 76016
rect 148652 75976 155592 76004
rect 148652 75964 148658 75976
rect 155586 75964 155592 75976
rect 155644 75964 155650 76016
rect 157426 75964 157432 76016
rect 157484 76004 157490 76016
rect 158346 76004 158352 76016
rect 157484 75976 158352 76004
rect 157484 75964 157490 75976
rect 158346 75964 158352 75976
rect 158404 75964 158410 76016
rect 161566 75964 161572 76016
rect 161624 76004 161630 76016
rect 161750 76004 161756 76016
rect 161624 75976 161756 76004
rect 161624 75964 161630 75976
rect 161750 75964 161756 75976
rect 161808 75964 161814 76016
rect 165798 75964 165804 76016
rect 165856 76004 165862 76016
rect 249794 76004 249800 76016
rect 165856 75976 249800 76004
rect 165856 75964 165862 75976
rect 249794 75964 249800 75976
rect 249852 75964 249858 76016
rect 129182 75936 129188 75948
rect 121426 75908 129188 75936
rect 121086 75828 121092 75880
rect 121144 75868 121150 75880
rect 121426 75868 121454 75908
rect 129182 75896 129188 75908
rect 129240 75896 129246 75948
rect 152826 75896 152832 75948
rect 152884 75936 152890 75948
rect 154114 75936 154120 75948
rect 152884 75908 154120 75936
rect 152884 75896 152890 75908
rect 154114 75896 154120 75908
rect 154172 75896 154178 75948
rect 157150 75896 157156 75948
rect 157208 75936 157214 75948
rect 157518 75936 157524 75948
rect 157208 75908 157524 75936
rect 157208 75896 157214 75908
rect 157518 75896 157524 75908
rect 157576 75896 157582 75948
rect 159174 75896 159180 75948
rect 159232 75936 159238 75948
rect 159358 75936 159364 75948
rect 159232 75908 159364 75936
rect 159232 75896 159238 75908
rect 159358 75896 159364 75908
rect 159416 75896 159422 75948
rect 162118 75896 162124 75948
rect 162176 75936 162182 75948
rect 288434 75936 288440 75948
rect 162176 75908 288440 75936
rect 162176 75896 162182 75908
rect 288434 75896 288440 75908
rect 288492 75896 288498 75948
rect 121144 75840 121454 75868
rect 121144 75828 121150 75840
rect 153470 75828 153476 75880
rect 153528 75868 153534 75880
rect 153930 75868 153936 75880
rect 153528 75840 153936 75868
rect 153528 75828 153534 75840
rect 153930 75828 153936 75840
rect 153988 75828 153994 75880
rect 154666 75828 154672 75880
rect 154724 75868 154730 75880
rect 155126 75868 155132 75880
rect 154724 75840 155132 75868
rect 154724 75828 154730 75840
rect 155126 75828 155132 75840
rect 155184 75828 155190 75880
rect 155954 75828 155960 75880
rect 156012 75868 156018 75880
rect 156322 75868 156328 75880
rect 156012 75840 156328 75868
rect 156012 75828 156018 75840
rect 156322 75828 156328 75840
rect 156380 75828 156386 75880
rect 156690 75828 156696 75880
rect 156748 75868 156754 75880
rect 161934 75868 161940 75880
rect 156748 75840 161940 75868
rect 156748 75828 156754 75840
rect 161934 75828 161940 75840
rect 161992 75828 161998 75880
rect 164878 75868 164884 75880
rect 163516 75840 164884 75868
rect 125226 75760 125232 75812
rect 125284 75800 125290 75812
rect 133506 75800 133512 75812
rect 125284 75772 133512 75800
rect 125284 75760 125290 75772
rect 133506 75760 133512 75772
rect 133564 75760 133570 75812
rect 141142 75760 141148 75812
rect 141200 75800 141206 75812
rect 163516 75800 163544 75840
rect 164878 75828 164884 75840
rect 164936 75828 164942 75880
rect 168346 75840 168742 75868
rect 141200 75772 163544 75800
rect 141200 75760 141206 75772
rect 163866 75760 163872 75812
rect 163924 75800 163930 75812
rect 164050 75800 164056 75812
rect 163924 75772 164056 75800
rect 163924 75760 163930 75772
rect 164050 75760 164056 75772
rect 164108 75760 164114 75812
rect 168346 75800 168374 75840
rect 164252 75772 168374 75800
rect 128538 75692 128544 75744
rect 128596 75732 128602 75744
rect 129366 75732 129372 75744
rect 128596 75704 129372 75732
rect 128596 75692 128602 75704
rect 129366 75692 129372 75704
rect 129424 75692 129430 75744
rect 139394 75692 139400 75744
rect 139452 75732 139458 75744
rect 164252 75732 164280 75772
rect 165798 75732 165804 75744
rect 139452 75704 164280 75732
rect 164390 75704 165804 75732
rect 139452 75692 139458 75704
rect 143626 75624 143632 75676
rect 143684 75664 143690 75676
rect 144086 75664 144092 75676
rect 143684 75636 144092 75664
rect 143684 75624 143690 75636
rect 144086 75624 144092 75636
rect 144144 75624 144150 75676
rect 145006 75624 145012 75676
rect 145064 75664 145070 75676
rect 164390 75664 164418 75704
rect 165798 75692 165804 75704
rect 165856 75692 165862 75744
rect 167914 75692 167920 75744
rect 167972 75732 167978 75744
rect 168098 75732 168104 75744
rect 167972 75704 168104 75732
rect 167972 75692 167978 75704
rect 168098 75692 168104 75704
rect 168156 75692 168162 75744
rect 168714 75732 168742 75840
rect 169018 75760 169024 75812
rect 169076 75800 169082 75812
rect 169662 75800 169668 75812
rect 169076 75772 169668 75800
rect 169076 75760 169082 75772
rect 169662 75760 169668 75772
rect 169720 75760 169726 75812
rect 172606 75760 172612 75812
rect 172664 75800 172670 75812
rect 284938 75800 284944 75812
rect 172664 75772 284944 75800
rect 172664 75760 172670 75772
rect 284938 75760 284944 75772
rect 284996 75760 285002 75812
rect 173158 75732 173164 75744
rect 168714 75704 173164 75732
rect 173158 75692 173164 75704
rect 173216 75692 173222 75744
rect 145064 75636 164418 75664
rect 145064 75624 145070 75636
rect 164510 75624 164516 75676
rect 164568 75664 164574 75676
rect 165522 75664 165528 75676
rect 164568 75636 165528 75664
rect 164568 75624 164574 75636
rect 165522 75624 165528 75636
rect 165580 75624 165586 75676
rect 167454 75624 167460 75676
rect 167512 75664 167518 75676
rect 167730 75664 167736 75676
rect 167512 75636 167736 75664
rect 167512 75624 167518 75636
rect 167730 75624 167736 75636
rect 167788 75624 167794 75676
rect 169018 75624 169024 75676
rect 169076 75664 169082 75676
rect 169478 75664 169484 75676
rect 169076 75636 169484 75664
rect 169076 75624 169082 75636
rect 169478 75624 169484 75636
rect 169536 75624 169542 75676
rect 169938 75624 169944 75676
rect 169996 75664 170002 75676
rect 170122 75664 170128 75676
rect 169996 75636 170128 75664
rect 169996 75624 170002 75636
rect 170122 75624 170128 75636
rect 170180 75624 170186 75676
rect 145190 75556 145196 75608
rect 145248 75596 145254 75608
rect 150434 75596 150440 75608
rect 145248 75568 150440 75596
rect 145248 75556 145254 75568
rect 150434 75556 150440 75568
rect 150492 75556 150498 75608
rect 150710 75556 150716 75608
rect 150768 75596 150774 75608
rect 151078 75596 151084 75608
rect 150768 75568 151084 75596
rect 150768 75556 150774 75568
rect 151078 75556 151084 75568
rect 151136 75556 151142 75608
rect 153470 75556 153476 75608
rect 153528 75596 153534 75608
rect 153746 75596 153752 75608
rect 153528 75568 153752 75596
rect 153528 75556 153534 75568
rect 153746 75556 153752 75568
rect 153804 75556 153810 75608
rect 153838 75556 153844 75608
rect 153896 75556 153902 75608
rect 155126 75556 155132 75608
rect 155184 75596 155190 75608
rect 155770 75596 155776 75608
rect 155184 75568 155776 75596
rect 155184 75556 155190 75568
rect 155770 75556 155776 75568
rect 155828 75556 155834 75608
rect 157334 75556 157340 75608
rect 157392 75596 157398 75608
rect 157886 75596 157892 75608
rect 157392 75568 157892 75596
rect 157392 75556 157398 75568
rect 157886 75556 157892 75568
rect 157944 75556 157950 75608
rect 158438 75556 158444 75608
rect 158496 75596 158502 75608
rect 159358 75596 159364 75608
rect 158496 75568 159364 75596
rect 158496 75556 158502 75568
rect 159358 75556 159364 75568
rect 159416 75556 159422 75608
rect 160278 75556 160284 75608
rect 160336 75596 160342 75608
rect 160462 75596 160468 75608
rect 160336 75568 160468 75596
rect 160336 75556 160342 75568
rect 160462 75556 160468 75568
rect 160520 75556 160526 75608
rect 160646 75556 160652 75608
rect 160704 75596 160710 75608
rect 242158 75596 242164 75608
rect 160704 75568 242164 75596
rect 160704 75556 160710 75568
rect 242158 75556 242164 75568
rect 242216 75556 242222 75608
rect 149146 75488 149152 75540
rect 149204 75528 149210 75540
rect 149882 75528 149888 75540
rect 149204 75500 149888 75528
rect 149204 75488 149210 75500
rect 149882 75488 149888 75500
rect 149940 75488 149946 75540
rect 150526 75488 150532 75540
rect 150584 75528 150590 75540
rect 150894 75528 150900 75540
rect 150584 75500 150900 75528
rect 150584 75488 150590 75500
rect 150894 75488 150900 75500
rect 150952 75488 150958 75540
rect 152918 75488 152924 75540
rect 152976 75528 152982 75540
rect 153856 75528 153884 75556
rect 152976 75500 153884 75528
rect 152976 75488 152982 75500
rect 154942 75488 154948 75540
rect 155000 75528 155006 75540
rect 155000 75500 157380 75528
rect 155000 75488 155006 75500
rect 155678 75420 155684 75472
rect 155736 75460 155742 75472
rect 156414 75460 156420 75472
rect 155736 75432 156420 75460
rect 155736 75420 155742 75432
rect 156414 75420 156420 75432
rect 156472 75420 156478 75472
rect 156598 75420 156604 75472
rect 156656 75460 156662 75472
rect 156874 75460 156880 75472
rect 156656 75432 156880 75460
rect 156656 75420 156662 75432
rect 156874 75420 156880 75432
rect 156932 75420 156938 75472
rect 157352 75460 157380 75500
rect 157426 75488 157432 75540
rect 157484 75528 157490 75540
rect 157978 75528 157984 75540
rect 157484 75500 157984 75528
rect 157484 75488 157490 75500
rect 157978 75488 157984 75500
rect 158036 75488 158042 75540
rect 158714 75488 158720 75540
rect 158772 75528 158778 75540
rect 158772 75500 161336 75528
rect 158772 75488 158778 75500
rect 161308 75472 161336 75500
rect 162394 75488 162400 75540
rect 162452 75528 162458 75540
rect 162452 75500 171134 75528
rect 162452 75488 162458 75500
rect 157352 75432 158300 75460
rect 110414 75352 110420 75404
rect 110472 75392 110478 75404
rect 133966 75392 133972 75404
rect 110472 75364 133972 75392
rect 110472 75352 110478 75364
rect 133966 75352 133972 75364
rect 134024 75352 134030 75404
rect 140406 75352 140412 75404
rect 140464 75392 140470 75404
rect 148594 75392 148600 75404
rect 140464 75364 148600 75392
rect 140464 75352 140470 75364
rect 148594 75352 148600 75364
rect 148652 75352 148658 75404
rect 153286 75352 153292 75404
rect 153344 75392 153350 75404
rect 153746 75392 153752 75404
rect 153344 75364 153752 75392
rect 153344 75352 153350 75364
rect 153746 75352 153752 75364
rect 153804 75352 153810 75404
rect 57238 75284 57244 75336
rect 57296 75324 57302 75336
rect 127434 75324 127440 75336
rect 57296 75296 127440 75324
rect 57296 75284 57302 75296
rect 127434 75284 127440 75296
rect 127492 75284 127498 75336
rect 128722 75284 128728 75336
rect 128780 75324 128786 75336
rect 129550 75324 129556 75336
rect 128780 75296 129556 75324
rect 128780 75284 128786 75296
rect 129550 75284 129556 75296
rect 129608 75284 129614 75336
rect 130102 75284 130108 75336
rect 130160 75324 130166 75336
rect 130654 75324 130660 75336
rect 130160 75296 130660 75324
rect 130160 75284 130166 75296
rect 130654 75284 130660 75296
rect 130712 75284 130718 75336
rect 143718 75284 143724 75336
rect 143776 75324 143782 75336
rect 143994 75324 144000 75336
rect 143776 75296 144000 75324
rect 143776 75284 143782 75296
rect 143994 75284 144000 75296
rect 144052 75284 144058 75336
rect 157610 75284 157616 75336
rect 157668 75324 157674 75336
rect 157886 75324 157892 75336
rect 157668 75296 157892 75324
rect 157668 75284 157674 75296
rect 157886 75284 157892 75296
rect 157944 75284 157950 75336
rect 158272 75324 158300 75432
rect 160278 75420 160284 75472
rect 160336 75460 160342 75472
rect 160554 75460 160560 75472
rect 160336 75432 160560 75460
rect 160336 75420 160342 75432
rect 160554 75420 160560 75432
rect 160612 75420 160618 75472
rect 161290 75420 161296 75472
rect 161348 75420 161354 75472
rect 162946 75420 162952 75472
rect 163004 75460 163010 75472
rect 163958 75460 163964 75472
rect 163004 75432 163964 75460
rect 163004 75420 163010 75432
rect 163958 75420 163964 75432
rect 164016 75420 164022 75472
rect 164142 75420 164148 75472
rect 164200 75460 164206 75472
rect 164602 75460 164608 75472
rect 164200 75432 164608 75460
rect 164200 75420 164206 75432
rect 164602 75420 164608 75432
rect 164660 75420 164666 75472
rect 171106 75460 171134 75500
rect 174722 75488 174728 75540
rect 174780 75528 174786 75540
rect 391198 75528 391204 75540
rect 174780 75500 391204 75528
rect 174780 75488 174786 75500
rect 391198 75488 391204 75500
rect 391256 75488 391262 75540
rect 471238 75460 471244 75472
rect 171106 75432 471244 75460
rect 471238 75420 471244 75432
rect 471296 75420 471302 75472
rect 158530 75352 158536 75404
rect 158588 75392 158594 75404
rect 161934 75392 161940 75404
rect 158588 75364 161940 75392
rect 158588 75352 158594 75364
rect 161934 75352 161940 75364
rect 161992 75352 161998 75404
rect 164234 75352 164240 75404
rect 164292 75392 164298 75404
rect 164786 75392 164792 75404
rect 164292 75364 164792 75392
rect 164292 75352 164298 75364
rect 164786 75352 164792 75364
rect 164844 75352 164850 75404
rect 165430 75352 165436 75404
rect 165488 75392 165494 75404
rect 478138 75392 478144 75404
rect 165488 75364 478144 75392
rect 165488 75352 165494 75364
rect 478138 75352 478144 75364
rect 478196 75352 478202 75404
rect 160554 75324 160560 75336
rect 158272 75296 160560 75324
rect 160554 75284 160560 75296
rect 160612 75284 160618 75336
rect 161658 75284 161664 75336
rect 161716 75324 161722 75336
rect 162210 75324 162216 75336
rect 161716 75296 162216 75324
rect 161716 75284 161722 75296
rect 162210 75284 162216 75296
rect 162268 75284 162274 75336
rect 163130 75284 163136 75336
rect 163188 75324 163194 75336
rect 483014 75324 483020 75336
rect 163188 75296 483020 75324
rect 163188 75284 163194 75296
rect 483014 75284 483020 75296
rect 483072 75284 483078 75336
rect 46198 75216 46204 75268
rect 46256 75256 46262 75268
rect 119798 75256 119804 75268
rect 46256 75228 119804 75256
rect 46256 75216 46262 75228
rect 119798 75216 119804 75228
rect 119856 75216 119862 75268
rect 129182 75216 129188 75268
rect 129240 75256 129246 75268
rect 130194 75256 130200 75268
rect 129240 75228 130200 75256
rect 129240 75216 129246 75228
rect 130194 75216 130200 75228
rect 130252 75216 130258 75268
rect 139210 75216 139216 75268
rect 139268 75256 139274 75268
rect 140406 75256 140412 75268
rect 139268 75228 140412 75256
rect 139268 75216 139274 75228
rect 140406 75216 140412 75228
rect 140464 75216 140470 75268
rect 140866 75216 140872 75268
rect 140924 75256 140930 75268
rect 153102 75256 153108 75268
rect 140924 75228 153108 75256
rect 140924 75216 140930 75228
rect 153102 75216 153108 75228
rect 153160 75216 153166 75268
rect 154390 75216 154396 75268
rect 154448 75256 154454 75268
rect 162394 75256 162400 75268
rect 154448 75228 162400 75256
rect 154448 75216 154454 75228
rect 162394 75216 162400 75228
rect 162452 75216 162458 75268
rect 162762 75216 162768 75268
rect 162820 75256 162826 75268
rect 163958 75256 163964 75268
rect 162820 75228 163964 75256
rect 162820 75216 162826 75228
rect 163958 75216 163964 75228
rect 164016 75216 164022 75268
rect 168742 75216 168748 75268
rect 168800 75256 168806 75268
rect 498194 75256 498200 75268
rect 168800 75228 498200 75256
rect 168800 75216 168806 75228
rect 498194 75216 498200 75228
rect 498252 75216 498258 75268
rect 22738 75148 22744 75200
rect 22796 75188 22802 75200
rect 123754 75188 123760 75200
rect 22796 75160 123760 75188
rect 22796 75148 22802 75160
rect 123754 75148 123760 75160
rect 123812 75148 123818 75200
rect 135070 75188 135076 75200
rect 126808 75160 135076 75188
rect 126808 75132 126836 75160
rect 135070 75148 135076 75160
rect 135128 75148 135134 75200
rect 137738 75148 137744 75200
rect 137796 75188 137802 75200
rect 152734 75188 152740 75200
rect 137796 75160 152740 75188
rect 137796 75148 137802 75160
rect 152734 75148 152740 75160
rect 152792 75148 152798 75200
rect 153838 75148 153844 75200
rect 153896 75188 153902 75200
rect 154022 75188 154028 75200
rect 153896 75160 154028 75188
rect 153896 75148 153902 75160
rect 154022 75148 154028 75160
rect 154080 75148 154086 75200
rect 156690 75148 156696 75200
rect 156748 75188 156754 75200
rect 156748 75160 157564 75188
rect 156748 75148 156754 75160
rect 126790 75080 126796 75132
rect 126848 75080 126854 75132
rect 127434 75080 127440 75132
rect 127492 75120 127498 75132
rect 128170 75120 128176 75132
rect 127492 75092 128176 75120
rect 127492 75080 127498 75092
rect 128170 75080 128176 75092
rect 128228 75080 128234 75132
rect 129366 75080 129372 75132
rect 129424 75120 129430 75132
rect 133874 75120 133880 75132
rect 129424 75092 133880 75120
rect 129424 75080 129430 75092
rect 133874 75080 133880 75092
rect 133932 75080 133938 75132
rect 133966 75080 133972 75132
rect 134024 75120 134030 75132
rect 136082 75120 136088 75132
rect 134024 75092 136088 75120
rect 134024 75080 134030 75092
rect 136082 75080 136088 75092
rect 136140 75080 136146 75132
rect 145006 75080 145012 75132
rect 145064 75120 145070 75132
rect 145374 75120 145380 75132
rect 145064 75092 145380 75120
rect 145064 75080 145070 75092
rect 145374 75080 145380 75092
rect 145432 75080 145438 75132
rect 149606 75080 149612 75132
rect 149664 75120 149670 75132
rect 149790 75120 149796 75132
rect 149664 75092 149796 75120
rect 149664 75080 149670 75092
rect 149790 75080 149796 75092
rect 149848 75080 149854 75132
rect 151814 75080 151820 75132
rect 151872 75120 151878 75132
rect 154482 75120 154488 75132
rect 151872 75092 154488 75120
rect 151872 75080 151878 75092
rect 154482 75080 154488 75092
rect 154540 75080 154546 75132
rect 155218 75080 155224 75132
rect 155276 75120 155282 75132
rect 157242 75120 157248 75132
rect 155276 75092 157248 75120
rect 155276 75080 155282 75092
rect 157242 75080 157248 75092
rect 157300 75080 157306 75132
rect 157536 75120 157564 75160
rect 157610 75148 157616 75200
rect 157668 75188 157674 75200
rect 158070 75188 158076 75200
rect 157668 75160 158076 75188
rect 157668 75148 157674 75160
rect 158070 75148 158076 75160
rect 158128 75148 158134 75200
rect 160370 75148 160376 75200
rect 160428 75188 160434 75200
rect 160646 75188 160652 75200
rect 160428 75160 160652 75188
rect 160428 75148 160434 75160
rect 160646 75148 160652 75160
rect 160704 75148 160710 75200
rect 161106 75148 161112 75200
rect 161164 75188 161170 75200
rect 161164 75160 168144 75188
rect 161164 75148 161170 75160
rect 164418 75120 164424 75132
rect 157536 75092 164424 75120
rect 164418 75080 164424 75092
rect 164476 75080 164482 75132
rect 164878 75080 164884 75132
rect 164936 75120 164942 75132
rect 165062 75120 165068 75132
rect 164936 75092 165068 75120
rect 164936 75080 164942 75092
rect 165062 75080 165068 75092
rect 165120 75080 165126 75132
rect 168116 75120 168144 75160
rect 169386 75148 169392 75200
rect 169444 75188 169450 75200
rect 532694 75188 532700 75200
rect 169444 75160 532700 75188
rect 169444 75148 169450 75160
rect 532694 75148 532700 75160
rect 532752 75148 532758 75200
rect 170398 75120 170404 75132
rect 168116 75092 170404 75120
rect 170398 75080 170404 75092
rect 170456 75080 170462 75132
rect 125318 75012 125324 75064
rect 125376 75052 125382 75064
rect 132954 75052 132960 75064
rect 125376 75024 132960 75052
rect 125376 75012 125382 75024
rect 132954 75012 132960 75024
rect 133012 75012 133018 75064
rect 133506 75012 133512 75064
rect 133564 75052 133570 75064
rect 135530 75052 135536 75064
rect 133564 75024 135536 75052
rect 133564 75012 133570 75024
rect 135530 75012 135536 75024
rect 135588 75012 135594 75064
rect 135714 75012 135720 75064
rect 135772 75052 135778 75064
rect 136542 75052 136548 75064
rect 135772 75024 136548 75052
rect 135772 75012 135778 75024
rect 136542 75012 136548 75024
rect 136600 75012 136606 75064
rect 137002 75052 137008 75064
rect 136652 75024 137008 75052
rect 123478 74944 123484 74996
rect 123536 74984 123542 74996
rect 134886 74984 134892 74996
rect 123536 74956 134892 74984
rect 123536 74944 123542 74956
rect 134886 74944 134892 74956
rect 134944 74944 134950 74996
rect 135070 74944 135076 74996
rect 135128 74984 135134 74996
rect 136652 74984 136680 75024
rect 137002 75012 137008 75024
rect 137060 75012 137066 75064
rect 147674 75012 147680 75064
rect 147732 75052 147738 75064
rect 148134 75052 148140 75064
rect 147732 75024 148140 75052
rect 147732 75012 147738 75024
rect 148134 75012 148140 75024
rect 148192 75012 148198 75064
rect 150434 75012 150440 75064
rect 150492 75052 150498 75064
rect 150986 75052 150992 75064
rect 150492 75024 150992 75052
rect 150492 75012 150498 75024
rect 150986 75012 150992 75024
rect 151044 75012 151050 75064
rect 158254 75012 158260 75064
rect 158312 75052 158318 75064
rect 158312 75024 166948 75052
rect 158312 75012 158318 75024
rect 135128 74956 136680 74984
rect 135128 74944 135134 74956
rect 136726 74944 136732 74996
rect 136784 74984 136790 74996
rect 137738 74984 137744 74996
rect 136784 74956 137744 74984
rect 136784 74944 136790 74956
rect 137738 74944 137744 74956
rect 137796 74944 137802 74996
rect 138658 74944 138664 74996
rect 138716 74984 138722 74996
rect 139026 74984 139032 74996
rect 138716 74956 139032 74984
rect 138716 74944 138722 74956
rect 139026 74944 139032 74956
rect 139084 74944 139090 74996
rect 143810 74944 143816 74996
rect 143868 74984 143874 74996
rect 144086 74984 144092 74996
rect 143868 74956 144092 74984
rect 143868 74944 143874 74956
rect 144086 74944 144092 74956
rect 144144 74944 144150 74996
rect 147950 74944 147956 74996
rect 148008 74984 148014 74996
rect 155218 74984 155224 74996
rect 148008 74956 155224 74984
rect 148008 74944 148014 74956
rect 155218 74944 155224 74956
rect 155276 74944 155282 74996
rect 158898 74944 158904 74996
rect 158956 74984 158962 74996
rect 159266 74984 159272 74996
rect 158956 74956 159272 74984
rect 158956 74944 158962 74956
rect 159266 74944 159272 74956
rect 159324 74944 159330 74996
rect 163222 74944 163228 74996
rect 163280 74984 163286 74996
rect 163498 74984 163504 74996
rect 163280 74956 163504 74984
rect 163280 74944 163286 74956
rect 163498 74944 163504 74956
rect 163556 74944 163562 74996
rect 166920 74984 166948 75024
rect 167546 75012 167552 75064
rect 167604 75052 167610 75064
rect 173434 75052 173440 75064
rect 167604 75024 173440 75052
rect 167604 75012 167610 75024
rect 173434 75012 173440 75024
rect 173492 75012 173498 75064
rect 173342 74984 173348 74996
rect 166920 74956 173348 74984
rect 173342 74944 173348 74956
rect 173400 74944 173406 74996
rect 127158 74876 127164 74928
rect 127216 74916 127222 74928
rect 128078 74916 128084 74928
rect 127216 74888 128084 74916
rect 127216 74876 127222 74888
rect 128078 74876 128084 74888
rect 128136 74876 128142 74928
rect 128446 74876 128452 74928
rect 128504 74916 128510 74928
rect 131482 74916 131488 74928
rect 128504 74888 131488 74916
rect 128504 74876 128510 74888
rect 131482 74876 131488 74888
rect 131540 74876 131546 74928
rect 135530 74876 135536 74928
rect 135588 74916 135594 74928
rect 135898 74916 135904 74928
rect 135588 74888 135904 74916
rect 135588 74876 135594 74888
rect 135898 74876 135904 74888
rect 135956 74876 135962 74928
rect 138106 74876 138112 74928
rect 138164 74916 138170 74928
rect 138750 74916 138756 74928
rect 138164 74888 138756 74916
rect 138164 74876 138170 74888
rect 138750 74876 138756 74888
rect 138808 74876 138814 74928
rect 139854 74876 139860 74928
rect 139912 74916 139918 74928
rect 140038 74916 140044 74928
rect 139912 74888 140044 74916
rect 139912 74876 139918 74888
rect 140038 74876 140044 74888
rect 140096 74876 140102 74928
rect 144914 74876 144920 74928
rect 144972 74916 144978 74928
rect 145466 74916 145472 74928
rect 144972 74888 145472 74916
rect 144972 74876 144978 74888
rect 145466 74876 145472 74888
rect 145524 74876 145530 74928
rect 147858 74876 147864 74928
rect 147916 74916 147922 74928
rect 148134 74916 148140 74928
rect 147916 74888 148140 74916
rect 147916 74876 147922 74888
rect 148134 74876 148140 74888
rect 148192 74876 148198 74928
rect 160094 74916 160100 74928
rect 150406 74888 160100 74916
rect 125134 74808 125140 74860
rect 125192 74848 125198 74860
rect 132310 74848 132316 74860
rect 125192 74820 132316 74848
rect 125192 74808 125198 74820
rect 132310 74808 132316 74820
rect 132368 74808 132374 74860
rect 134058 74808 134064 74860
rect 134116 74848 134122 74860
rect 134518 74848 134524 74860
rect 134116 74820 134524 74848
rect 134116 74808 134122 74820
rect 134518 74808 134524 74820
rect 134576 74808 134582 74860
rect 135438 74808 135444 74860
rect 135496 74848 135502 74860
rect 136174 74848 136180 74860
rect 135496 74820 136180 74848
rect 135496 74808 135502 74820
rect 136174 74808 136180 74820
rect 136232 74808 136238 74860
rect 136634 74808 136640 74860
rect 136692 74848 136698 74860
rect 137002 74848 137008 74860
rect 136692 74820 137008 74848
rect 136692 74808 136698 74820
rect 137002 74808 137008 74820
rect 137060 74808 137066 74860
rect 140774 74808 140780 74860
rect 140832 74848 140838 74860
rect 141418 74848 141424 74860
rect 140832 74820 141424 74848
rect 140832 74808 140838 74820
rect 141418 74808 141424 74820
rect 141476 74808 141482 74860
rect 145282 74808 145288 74860
rect 145340 74848 145346 74860
rect 145742 74848 145748 74860
rect 145340 74820 145748 74848
rect 145340 74808 145346 74820
rect 145742 74808 145748 74820
rect 145800 74808 145806 74860
rect 129734 74740 129740 74792
rect 129792 74780 129798 74792
rect 135622 74780 135628 74792
rect 129792 74752 135628 74780
rect 129792 74740 129798 74752
rect 135622 74740 135628 74752
rect 135680 74740 135686 74792
rect 135898 74740 135904 74792
rect 135956 74780 135962 74792
rect 136450 74780 136456 74792
rect 135956 74752 136456 74780
rect 135956 74740 135962 74752
rect 136450 74740 136456 74752
rect 136508 74740 136514 74792
rect 145466 74740 145472 74792
rect 145524 74780 145530 74792
rect 146018 74780 146024 74792
rect 145524 74752 146024 74780
rect 145524 74740 145530 74752
rect 146018 74740 146024 74752
rect 146076 74740 146082 74792
rect 150406 74780 150434 74888
rect 160094 74876 160100 74888
rect 160152 74876 160158 74928
rect 160554 74876 160560 74928
rect 160612 74916 160618 74928
rect 161382 74916 161388 74928
rect 160612 74888 161388 74916
rect 160612 74876 160618 74888
rect 161382 74876 161388 74888
rect 161440 74876 161446 74928
rect 167546 74876 167552 74928
rect 167604 74916 167610 74928
rect 167822 74916 167828 74928
rect 167604 74888 167828 74916
rect 167604 74876 167610 74888
rect 167822 74876 167828 74888
rect 167880 74876 167886 74928
rect 170122 74876 170128 74928
rect 170180 74916 170186 74928
rect 170950 74916 170956 74928
rect 170180 74888 170956 74916
rect 170180 74876 170186 74888
rect 170950 74876 170956 74888
rect 171008 74876 171014 74928
rect 171778 74876 171784 74928
rect 171836 74916 171842 74928
rect 183002 74916 183008 74928
rect 171836 74888 183008 74916
rect 171836 74876 171842 74888
rect 183002 74876 183008 74888
rect 183060 74876 183066 74928
rect 155218 74808 155224 74860
rect 155276 74848 155282 74860
rect 162118 74848 162124 74860
rect 155276 74820 162124 74848
rect 155276 74808 155282 74820
rect 162118 74808 162124 74820
rect 162176 74808 162182 74860
rect 162854 74808 162860 74860
rect 162912 74848 162918 74860
rect 163498 74848 163504 74860
rect 162912 74820 163504 74848
rect 162912 74808 162918 74820
rect 163498 74808 163504 74820
rect 163556 74808 163562 74860
rect 164418 74808 164424 74860
rect 164476 74848 164482 74860
rect 172238 74848 172244 74860
rect 164476 74820 172244 74848
rect 164476 74808 164482 74820
rect 172238 74808 172244 74820
rect 172296 74808 172302 74860
rect 149026 74752 150434 74780
rect 120718 74672 120724 74724
rect 120776 74712 120782 74724
rect 128630 74712 128636 74724
rect 120776 74684 128636 74712
rect 120776 74672 120782 74684
rect 128630 74672 128636 74684
rect 128688 74672 128694 74724
rect 135254 74672 135260 74724
rect 135312 74712 135318 74724
rect 136266 74712 136272 74724
rect 135312 74684 136272 74712
rect 135312 74672 135318 74684
rect 136266 74672 136272 74684
rect 136324 74672 136330 74724
rect 140866 74672 140872 74724
rect 140924 74712 140930 74724
rect 149026 74712 149054 74752
rect 158806 74740 158812 74792
rect 158864 74780 158870 74792
rect 159542 74780 159548 74792
rect 158864 74752 159548 74780
rect 158864 74740 158870 74752
rect 159542 74740 159548 74752
rect 159600 74740 159606 74792
rect 160370 74740 160376 74792
rect 160428 74780 160434 74792
rect 161014 74780 161020 74792
rect 160428 74752 161020 74780
rect 160428 74740 160434 74752
rect 161014 74740 161020 74752
rect 161072 74740 161078 74792
rect 165246 74740 165252 74792
rect 165304 74780 165310 74792
rect 170490 74780 170496 74792
rect 165304 74752 170496 74780
rect 165304 74740 165310 74752
rect 170490 74740 170496 74752
rect 170548 74740 170554 74792
rect 171870 74740 171876 74792
rect 171928 74780 171934 74792
rect 580718 74780 580724 74792
rect 171928 74752 580724 74780
rect 171928 74740 171934 74752
rect 580718 74740 580724 74752
rect 580776 74740 580782 74792
rect 140924 74684 149054 74712
rect 140924 74672 140930 74684
rect 154574 74672 154580 74724
rect 154632 74712 154638 74724
rect 155218 74712 155224 74724
rect 154632 74684 155224 74712
rect 154632 74672 154638 74684
rect 155218 74672 155224 74684
rect 155276 74672 155282 74724
rect 164418 74672 164424 74724
rect 164476 74712 164482 74724
rect 165154 74712 165160 74724
rect 164476 74684 165160 74712
rect 164476 74672 164482 74684
rect 165154 74672 165160 74684
rect 165212 74672 165218 74724
rect 165798 74672 165804 74724
rect 165856 74712 165862 74724
rect 166258 74712 166264 74724
rect 165856 74684 166264 74712
rect 165856 74672 165862 74684
rect 166258 74672 166264 74684
rect 166316 74672 166322 74724
rect 170398 74672 170404 74724
rect 170456 74712 170462 74724
rect 215938 74712 215944 74724
rect 170456 74684 215944 74712
rect 170456 74672 170462 74684
rect 215938 74672 215944 74684
rect 215996 74672 216002 74724
rect 134794 74644 134800 74656
rect 127360 74616 134800 74644
rect 124950 74468 124956 74520
rect 125008 74508 125014 74520
rect 127360 74508 127388 74616
rect 134794 74604 134800 74616
rect 134852 74604 134858 74656
rect 135622 74604 135628 74656
rect 135680 74644 135686 74656
rect 136358 74644 136364 74656
rect 135680 74616 136364 74644
rect 135680 74604 135686 74616
rect 136358 74604 136364 74616
rect 136416 74604 136422 74656
rect 162854 74604 162860 74656
rect 162912 74644 162918 74656
rect 163682 74644 163688 74656
rect 162912 74616 163688 74644
rect 162912 74604 162918 74616
rect 163682 74604 163688 74616
rect 163740 74604 163746 74656
rect 165614 74604 165620 74656
rect 165672 74644 165678 74656
rect 171502 74644 171508 74656
rect 165672 74616 171508 74644
rect 165672 74604 165678 74616
rect 171502 74604 171508 74616
rect 171560 74604 171566 74656
rect 131206 74536 131212 74588
rect 131264 74576 131270 74588
rect 131850 74576 131856 74588
rect 131264 74548 131856 74576
rect 131264 74536 131270 74548
rect 131850 74536 131856 74548
rect 131908 74536 131914 74588
rect 168558 74536 168564 74588
rect 168616 74576 168622 74588
rect 170766 74576 170772 74588
rect 168616 74548 170772 74576
rect 168616 74536 168622 74548
rect 170766 74536 170772 74548
rect 170824 74536 170830 74588
rect 171134 74508 171140 74520
rect 125008 74480 127388 74508
rect 127636 74480 171140 74508
rect 125008 74468 125014 74480
rect 122834 74400 122840 74452
rect 122892 74440 122898 74452
rect 126790 74440 126796 74452
rect 122892 74412 126796 74440
rect 122892 74400 122898 74412
rect 126790 74400 126796 74412
rect 126848 74400 126854 74452
rect 127636 74372 127664 74480
rect 171134 74468 171140 74480
rect 171192 74468 171198 74520
rect 130286 74400 130292 74452
rect 130344 74440 130350 74452
rect 131022 74440 131028 74452
rect 130344 74412 131028 74440
rect 130344 74400 130350 74412
rect 131022 74400 131028 74412
rect 131080 74400 131086 74452
rect 131114 74400 131120 74452
rect 131172 74440 131178 74452
rect 166994 74440 167000 74452
rect 131172 74412 167000 74440
rect 131172 74400 131178 74412
rect 166994 74400 167000 74412
rect 167052 74400 167058 74452
rect 168282 74440 168288 74452
rect 167104 74412 168288 74440
rect 127452 74344 127664 74372
rect 120994 74196 121000 74248
rect 121052 74236 121058 74248
rect 127452 74236 127480 74344
rect 128078 74332 128084 74384
rect 128136 74372 128142 74384
rect 167104 74372 167132 74412
rect 168282 74400 168288 74412
rect 168340 74400 168346 74452
rect 169386 74400 169392 74452
rect 169444 74440 169450 74452
rect 172974 74440 172980 74452
rect 169444 74412 172980 74440
rect 169444 74400 169450 74412
rect 172974 74400 172980 74412
rect 173032 74400 173038 74452
rect 128136 74344 167132 74372
rect 128136 74332 128142 74344
rect 168558 74332 168564 74384
rect 168616 74372 168622 74384
rect 168926 74372 168932 74384
rect 168616 74344 168932 74372
rect 168616 74332 168622 74344
rect 168926 74332 168932 74344
rect 168984 74332 168990 74384
rect 169754 74332 169760 74384
rect 169812 74372 169818 74384
rect 170398 74372 170404 74384
rect 169812 74344 170404 74372
rect 169812 74332 169818 74344
rect 170398 74332 170404 74344
rect 170456 74332 170462 74384
rect 128464 74276 132356 74304
rect 128464 74236 128492 74276
rect 121052 74208 127480 74236
rect 128234 74208 128492 74236
rect 121052 74196 121058 74208
rect 102134 74128 102140 74180
rect 102192 74168 102198 74180
rect 128234 74168 128262 74208
rect 131850 74196 131856 74248
rect 131908 74236 131914 74248
rect 132218 74236 132224 74248
rect 131908 74208 132224 74236
rect 131908 74196 131914 74208
rect 132218 74196 132224 74208
rect 132276 74196 132282 74248
rect 131942 74168 131948 74180
rect 102192 74140 128262 74168
rect 128740 74140 131948 74168
rect 102192 74128 102198 74140
rect 93854 74060 93860 74112
rect 93912 74100 93918 74112
rect 128630 74100 128636 74112
rect 93912 74072 128636 74100
rect 93912 74060 93918 74072
rect 128630 74060 128636 74072
rect 128688 74060 128694 74112
rect 86954 73992 86960 74044
rect 87012 74032 87018 74044
rect 128740 74032 128768 74140
rect 131942 74128 131948 74140
rect 132000 74128 132006 74180
rect 132328 74168 132356 74276
rect 133046 74264 133052 74316
rect 133104 74304 133110 74316
rect 133782 74304 133788 74316
rect 133104 74276 133788 74304
rect 133104 74264 133110 74276
rect 133782 74264 133788 74276
rect 133840 74264 133846 74316
rect 137094 74264 137100 74316
rect 137152 74304 137158 74316
rect 137462 74304 137468 74316
rect 137152 74276 137468 74304
rect 137152 74264 137158 74276
rect 137462 74264 137468 74276
rect 137520 74264 137526 74316
rect 143810 74264 143816 74316
rect 143868 74304 143874 74316
rect 144454 74304 144460 74316
rect 143868 74276 144460 74304
rect 143868 74264 143874 74276
rect 144454 74264 144460 74276
rect 144512 74264 144518 74316
rect 147674 74264 147680 74316
rect 147732 74304 147738 74316
rect 148410 74304 148416 74316
rect 147732 74276 148416 74304
rect 147732 74264 147738 74276
rect 148410 74264 148416 74276
rect 148468 74264 148474 74316
rect 153102 74264 153108 74316
rect 153160 74304 153166 74316
rect 197354 74304 197360 74316
rect 153160 74276 197360 74304
rect 153160 74264 153166 74276
rect 197354 74264 197360 74276
rect 197412 74264 197418 74316
rect 132770 74196 132776 74248
rect 132828 74236 132834 74248
rect 133690 74236 133696 74248
rect 132828 74208 133696 74236
rect 132828 74196 132834 74208
rect 133690 74196 133696 74208
rect 133748 74196 133754 74248
rect 133966 74196 133972 74248
rect 134024 74236 134030 74248
rect 134426 74236 134432 74248
rect 134024 74208 134432 74236
rect 134024 74196 134030 74208
rect 134426 74196 134432 74208
rect 134484 74196 134490 74248
rect 134610 74196 134616 74248
rect 134668 74236 134674 74248
rect 135162 74236 135168 74248
rect 134668 74208 135168 74236
rect 134668 74196 134674 74208
rect 135162 74196 135168 74208
rect 135220 74196 135226 74248
rect 142246 74196 142252 74248
rect 142304 74236 142310 74248
rect 142706 74236 142712 74248
rect 142304 74208 142712 74236
rect 142304 74196 142310 74208
rect 142706 74196 142712 74208
rect 142764 74196 142770 74248
rect 147490 74196 147496 74248
rect 147548 74236 147554 74248
rect 226334 74236 226340 74248
rect 147548 74208 226340 74236
rect 147548 74196 147554 74208
rect 226334 74196 226340 74208
rect 226392 74196 226398 74248
rect 133414 74168 133420 74180
rect 132328 74140 133420 74168
rect 133414 74128 133420 74140
rect 133472 74128 133478 74180
rect 139946 74128 139952 74180
rect 140004 74168 140010 74180
rect 140314 74168 140320 74180
rect 140004 74140 140320 74168
rect 140004 74128 140010 74140
rect 140314 74128 140320 74140
rect 140372 74128 140378 74180
rect 144546 74128 144552 74180
rect 144604 74168 144610 74180
rect 240134 74168 240140 74180
rect 144604 74140 240140 74168
rect 144604 74128 144610 74140
rect 240134 74128 240140 74140
rect 240192 74128 240198 74180
rect 131390 74060 131396 74112
rect 131448 74100 131454 74112
rect 132402 74100 132408 74112
rect 131448 74072 132408 74100
rect 131448 74060 131454 74072
rect 132402 74060 132408 74072
rect 132460 74060 132466 74112
rect 132678 74060 132684 74112
rect 132736 74100 132742 74112
rect 133598 74100 133604 74112
rect 132736 74072 133604 74100
rect 132736 74060 132742 74072
rect 133598 74060 133604 74072
rect 133656 74060 133662 74112
rect 138290 74060 138296 74112
rect 138348 74100 138354 74112
rect 138658 74100 138664 74112
rect 138348 74072 138664 74100
rect 138348 74060 138354 74072
rect 138658 74060 138664 74072
rect 138716 74060 138722 74112
rect 142338 74060 142344 74112
rect 142396 74100 142402 74112
rect 142706 74100 142712 74112
rect 142396 74072 142712 74100
rect 142396 74060 142402 74072
rect 142706 74060 142712 74072
rect 142764 74060 142770 74112
rect 145926 74060 145932 74112
rect 145984 74100 145990 74112
rect 260834 74100 260840 74112
rect 145984 74072 260840 74100
rect 145984 74060 145990 74072
rect 260834 74060 260840 74072
rect 260892 74060 260898 74112
rect 87012 74004 128768 74032
rect 87012 73992 87018 74004
rect 131482 73992 131488 74044
rect 131540 74032 131546 74044
rect 132126 74032 132132 74044
rect 131540 74004 132132 74032
rect 131540 73992 131546 74004
rect 132126 73992 132132 74004
rect 132184 73992 132190 74044
rect 138566 73992 138572 74044
rect 138624 74032 138630 74044
rect 138842 74032 138848 74044
rect 138624 74004 138848 74032
rect 138624 73992 138630 74004
rect 138842 73992 138848 74004
rect 138900 73992 138906 74044
rect 139394 73992 139400 74044
rect 139452 74032 139458 74044
rect 140222 74032 140228 74044
rect 139452 74004 140228 74032
rect 139452 73992 139458 74004
rect 140222 73992 140228 74004
rect 140280 73992 140286 74044
rect 160186 73992 160192 74044
rect 160244 74032 160250 74044
rect 160830 74032 160836 74044
rect 160244 74004 160836 74032
rect 160244 73992 160250 74004
rect 160830 73992 160836 74004
rect 160888 73992 160894 74044
rect 296714 74032 296720 74044
rect 166184 74004 296720 74032
rect 69014 73924 69020 73976
rect 69072 73964 69078 73976
rect 124766 73964 124772 73976
rect 69072 73936 124772 73964
rect 69072 73924 69078 73936
rect 124766 73924 124772 73936
rect 124824 73924 124830 73976
rect 134518 73924 134524 73976
rect 134576 73964 134582 73976
rect 135346 73964 135352 73976
rect 134576 73936 135352 73964
rect 134576 73924 134582 73936
rect 135346 73924 135352 73936
rect 135404 73924 135410 73976
rect 136818 73924 136824 73976
rect 136876 73964 136882 73976
rect 137830 73964 137836 73976
rect 136876 73936 137836 73964
rect 136876 73924 136882 73936
rect 137830 73924 137836 73936
rect 137888 73924 137894 73976
rect 146386 73924 146392 73976
rect 146444 73964 146450 73976
rect 146662 73964 146668 73976
rect 146444 73936 146668 73964
rect 146444 73924 146450 73936
rect 146662 73924 146668 73936
rect 146720 73924 146726 73976
rect 44174 73856 44180 73908
rect 44232 73896 44238 73908
rect 44232 73868 120120 73896
rect 44232 73856 44238 73868
rect 30374 73788 30380 73840
rect 30432 73828 30438 73840
rect 120092 73828 120120 73868
rect 122190 73856 122196 73908
rect 122248 73896 122254 73908
rect 127526 73896 127532 73908
rect 122248 73868 127532 73896
rect 122248 73856 122254 73868
rect 127526 73856 127532 73868
rect 127584 73856 127590 73908
rect 143074 73856 143080 73908
rect 143132 73896 143138 73908
rect 147490 73896 147496 73908
rect 143132 73868 147496 73896
rect 143132 73856 143138 73868
rect 147490 73856 147496 73868
rect 147548 73856 147554 73908
rect 159082 73856 159088 73908
rect 159140 73896 159146 73908
rect 159266 73896 159272 73908
rect 159140 73868 159272 73896
rect 159140 73856 159146 73868
rect 159266 73856 159272 73868
rect 159324 73856 159330 73908
rect 128354 73828 128360 73840
rect 30432 73800 118694 73828
rect 120092 73800 128360 73828
rect 30432 73788 30438 73800
rect 118666 73760 118694 73800
rect 128354 73788 128360 73800
rect 128412 73788 128418 73840
rect 127986 73760 127992 73772
rect 118666 73732 127992 73760
rect 127986 73720 127992 73732
rect 128044 73720 128050 73772
rect 143718 73720 143724 73772
rect 143776 73760 143782 73772
rect 144362 73760 144368 73772
rect 143776 73732 144368 73760
rect 143776 73720 143782 73732
rect 144362 73720 144368 73732
rect 144420 73720 144426 73772
rect 151906 73720 151912 73772
rect 151964 73760 151970 73772
rect 152642 73760 152648 73772
rect 151964 73732 152648 73760
rect 151964 73720 151970 73732
rect 152642 73720 152648 73732
rect 152700 73720 152706 73772
rect 155586 73720 155592 73772
rect 155644 73760 155650 73772
rect 166184 73760 166212 74004
rect 296714 73992 296720 74004
rect 296772 73992 296778 74044
rect 382274 73964 382280 73976
rect 155644 73732 166212 73760
rect 166644 73936 382280 73964
rect 155644 73720 155650 73732
rect 120902 73652 120908 73704
rect 120960 73692 120966 73704
rect 127066 73692 127072 73704
rect 120960 73664 127072 73692
rect 120960 73652 120966 73664
rect 127066 73652 127072 73664
rect 127124 73652 127130 73704
rect 136726 73652 136732 73704
rect 136784 73692 136790 73704
rect 138934 73692 138940 73704
rect 136784 73664 138940 73692
rect 136784 73652 136790 73664
rect 138934 73652 138940 73664
rect 138992 73652 138998 73704
rect 161934 73652 161940 73704
rect 161992 73692 161998 73704
rect 162302 73692 162308 73704
rect 161992 73664 162308 73692
rect 161992 73652 161998 73664
rect 162302 73652 162308 73664
rect 162360 73652 162366 73704
rect 165706 73652 165712 73704
rect 165764 73692 165770 73704
rect 166258 73692 166264 73704
rect 165764 73664 166264 73692
rect 165764 73652 165770 73664
rect 166258 73652 166264 73664
rect 166316 73652 166322 73704
rect 120810 73584 120816 73636
rect 120868 73624 120874 73636
rect 128078 73624 128084 73636
rect 120868 73596 128084 73624
rect 120868 73584 120874 73596
rect 128078 73584 128084 73596
rect 128136 73584 128142 73636
rect 157242 73584 157248 73636
rect 157300 73624 157306 73636
rect 166644 73624 166672 73936
rect 382274 73924 382280 73936
rect 382332 73924 382338 73976
rect 166902 73856 166908 73908
rect 166960 73896 166966 73908
rect 390554 73896 390560 73908
rect 166960 73868 390560 73896
rect 166960 73856 166966 73868
rect 390554 73856 390560 73868
rect 390612 73856 390618 73908
rect 168374 73788 168380 73840
rect 168432 73828 168438 73840
rect 168926 73828 168932 73840
rect 168432 73800 168932 73828
rect 168432 73788 168438 73800
rect 168926 73788 168932 73800
rect 168984 73788 168990 73840
rect 169754 73788 169760 73840
rect 169812 73828 169818 73840
rect 170674 73828 170680 73840
rect 169812 73800 170680 73828
rect 169812 73788 169818 73800
rect 170674 73788 170680 73800
rect 170732 73788 170738 73840
rect 558914 73828 558920 73840
rect 176626 73800 558920 73828
rect 166718 73720 166724 73772
rect 166776 73760 166782 73772
rect 171870 73760 171876 73772
rect 166776 73732 171876 73760
rect 166776 73720 166782 73732
rect 171870 73720 171876 73732
rect 171928 73720 171934 73772
rect 169662 73652 169668 73704
rect 169720 73692 169726 73704
rect 176626 73692 176654 73800
rect 558914 73788 558920 73800
rect 558972 73788 558978 73840
rect 169720 73664 176654 73692
rect 169720 73652 169726 73664
rect 157300 73596 166672 73624
rect 157300 73584 157306 73596
rect 168282 73584 168288 73636
rect 168340 73624 168346 73636
rect 172698 73624 172704 73636
rect 168340 73596 172704 73624
rect 168340 73584 168346 73596
rect 172698 73584 172704 73596
rect 172756 73584 172762 73636
rect 125870 73516 125876 73568
rect 125928 73556 125934 73568
rect 126330 73556 126336 73568
rect 125928 73528 126336 73556
rect 125928 73516 125934 73528
rect 126330 73516 126336 73528
rect 126388 73516 126394 73568
rect 127066 73516 127072 73568
rect 127124 73556 127130 73568
rect 131114 73556 131120 73568
rect 127124 73528 131120 73556
rect 127124 73516 127130 73528
rect 131114 73516 131120 73528
rect 131172 73516 131178 73568
rect 165614 73516 165620 73568
rect 165672 73556 165678 73568
rect 166626 73556 166632 73568
rect 165672 73528 166632 73556
rect 165672 73516 165678 73528
rect 166626 73516 166632 73528
rect 166684 73516 166690 73568
rect 136726 73448 136732 73500
rect 136784 73488 136790 73500
rect 137278 73488 137284 73500
rect 136784 73460 137284 73488
rect 136784 73448 136790 73460
rect 137278 73448 137284 73460
rect 137336 73448 137342 73500
rect 139578 73448 139584 73500
rect 139636 73488 139642 73500
rect 140130 73488 140136 73500
rect 139636 73460 140136 73488
rect 139636 73448 139642 73460
rect 140130 73448 140136 73460
rect 140188 73448 140194 73500
rect 152826 73448 152832 73500
rect 152884 73488 152890 73500
rect 161014 73488 161020 73500
rect 152884 73460 161020 73488
rect 152884 73448 152890 73460
rect 161014 73448 161020 73460
rect 161072 73448 161078 73500
rect 161290 73448 161296 73500
rect 161348 73488 161354 73500
rect 172422 73488 172428 73500
rect 161348 73460 172428 73488
rect 161348 73448 161354 73460
rect 172422 73448 172428 73460
rect 172480 73448 172486 73500
rect 146570 73380 146576 73432
rect 146628 73420 146634 73432
rect 147214 73420 147220 73432
rect 146628 73392 147220 73420
rect 146628 73380 146634 73392
rect 147214 73380 147220 73392
rect 147272 73380 147278 73432
rect 149238 73380 149244 73432
rect 149296 73420 149302 73432
rect 152642 73420 152648 73432
rect 149296 73392 152648 73420
rect 149296 73380 149302 73392
rect 152642 73380 152648 73392
rect 152700 73380 152706 73432
rect 166166 73380 166172 73432
rect 166224 73420 166230 73432
rect 166810 73420 166816 73432
rect 166224 73392 166816 73420
rect 166224 73380 166230 73392
rect 166810 73380 166816 73392
rect 166868 73380 166874 73432
rect 127526 73312 127532 73364
rect 127584 73352 127590 73364
rect 127894 73352 127900 73364
rect 127584 73324 127900 73352
rect 127584 73312 127590 73324
rect 127894 73312 127900 73324
rect 127952 73312 127958 73364
rect 152182 73312 152188 73364
rect 152240 73352 152246 73364
rect 152550 73352 152556 73364
rect 152240 73324 152556 73352
rect 152240 73312 152246 73324
rect 152550 73312 152556 73324
rect 152608 73312 152614 73364
rect 163038 73312 163044 73364
rect 163096 73352 163102 73364
rect 163774 73352 163780 73364
rect 163096 73324 163780 73352
rect 163096 73312 163102 73324
rect 163774 73312 163780 73324
rect 163832 73312 163838 73364
rect 137370 73244 137376 73296
rect 137428 73284 137434 73296
rect 144454 73284 144460 73296
rect 137428 73256 144460 73284
rect 137428 73244 137434 73256
rect 144454 73244 144460 73256
rect 144512 73244 144518 73296
rect 149238 73244 149244 73296
rect 149296 73284 149302 73296
rect 150066 73284 150072 73296
rect 149296 73256 150072 73284
rect 149296 73244 149302 73256
rect 150066 73244 150072 73256
rect 150124 73244 150130 73296
rect 132586 73176 132592 73228
rect 132644 73216 132650 73228
rect 132954 73216 132960 73228
rect 132644 73188 132960 73216
rect 132644 73176 132650 73188
rect 132954 73176 132960 73188
rect 133012 73176 133018 73228
rect 128354 73108 128360 73160
rect 128412 73148 128418 73160
rect 133506 73148 133512 73160
rect 128412 73120 133512 73148
rect 128412 73108 128418 73120
rect 133506 73108 133512 73120
rect 133564 73108 133570 73160
rect 431954 73108 431960 73160
rect 432012 73148 432018 73160
rect 580166 73148 580172 73160
rect 432012 73120 580172 73148
rect 432012 73108 432018 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 140958 73040 140964 73092
rect 141016 73080 141022 73092
rect 141510 73080 141516 73092
rect 141016 73052 141516 73080
rect 141016 73040 141022 73052
rect 141510 73040 141516 73052
rect 141568 73040 141574 73092
rect 132954 72972 132960 73024
rect 133012 73012 133018 73024
rect 133322 73012 133328 73024
rect 133012 72984 133328 73012
rect 133012 72972 133018 72984
rect 133322 72972 133328 72984
rect 133380 72972 133386 73024
rect 121454 72836 121460 72888
rect 121512 72876 121518 72888
rect 134978 72876 134984 72888
rect 121512 72848 134984 72876
rect 121512 72836 121518 72848
rect 134978 72836 134984 72848
rect 135036 72836 135042 72888
rect 107654 72768 107660 72820
rect 107712 72808 107718 72820
rect 129366 72808 129372 72820
rect 107712 72780 129372 72808
rect 107712 72768 107718 72780
rect 129366 72768 129372 72780
rect 129424 72768 129430 72820
rect 162670 72768 162676 72820
rect 162728 72808 162734 72820
rect 172054 72808 172060 72820
rect 162728 72780 172060 72808
rect 162728 72768 162734 72780
rect 172054 72768 172060 72780
rect 172112 72768 172118 72820
rect 51074 72700 51080 72752
rect 51132 72740 51138 72752
rect 129458 72740 129464 72752
rect 51132 72712 129464 72740
rect 51132 72700 51138 72712
rect 129458 72700 129464 72712
rect 129516 72700 129522 72752
rect 159910 72700 159916 72752
rect 159968 72740 159974 72752
rect 431954 72740 431960 72752
rect 159968 72712 431960 72740
rect 159968 72700 159974 72712
rect 431954 72700 431960 72712
rect 432012 72700 432018 72752
rect 60734 72632 60740 72684
rect 60792 72672 60798 72684
rect 130746 72672 130752 72684
rect 60792 72644 130752 72672
rect 60792 72632 60798 72644
rect 130746 72632 130752 72644
rect 130804 72632 130810 72684
rect 152918 72632 152924 72684
rect 152976 72672 152982 72684
rect 158346 72672 158352 72684
rect 152976 72644 158352 72672
rect 152976 72632 152982 72644
rect 158346 72632 158352 72644
rect 158404 72632 158410 72684
rect 163866 72632 163872 72684
rect 163924 72672 163930 72684
rect 438854 72672 438860 72684
rect 163924 72644 438860 72672
rect 163924 72632 163930 72644
rect 438854 72632 438860 72644
rect 438912 72632 438918 72684
rect 42794 72564 42800 72616
rect 42852 72604 42858 72616
rect 128906 72604 128912 72616
rect 42852 72576 128912 72604
rect 42852 72564 42858 72576
rect 128906 72564 128912 72576
rect 128964 72564 128970 72616
rect 150710 72564 150716 72616
rect 150768 72604 150774 72616
rect 151262 72604 151268 72616
rect 150768 72576 151268 72604
rect 150768 72564 150774 72576
rect 151262 72564 151268 72576
rect 151320 72564 151326 72616
rect 161198 72564 161204 72616
rect 161256 72604 161262 72616
rect 454034 72604 454040 72616
rect 161256 72576 454040 72604
rect 161256 72564 161262 72576
rect 454034 72564 454040 72576
rect 454092 72564 454098 72616
rect 16574 72496 16580 72548
rect 16632 72536 16638 72548
rect 16632 72508 123432 72536
rect 16632 72496 16638 72508
rect 6914 72428 6920 72480
rect 6972 72468 6978 72480
rect 121638 72468 121644 72480
rect 6972 72440 121644 72468
rect 6972 72428 6978 72440
rect 121638 72428 121644 72440
rect 121696 72428 121702 72480
rect 123404 72468 123432 72508
rect 126330 72496 126336 72548
rect 126388 72536 126394 72548
rect 126606 72536 126612 72548
rect 126388 72508 126612 72536
rect 126388 72496 126394 72508
rect 126606 72496 126612 72508
rect 126664 72496 126670 72548
rect 154942 72496 154948 72548
rect 155000 72536 155006 72548
rect 155494 72536 155500 72548
rect 155000 72508 155500 72536
rect 155000 72496 155006 72508
rect 155494 72496 155500 72508
rect 155552 72496 155558 72548
rect 164050 72496 164056 72548
rect 164108 72536 164114 72548
rect 489914 72536 489920 72548
rect 164108 72508 489920 72536
rect 164108 72496 164114 72508
rect 489914 72496 489920 72508
rect 489972 72496 489978 72548
rect 126882 72468 126888 72480
rect 123404 72440 126888 72468
rect 126882 72428 126888 72440
rect 126940 72428 126946 72480
rect 128630 72428 128636 72480
rect 128688 72468 128694 72480
rect 129642 72468 129648 72480
rect 128688 72440 129648 72468
rect 128688 72428 128694 72440
rect 129642 72428 129648 72440
rect 129700 72428 129706 72480
rect 138750 72428 138756 72480
rect 138808 72468 138814 72480
rect 138808 72440 157334 72468
rect 138808 72428 138814 72440
rect 124214 72360 124220 72412
rect 124272 72400 124278 72412
rect 125410 72400 125416 72412
rect 124272 72372 125416 72400
rect 124272 72360 124278 72372
rect 125410 72360 125416 72372
rect 125468 72360 125474 72412
rect 157306 72332 157334 72440
rect 167822 72428 167828 72480
rect 167880 72468 167886 72480
rect 535454 72468 535460 72480
rect 167880 72440 535460 72468
rect 167880 72428 167886 72440
rect 535454 72428 535460 72440
rect 535512 72428 535518 72480
rect 168650 72360 168656 72412
rect 168708 72400 168714 72412
rect 169110 72400 169116 72412
rect 168708 72372 169116 72400
rect 168708 72360 168714 72372
rect 169110 72360 169116 72372
rect 169168 72360 169174 72412
rect 174262 72360 174268 72412
rect 174320 72400 174326 72412
rect 174630 72400 174636 72412
rect 174320 72372 174636 72400
rect 174320 72360 174326 72372
rect 174630 72360 174636 72372
rect 174688 72360 174694 72412
rect 163774 72332 163780 72344
rect 157306 72304 163780 72332
rect 163774 72292 163780 72304
rect 163832 72292 163838 72344
rect 168374 72292 168380 72344
rect 168432 72332 168438 72344
rect 169202 72332 169208 72344
rect 168432 72304 169208 72332
rect 168432 72292 168438 72304
rect 169202 72292 169208 72304
rect 169260 72292 169266 72344
rect 168742 72224 168748 72276
rect 168800 72264 168806 72276
rect 169110 72264 169116 72276
rect 168800 72236 169116 72264
rect 168800 72224 168806 72236
rect 169110 72224 169116 72236
rect 169168 72224 169174 72276
rect 151446 72088 151452 72140
rect 151504 72128 151510 72140
rect 154206 72128 154212 72140
rect 151504 72100 154212 72128
rect 151504 72088 151510 72100
rect 154206 72088 154212 72100
rect 154264 72088 154270 72140
rect 168742 72088 168748 72140
rect 168800 72128 168806 72140
rect 169294 72128 169300 72140
rect 168800 72100 169300 72128
rect 168800 72088 168806 72100
rect 169294 72088 169300 72100
rect 169352 72088 169358 72140
rect 159082 71952 159088 72004
rect 159140 71992 159146 72004
rect 159450 71992 159456 72004
rect 159140 71964 159456 71992
rect 159140 71952 159146 71964
rect 159450 71952 159456 71964
rect 159508 71952 159514 72004
rect 154666 71816 154672 71868
rect 154724 71856 154730 71868
rect 155402 71856 155408 71868
rect 154724 71828 155408 71856
rect 154724 71816 154730 71828
rect 155402 71816 155408 71828
rect 155460 71816 155466 71868
rect 163958 71748 163964 71800
rect 164016 71788 164022 71800
rect 170674 71788 170680 71800
rect 164016 71760 170680 71788
rect 164016 71748 164022 71760
rect 170674 71748 170680 71760
rect 170732 71748 170738 71800
rect 3510 71680 3516 71732
rect 3568 71720 3574 71732
rect 171778 71720 171784 71732
rect 3568 71692 171784 71720
rect 3568 71680 3574 71692
rect 171778 71680 171784 71692
rect 171836 71680 171842 71732
rect 137646 71612 137652 71664
rect 137704 71652 137710 71664
rect 142982 71652 142988 71664
rect 137704 71624 142988 71652
rect 137704 71612 137710 71624
rect 142982 71612 142988 71624
rect 143040 71612 143046 71664
rect 149606 71544 149612 71596
rect 149664 71584 149670 71596
rect 150250 71584 150256 71596
rect 149664 71556 150256 71584
rect 149664 71544 149670 71556
rect 150250 71544 150256 71556
rect 150308 71544 150314 71596
rect 171042 71544 171048 71596
rect 171100 71584 171106 71596
rect 171778 71584 171784 71596
rect 171100 71556 171784 71584
rect 171100 71544 171106 71556
rect 171778 71544 171784 71556
rect 171836 71544 171842 71596
rect 140682 71408 140688 71460
rect 140740 71448 140746 71460
rect 184934 71448 184940 71460
rect 140740 71420 184940 71448
rect 140740 71408 140746 71420
rect 184934 71408 184940 71420
rect 184992 71408 184998 71460
rect 118694 71340 118700 71392
rect 118752 71380 118758 71392
rect 134058 71380 134064 71392
rect 118752 71352 134064 71380
rect 118752 71340 118758 71352
rect 134058 71340 134064 71352
rect 134116 71340 134122 71392
rect 154114 71340 154120 71392
rect 154172 71380 154178 71392
rect 211798 71380 211804 71392
rect 154172 71352 211804 71380
rect 154172 71340 154178 71352
rect 211798 71340 211804 71352
rect 211856 71340 211862 71392
rect 93946 71272 93952 71324
rect 94004 71312 94010 71324
rect 132586 71312 132592 71324
rect 94004 71284 132592 71312
rect 94004 71272 94010 71284
rect 132586 71272 132592 71284
rect 132644 71272 132650 71324
rect 141786 71272 141792 71324
rect 141844 71312 141850 71324
rect 209774 71312 209780 71324
rect 141844 71284 209780 71312
rect 141844 71272 141850 71284
rect 209774 71272 209780 71284
rect 209832 71272 209838 71324
rect 75914 71204 75920 71256
rect 75972 71244 75978 71256
rect 131206 71244 131212 71256
rect 75972 71216 131212 71244
rect 75972 71204 75978 71216
rect 131206 71204 131212 71216
rect 131264 71204 131270 71256
rect 142890 71204 142896 71256
rect 142948 71244 142954 71256
rect 216674 71244 216680 71256
rect 142948 71216 216680 71244
rect 142948 71204 142954 71216
rect 216674 71204 216680 71216
rect 216732 71204 216738 71256
rect 64874 71136 64880 71188
rect 64932 71176 64938 71188
rect 130838 71176 130844 71188
rect 64932 71148 130844 71176
rect 64932 71136 64938 71148
rect 130838 71136 130844 71148
rect 130896 71136 130902 71188
rect 143074 71136 143080 71188
rect 143132 71176 143138 71188
rect 223574 71176 223580 71188
rect 143132 71148 223580 71176
rect 143132 71136 143138 71148
rect 223574 71136 223580 71148
rect 223632 71136 223638 71188
rect 46934 71068 46940 71120
rect 46992 71108 46998 71120
rect 127618 71108 127624 71120
rect 46992 71080 127624 71108
rect 46992 71068 46998 71080
rect 127618 71068 127624 71080
rect 127676 71068 127682 71120
rect 147858 71068 147864 71120
rect 147916 71108 147922 71120
rect 148226 71108 148232 71120
rect 147916 71080 148232 71108
rect 147916 71068 147922 71080
rect 148226 71068 148232 71080
rect 148284 71068 148290 71120
rect 161382 71068 161388 71120
rect 161440 71108 161446 71120
rect 375374 71108 375380 71120
rect 161440 71080 375380 71108
rect 161440 71068 161446 71080
rect 375374 71068 375380 71080
rect 375432 71068 375438 71120
rect 26234 71000 26240 71052
rect 26292 71040 26298 71052
rect 126606 71040 126612 71052
rect 26292 71012 126612 71040
rect 26292 71000 26298 71012
rect 126606 71000 126612 71012
rect 126664 71000 126670 71052
rect 169110 71000 169116 71052
rect 169168 71040 169174 71052
rect 564434 71040 564440 71052
rect 169168 71012 564440 71040
rect 169168 71000 169174 71012
rect 564434 71000 564440 71012
rect 564492 71000 564498 71052
rect 141142 70864 141148 70916
rect 141200 70904 141206 70916
rect 141694 70904 141700 70916
rect 141200 70876 141700 70904
rect 141200 70864 141206 70876
rect 141694 70864 141700 70876
rect 141752 70864 141758 70916
rect 142338 70864 142344 70916
rect 142396 70904 142402 70916
rect 142798 70904 142804 70916
rect 142396 70876 142804 70904
rect 142396 70864 142402 70876
rect 142798 70864 142804 70876
rect 142856 70864 142862 70916
rect 146846 70728 146852 70780
rect 146904 70768 146910 70780
rect 147122 70768 147128 70780
rect 146904 70740 147128 70768
rect 146904 70728 146910 70740
rect 147122 70728 147128 70740
rect 147180 70728 147186 70780
rect 148226 70728 148232 70780
rect 148284 70768 148290 70780
rect 148502 70768 148508 70780
rect 148284 70740 148508 70768
rect 148284 70728 148290 70740
rect 148502 70728 148508 70740
rect 148560 70728 148566 70780
rect 150986 70456 150992 70508
rect 151044 70496 151050 70508
rect 151354 70496 151360 70508
rect 151044 70468 151360 70496
rect 151044 70456 151050 70468
rect 151354 70456 151360 70468
rect 151412 70456 151418 70508
rect 151814 70456 151820 70508
rect 151872 70496 151878 70508
rect 152458 70496 152464 70508
rect 151872 70468 152464 70496
rect 151872 70456 151878 70468
rect 152458 70456 152464 70468
rect 152516 70456 152522 70508
rect 152642 69980 152648 70032
rect 152700 70020 152706 70032
rect 304994 70020 305000 70032
rect 152700 69992 305000 70020
rect 152700 69980 152706 69992
rect 304994 69980 305000 69992
rect 305052 69980 305058 70032
rect 149882 69912 149888 69964
rect 149940 69952 149946 69964
rect 311894 69952 311900 69964
rect 149940 69924 311900 69952
rect 149940 69912 149946 69924
rect 311894 69912 311900 69924
rect 311952 69912 311958 69964
rect 151170 69844 151176 69896
rect 151228 69884 151234 69896
rect 325694 69884 325700 69896
rect 151228 69856 325700 69884
rect 151228 69844 151234 69856
rect 325694 69844 325700 69856
rect 325752 69844 325758 69896
rect 154482 69776 154488 69828
rect 154540 69816 154546 69828
rect 332594 69816 332600 69828
rect 154540 69788 332600 69816
rect 154540 69776 154546 69788
rect 332594 69776 332600 69788
rect 332652 69776 332658 69828
rect 154022 69708 154028 69760
rect 154080 69748 154086 69760
rect 340874 69748 340880 69760
rect 154080 69720 340880 69748
rect 154080 69708 154086 69720
rect 340874 69708 340880 69720
rect 340932 69708 340938 69760
rect 114554 69640 114560 69692
rect 114612 69680 114618 69692
rect 133966 69680 133972 69692
rect 114612 69652 133972 69680
rect 114612 69640 114618 69652
rect 133966 69640 133972 69652
rect 134024 69640 134030 69692
rect 138658 69640 138664 69692
rect 138716 69680 138722 69692
rect 149974 69680 149980 69692
rect 138716 69652 149980 69680
rect 138716 69640 138722 69652
rect 149974 69640 149980 69652
rect 150032 69640 150038 69692
rect 156782 69640 156788 69692
rect 156840 69680 156846 69692
rect 382366 69680 382372 69692
rect 156840 69652 382372 69680
rect 156840 69640 156846 69652
rect 382366 69640 382372 69652
rect 382424 69640 382430 69692
rect 149054 69572 149060 69624
rect 149112 69612 149118 69624
rect 149790 69612 149796 69624
rect 149112 69584 149796 69612
rect 149112 69572 149118 69584
rect 149790 69572 149796 69584
rect 149848 69572 149854 69624
rect 138566 68960 138572 69012
rect 138624 69000 138630 69012
rect 142798 69000 142804 69012
rect 138624 68972 142804 69000
rect 138624 68960 138630 68972
rect 142798 68960 142804 68972
rect 142856 68960 142862 69012
rect 148962 68552 148968 68604
rect 149020 68592 149026 68604
rect 190454 68592 190460 68604
rect 149020 68564 190460 68592
rect 149020 68552 149026 68564
rect 190454 68552 190460 68564
rect 190512 68552 190518 68604
rect 163590 68484 163596 68536
rect 163648 68524 163654 68536
rect 487154 68524 487160 68536
rect 163648 68496 487160 68524
rect 163648 68484 163654 68496
rect 487154 68484 487160 68496
rect 487212 68484 487218 68536
rect 165522 68416 165528 68468
rect 165580 68456 165586 68468
rect 500954 68456 500960 68468
rect 165580 68428 500960 68456
rect 165580 68416 165586 68428
rect 500954 68416 500960 68428
rect 501012 68416 501018 68468
rect 164970 68348 164976 68400
rect 165028 68388 165034 68400
rect 505094 68388 505100 68400
rect 165028 68360 505100 68388
rect 165028 68348 165034 68360
rect 505094 68348 505100 68360
rect 505152 68348 505158 68400
rect 169018 68280 169024 68332
rect 169076 68320 169082 68332
rect 564526 68320 564532 68332
rect 169076 68292 564532 68320
rect 169076 68280 169082 68292
rect 564526 68280 564532 68292
rect 564584 68280 564590 68332
rect 140038 67192 140044 67244
rect 140096 67232 140102 67244
rect 182174 67232 182180 67244
rect 140096 67204 182180 67232
rect 140096 67192 140102 67204
rect 182174 67192 182180 67204
rect 182232 67192 182238 67244
rect 141510 67124 141516 67176
rect 141568 67164 141574 67176
rect 209866 67164 209872 67176
rect 141568 67136 209872 67164
rect 141568 67124 141574 67136
rect 209866 67124 209872 67136
rect 209924 67124 209930 67176
rect 156690 67056 156696 67108
rect 156748 67096 156754 67108
rect 396074 67096 396080 67108
rect 156748 67068 396080 67096
rect 156748 67056 156754 67068
rect 396074 67056 396080 67068
rect 396132 67056 396138 67108
rect 166350 66988 166356 67040
rect 166408 67028 166414 67040
rect 523034 67028 523040 67040
rect 166408 67000 523040 67028
rect 166408 66988 166414 67000
rect 523034 66988 523040 67000
rect 523092 66988 523098 67040
rect 167730 66920 167736 66972
rect 167788 66960 167794 66972
rect 536834 66960 536840 66972
rect 167788 66932 536840 66960
rect 167788 66920 167794 66932
rect 536834 66920 536840 66932
rect 536892 66920 536898 66972
rect 170766 66852 170772 66904
rect 170824 66892 170830 66904
rect 550634 66892 550640 66904
rect 170824 66864 550640 66892
rect 170824 66852 170830 66864
rect 550634 66852 550640 66864
rect 550692 66852 550698 66904
rect 142706 65832 142712 65884
rect 142764 65872 142770 65884
rect 218054 65872 218060 65884
rect 142764 65844 218060 65872
rect 142764 65832 142770 65844
rect 218054 65832 218060 65844
rect 218112 65832 218118 65884
rect 154206 65764 154212 65816
rect 154264 65804 154270 65816
rect 332686 65804 332692 65816
rect 154264 65776 332692 65804
rect 154264 65764 154270 65776
rect 332686 65764 332692 65776
rect 332744 65764 332750 65816
rect 157978 65696 157984 65748
rect 158036 65736 158042 65748
rect 408494 65736 408500 65748
rect 158036 65708 408500 65736
rect 158036 65696 158042 65708
rect 408494 65696 408500 65708
rect 408552 65696 408558 65748
rect 167638 65628 167644 65680
rect 167696 65668 167702 65680
rect 539594 65668 539600 65680
rect 167696 65640 539600 65668
rect 167696 65628 167702 65640
rect 539594 65628 539600 65640
rect 539652 65628 539658 65680
rect 167546 65560 167552 65612
rect 167604 65600 167610 65612
rect 543734 65600 543740 65612
rect 167604 65572 543740 65600
rect 167604 65560 167610 65572
rect 543734 65560 543740 65572
rect 543792 65560 543798 65612
rect 170398 65492 170404 65544
rect 170456 65532 170462 65544
rect 568574 65532 568580 65544
rect 170456 65504 568580 65532
rect 170456 65492 170462 65504
rect 568574 65492 568580 65504
rect 568632 65492 568638 65544
rect 139946 64540 139952 64592
rect 140004 64580 140010 64592
rect 189074 64580 189080 64592
rect 140004 64552 189080 64580
rect 140004 64540 140010 64552
rect 189074 64540 189080 64552
rect 189132 64540 189138 64592
rect 141418 64472 141424 64524
rect 141476 64512 141482 64524
rect 207014 64512 207020 64524
rect 141476 64484 207020 64512
rect 141476 64472 141482 64484
rect 207014 64472 207020 64484
rect 207072 64472 207078 64524
rect 145650 64404 145656 64456
rect 145708 64444 145714 64456
rect 256694 64444 256700 64456
rect 145708 64416 256700 64444
rect 145708 64404 145714 64416
rect 256694 64404 256700 64416
rect 256752 64404 256758 64456
rect 147122 64336 147128 64388
rect 147180 64376 147186 64388
rect 270494 64376 270500 64388
rect 147180 64348 270500 64376
rect 147180 64336 147186 64348
rect 270494 64336 270500 64348
rect 270552 64336 270558 64388
rect 151078 64268 151084 64320
rect 151136 64308 151142 64320
rect 324314 64308 324320 64320
rect 151136 64280 324320 64308
rect 151136 64268 151142 64280
rect 324314 64268 324320 64280
rect 324372 64268 324378 64320
rect 162210 64200 162216 64252
rect 162268 64240 162274 64252
rect 368474 64240 368480 64252
rect 162268 64212 368480 64240
rect 162268 64200 162274 64212
rect 368474 64200 368480 64212
rect 368532 64200 368538 64252
rect 159358 64132 159364 64184
rect 159416 64172 159422 64184
rect 437474 64172 437480 64184
rect 159416 64144 437480 64172
rect 159416 64132 159422 64144
rect 437474 64132 437480 64144
rect 437532 64132 437538 64184
rect 139854 63112 139860 63164
rect 139912 63152 139918 63164
rect 185026 63152 185032 63164
rect 139912 63124 185032 63152
rect 139912 63112 139918 63124
rect 185026 63112 185032 63124
rect 185084 63112 185090 63164
rect 145558 63044 145564 63096
rect 145616 63084 145622 63096
rect 259454 63084 259460 63096
rect 145616 63056 259460 63084
rect 145616 63044 145622 63056
rect 259454 63044 259460 63056
rect 259512 63044 259518 63096
rect 161014 62976 161020 63028
rect 161072 63016 161078 63028
rect 347774 63016 347780 63028
rect 161072 62988 347780 63016
rect 161072 62976 161078 62988
rect 347774 62976 347780 62988
rect 347832 62976 347838 63028
rect 152366 62908 152372 62960
rect 152424 62948 152430 62960
rect 340966 62948 340972 62960
rect 152424 62920 340972 62948
rect 152424 62908 152430 62920
rect 340966 62908 340972 62920
rect 341024 62908 341030 62960
rect 155310 62840 155316 62892
rect 155368 62880 155374 62892
rect 376754 62880 376760 62892
rect 155368 62852 376760 62880
rect 155368 62840 155374 62852
rect 376754 62840 376760 62852
rect 376812 62840 376818 62892
rect 157886 62772 157892 62824
rect 157944 62812 157950 62824
rect 412634 62812 412640 62824
rect 157944 62784 412640 62812
rect 157944 62772 157950 62784
rect 412634 62772 412640 62784
rect 412692 62772 412698 62824
rect 138474 62160 138480 62212
rect 138532 62200 138538 62212
rect 140038 62200 140044 62212
rect 138532 62172 140044 62200
rect 138532 62160 138538 62172
rect 140038 62160 140044 62172
rect 140096 62160 140102 62212
rect 137278 62092 137284 62144
rect 137336 62132 137342 62144
rect 138658 62132 138664 62144
rect 137336 62104 138664 62132
rect 137336 62092 137342 62104
rect 138658 62092 138664 62104
rect 138716 62092 138722 62144
rect 144178 61820 144184 61872
rect 144236 61860 144242 61872
rect 234614 61860 234620 61872
rect 144236 61832 234620 61860
rect 144236 61820 144242 61832
rect 234614 61820 234620 61832
rect 234672 61820 234678 61872
rect 144270 61752 144276 61804
rect 144328 61792 144334 61804
rect 238754 61792 238760 61804
rect 144328 61764 238760 61792
rect 144328 61752 144334 61764
rect 238754 61752 238760 61764
rect 238812 61752 238818 61804
rect 147030 61684 147036 61736
rect 147088 61724 147094 61736
rect 274634 61724 274640 61736
rect 147088 61696 274640 61724
rect 147088 61684 147094 61696
rect 274634 61684 274640 61696
rect 274692 61684 274698 61736
rect 150986 61616 150992 61668
rect 151044 61656 151050 61668
rect 331214 61656 331220 61668
rect 151044 61628 331220 61656
rect 151044 61616 151050 61628
rect 331214 61616 331220 61628
rect 331272 61616 331278 61668
rect 153930 61548 153936 61600
rect 153988 61588 153994 61600
rect 358814 61588 358820 61600
rect 153988 61560 358820 61588
rect 153988 61548 153994 61560
rect 358814 61548 358820 61560
rect 358872 61548 358878 61600
rect 159266 61480 159272 61532
rect 159324 61520 159330 61532
rect 430574 61520 430580 61532
rect 159324 61492 430580 61520
rect 159324 61480 159330 61492
rect 430574 61480 430580 61492
rect 430632 61480 430638 61532
rect 166258 61412 166264 61464
rect 166316 61452 166322 61464
rect 516134 61452 516140 61464
rect 166316 61424 516140 61452
rect 166316 61412 166322 61424
rect 516134 61412 516140 61424
rect 516192 61412 516198 61464
rect 170306 61344 170312 61396
rect 170364 61384 170370 61396
rect 572714 61384 572720 61396
rect 170364 61356 572720 61384
rect 170364 61344 170370 61356
rect 572714 61344 572720 61356
rect 572772 61344 572778 61396
rect 118510 60664 118516 60716
rect 118568 60704 118574 60716
rect 580166 60704 580172 60716
rect 118568 60676 580172 60704
rect 118568 60664 118574 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 142614 60256 142620 60308
rect 142672 60296 142678 60308
rect 220814 60296 220820 60308
rect 142672 60268 220820 60296
rect 142672 60256 142678 60268
rect 220814 60256 220820 60268
rect 220872 60256 220878 60308
rect 148318 60188 148324 60240
rect 148376 60228 148382 60240
rect 292574 60228 292580 60240
rect 148376 60200 292580 60228
rect 148376 60188 148382 60200
rect 292574 60188 292580 60200
rect 292632 60188 292638 60240
rect 149698 60120 149704 60172
rect 149756 60160 149762 60172
rect 309134 60160 309140 60172
rect 149756 60132 309140 60160
rect 149756 60120 149762 60132
rect 309134 60120 309140 60132
rect 309192 60120 309198 60172
rect 153838 60052 153844 60104
rect 153896 60092 153902 60104
rect 356054 60092 356060 60104
rect 153896 60064 356060 60092
rect 153896 60052 153902 60064
rect 356054 60052 356060 60064
rect 356112 60052 356118 60104
rect 157794 59984 157800 60036
rect 157852 60024 157858 60036
rect 415394 60024 415400 60036
rect 157852 59996 415400 60024
rect 157852 59984 157858 59996
rect 415394 59984 415400 59996
rect 415452 59984 415458 60036
rect 162302 58760 162308 58812
rect 162360 58800 162366 58812
rect 354674 58800 354680 58812
rect 162360 58772 354680 58800
rect 162360 58760 162366 58772
rect 354674 58760 354680 58772
rect 354732 58760 354738 58812
rect 160646 58692 160652 58744
rect 160704 58732 160710 58744
rect 448514 58732 448520 58744
rect 160704 58704 448520 58732
rect 160704 58692 160710 58704
rect 448514 58692 448520 58704
rect 448572 58692 448578 58744
rect 163498 58624 163504 58676
rect 163556 58664 163562 58676
rect 481634 58664 481640 58676
rect 163556 58636 481640 58664
rect 163556 58624 163562 58636
rect 481634 58624 481640 58636
rect 481692 58624 481698 58676
rect 137186 57876 137192 57928
rect 137244 57916 137250 57928
rect 140130 57916 140136 57928
rect 137244 57888 140136 57916
rect 137244 57876 137250 57888
rect 140130 57876 140136 57888
rect 140188 57876 140194 57928
rect 155218 57332 155224 57384
rect 155276 57372 155282 57384
rect 373994 57372 374000 57384
rect 155276 57344 374000 57372
rect 155276 57332 155282 57344
rect 373994 57332 374000 57344
rect 374052 57332 374058 57384
rect 164878 57264 164884 57316
rect 164936 57304 164942 57316
rect 507854 57304 507860 57316
rect 164936 57276 507860 57304
rect 164936 57264 164942 57276
rect 507854 57264 507860 57276
rect 507912 57264 507918 57316
rect 166166 57196 166172 57248
rect 166224 57236 166230 57248
rect 525794 57236 525800 57248
rect 166224 57208 525800 57236
rect 166224 57196 166230 57208
rect 525794 57196 525800 57208
rect 525852 57196 525858 57248
rect 95234 55836 95240 55888
rect 95292 55876 95298 55888
rect 125318 55876 125324 55888
rect 95292 55848 125324 55876
rect 95292 55836 95298 55848
rect 125318 55836 125324 55848
rect 125376 55836 125382 55888
rect 152274 55836 152280 55888
rect 152332 55876 152338 55888
rect 338114 55876 338120 55888
rect 152332 55848 338120 55876
rect 152332 55836 152338 55848
rect 338114 55836 338120 55848
rect 338172 55836 338178 55888
rect 148226 54544 148232 54596
rect 148284 54584 148290 54596
rect 295334 54584 295340 54596
rect 148284 54556 295340 54584
rect 148284 54544 148290 54556
rect 295334 54544 295340 54556
rect 295392 54544 295398 54596
rect 102226 54476 102232 54528
rect 102284 54516 102290 54528
rect 125226 54516 125232 54528
rect 102284 54488 125232 54516
rect 102284 54476 102290 54488
rect 125226 54476 125232 54488
rect 125284 54476 125290 54528
rect 156598 54476 156604 54528
rect 156656 54516 156662 54528
rect 401594 54516 401600 54528
rect 156656 54488 401600 54516
rect 156656 54476 156662 54488
rect 401594 54476 401600 54488
rect 401652 54476 401658 54528
rect 149606 53048 149612 53100
rect 149664 53088 149670 53100
rect 316034 53088 316040 53100
rect 149664 53060 316040 53088
rect 149664 53048 149670 53060
rect 316034 53048 316040 53060
rect 316092 53048 316098 53100
rect 156506 50464 156512 50516
rect 156564 50504 156570 50516
rect 398834 50504 398840 50516
rect 156564 50476 398840 50504
rect 156564 50464 156570 50476
rect 398834 50464 398840 50476
rect 398892 50464 398898 50516
rect 161934 50396 161940 50448
rect 161992 50436 161998 50448
rect 469214 50436 469220 50448
rect 161992 50408 469220 50436
rect 161992 50396 161998 50408
rect 469214 50396 469220 50408
rect 469272 50396 469278 50448
rect 163406 50328 163412 50380
rect 163464 50368 163470 50380
rect 481726 50368 481732 50380
rect 163464 50340 481732 50368
rect 163464 50328 163470 50340
rect 481726 50328 481732 50340
rect 481784 50328 481790 50380
rect 182818 46860 182824 46912
rect 182876 46900 182882 46912
rect 580166 46900 580172 46912
rect 182876 46872 580172 46900
rect 182876 46860 182882 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 139762 46180 139768 46232
rect 139820 46220 139826 46232
rect 180794 46220 180800 46232
rect 139820 46192 180800 46220
rect 139820 46180 139826 46192
rect 180794 46180 180800 46192
rect 180852 46180 180858 46232
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 174630 45540 174636 45552
rect 3568 45512 174636 45540
rect 3568 45500 3574 45512
rect 174630 45500 174636 45512
rect 174688 45500 174694 45552
rect 35986 44820 35992 44872
rect 36044 44860 36050 44872
rect 127434 44860 127440 44872
rect 36044 44832 127440 44860
rect 36044 44820 36050 44832
rect 127434 44820 127440 44832
rect 127492 44820 127498 44872
rect 171502 42032 171508 42084
rect 171560 42072 171566 42084
rect 514846 42072 514852 42084
rect 171560 42044 514852 42072
rect 171560 42032 171566 42044
rect 514846 42032 514852 42044
rect 514904 42032 514910 42084
rect 120074 40264 120080 40316
rect 120132 40304 120138 40316
rect 123478 40304 123484 40316
rect 120132 40276 123484 40304
rect 120132 40264 120138 40276
rect 123478 40264 123484 40276
rect 123536 40264 123542 40316
rect 88334 36524 88340 36576
rect 88392 36564 88398 36576
rect 125134 36564 125140 36576
rect 88392 36536 125140 36564
rect 88392 36524 88398 36536
rect 125134 36524 125140 36536
rect 125192 36524 125198 36576
rect 145466 35572 145472 35624
rect 145524 35612 145530 35624
rect 262214 35612 262220 35624
rect 145524 35584 262220 35612
rect 145524 35572 145530 35584
rect 262214 35572 262220 35584
rect 262272 35572 262278 35624
rect 146938 35504 146944 35556
rect 146996 35544 147002 35556
rect 273254 35544 273260 35556
rect 146996 35516 273260 35544
rect 146996 35504 147002 35516
rect 273254 35504 273260 35516
rect 273312 35504 273318 35556
rect 146846 35436 146852 35488
rect 146904 35476 146910 35488
rect 276014 35476 276020 35488
rect 146904 35448 276020 35476
rect 146904 35436 146910 35448
rect 276014 35436 276020 35448
rect 276072 35436 276078 35488
rect 148134 35368 148140 35420
rect 148192 35408 148198 35420
rect 287054 35408 287060 35420
rect 148192 35380 287060 35408
rect 148192 35368 148198 35380
rect 287054 35368 287060 35380
rect 287112 35368 287118 35420
rect 149514 35300 149520 35352
rect 149572 35340 149578 35352
rect 307754 35340 307760 35352
rect 149572 35312 307760 35340
rect 149572 35300 149578 35312
rect 307754 35300 307760 35312
rect 307812 35300 307818 35352
rect 155034 35232 155040 35284
rect 155092 35272 155098 35284
rect 379514 35272 379520 35284
rect 155092 35244 379520 35272
rect 155092 35232 155098 35244
rect 379514 35232 379520 35244
rect 379572 35232 379578 35284
rect 155126 35164 155132 35216
rect 155184 35204 155190 35216
rect 386414 35204 386420 35216
rect 155184 35176 386420 35204
rect 155184 35164 155190 35176
rect 386414 35164 386420 35176
rect 386472 35164 386478 35216
rect 141234 34144 141240 34196
rect 141292 34184 141298 34196
rect 198734 34184 198740 34196
rect 141292 34156 198740 34184
rect 141292 34144 141298 34156
rect 198734 34144 198740 34156
rect 198792 34144 198798 34196
rect 142522 34076 142528 34128
rect 142580 34116 142586 34128
rect 219434 34116 219440 34128
rect 142580 34088 219440 34116
rect 142580 34076 142586 34088
rect 219434 34076 219440 34088
rect 219492 34076 219498 34128
rect 144086 34008 144092 34060
rect 144144 34048 144150 34060
rect 234706 34048 234712 34060
rect 144144 34020 234712 34048
rect 144144 34008 144150 34020
rect 234706 34008 234712 34020
rect 234764 34008 234770 34060
rect 145374 33940 145380 33992
rect 145432 33980 145438 33992
rect 251174 33980 251180 33992
rect 145432 33952 251180 33980
rect 145432 33940 145438 33952
rect 251174 33940 251180 33952
rect 251232 33940 251238 33992
rect 145282 33872 145288 33924
rect 145340 33912 145346 33924
rect 259546 33912 259552 33924
rect 145340 33884 259552 33912
rect 145340 33872 145346 33884
rect 259546 33872 259552 33884
rect 259604 33872 259610 33924
rect 141326 33804 141332 33856
rect 141384 33844 141390 33856
rect 201494 33844 201500 33856
rect 141384 33816 201500 33844
rect 141384 33804 141390 33816
rect 201494 33804 201500 33816
rect 201552 33804 201558 33856
rect 215938 33804 215944 33856
rect 215996 33844 216002 33856
rect 456794 33844 456800 33856
rect 215996 33816 456800 33844
rect 215996 33804 216002 33816
rect 456794 33804 456800 33816
rect 456852 33804 456858 33856
rect 170214 33736 170220 33788
rect 170272 33776 170278 33788
rect 574094 33776 574100 33788
rect 170272 33748 574100 33776
rect 170272 33736 170278 33748
rect 574094 33736 574100 33748
rect 574152 33736 574158 33788
rect 170122 33056 170128 33108
rect 170180 33096 170186 33108
rect 580166 33096 580172 33108
rect 170180 33068 580172 33096
rect 170180 33056 170186 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 3510 32988 3516 33040
rect 3568 33028 3574 33040
rect 180886 33028 180892 33040
rect 3568 33000 180892 33028
rect 3568 32988 3574 33000
rect 180886 32988 180892 33000
rect 180944 32988 180950 33040
rect 174538 32580 174544 32632
rect 174596 32620 174602 32632
rect 425054 32620 425060 32632
rect 174596 32592 425060 32620
rect 174596 32580 174602 32592
rect 425054 32580 425060 32592
rect 425112 32580 425118 32632
rect 163314 32512 163320 32564
rect 163372 32552 163378 32564
rect 485774 32552 485780 32564
rect 163372 32524 485780 32552
rect 163372 32512 163378 32524
rect 485774 32512 485780 32524
rect 485832 32512 485838 32564
rect 167454 32444 167460 32496
rect 167512 32484 167518 32496
rect 542354 32484 542360 32496
rect 167512 32456 542360 32484
rect 167512 32444 167518 32456
rect 542354 32444 542360 32456
rect 542412 32444 542418 32496
rect 170030 32376 170036 32428
rect 170088 32416 170094 32428
rect 571334 32416 571340 32428
rect 170088 32388 571340 32416
rect 170088 32376 170094 32388
rect 571334 32376 571340 32388
rect 571392 32376 571398 32428
rect 149330 31492 149336 31544
rect 149388 31532 149394 31544
rect 303614 31532 303620 31544
rect 149388 31504 303620 31532
rect 149388 31492 149394 31504
rect 303614 31492 303620 31504
rect 303672 31492 303678 31544
rect 149422 31424 149428 31476
rect 149480 31464 149486 31476
rect 307846 31464 307852 31476
rect 149480 31436 307852 31464
rect 149480 31424 149486 31436
rect 307846 31424 307852 31436
rect 307904 31424 307910 31476
rect 150894 31356 150900 31408
rect 150952 31396 150958 31408
rect 321554 31396 321560 31408
rect 150952 31368 321560 31396
rect 150952 31356 150958 31368
rect 321554 31356 321560 31368
rect 321612 31356 321618 31408
rect 154942 31288 154948 31340
rect 155000 31328 155006 31340
rect 385034 31328 385040 31340
rect 155000 31300 385040 31328
rect 155000 31288 155006 31300
rect 385034 31288 385040 31300
rect 385092 31288 385098 31340
rect 159174 31220 159180 31272
rect 159232 31260 159238 31272
rect 434714 31260 434720 31272
rect 159232 31232 434720 31260
rect 159232 31220 159238 31232
rect 434714 31220 434720 31232
rect 434772 31220 434778 31272
rect 164786 31152 164792 31204
rect 164844 31192 164850 31204
rect 506474 31192 506480 31204
rect 164844 31164 506480 31192
rect 164844 31152 164850 31164
rect 506474 31152 506480 31164
rect 506532 31152 506538 31204
rect 166074 31084 166080 31136
rect 166132 31124 166138 31136
rect 517514 31124 517520 31136
rect 166132 31096 517520 31124
rect 166132 31084 166138 31096
rect 517514 31084 517520 31096
rect 517572 31084 517578 31136
rect 165982 31016 165988 31068
rect 166040 31056 166046 31068
rect 521654 31056 521660 31068
rect 166040 31028 521660 31056
rect 166040 31016 166046 31028
rect 521654 31016 521660 31028
rect 521712 31016 521718 31068
rect 143994 30064 144000 30116
rect 144052 30104 144058 30116
rect 233234 30104 233240 30116
rect 144052 30076 233240 30104
rect 144052 30064 144058 30076
rect 233234 30064 233240 30076
rect 233292 30064 233298 30116
rect 143902 29996 143908 30048
rect 143960 30036 143966 30048
rect 235994 30036 236000 30048
rect 143960 30008 236000 30036
rect 143960 29996 143966 30008
rect 235994 29996 236000 30008
rect 236052 29996 236058 30048
rect 145190 29928 145196 29980
rect 145248 29968 145254 29980
rect 251266 29968 251272 29980
rect 145248 29940 251272 29968
rect 145248 29928 145254 29940
rect 251266 29928 251272 29940
rect 251324 29928 251330 29980
rect 146754 29860 146760 29912
rect 146812 29900 146818 29912
rect 267826 29900 267832 29912
rect 146812 29872 267832 29900
rect 146812 29860 146818 29872
rect 267826 29860 267832 29872
rect 267884 29860 267890 29912
rect 147950 29792 147956 29844
rect 148008 29832 148014 29844
rect 285674 29832 285680 29844
rect 148008 29804 285680 29832
rect 148008 29792 148014 29804
rect 285674 29792 285680 29804
rect 285732 29792 285738 29844
rect 148042 29724 148048 29776
rect 148100 29764 148106 29776
rect 289814 29764 289820 29776
rect 148100 29736 289820 29764
rect 148100 29724 148106 29736
rect 289814 29724 289820 29736
rect 289872 29724 289878 29776
rect 154850 29656 154856 29708
rect 154908 29696 154914 29708
rect 374086 29696 374092 29708
rect 154908 29668 374092 29696
rect 154908 29656 154914 29668
rect 374086 29656 374092 29668
rect 374144 29656 374150 29708
rect 161842 29588 161848 29640
rect 161900 29628 161906 29640
rect 466454 29628 466460 29640
rect 161900 29600 466460 29628
rect 161900 29588 161906 29600
rect 466454 29588 466460 29600
rect 466512 29588 466518 29640
rect 141142 28704 141148 28756
rect 141200 28744 141206 28756
rect 208394 28744 208400 28756
rect 141200 28716 208400 28744
rect 141200 28704 141206 28716
rect 208394 28704 208400 28716
rect 208452 28704 208458 28756
rect 142430 28636 142436 28688
rect 142488 28676 142494 28688
rect 215294 28676 215300 28688
rect 142488 28648 215300 28676
rect 142488 28636 142494 28648
rect 215294 28636 215300 28648
rect 215352 28636 215358 28688
rect 142246 28568 142252 28620
rect 142304 28608 142310 28620
rect 218146 28608 218152 28620
rect 142304 28580 218152 28608
rect 142304 28568 142310 28580
rect 218146 28568 218152 28580
rect 218204 28568 218210 28620
rect 142338 28500 142344 28552
rect 142396 28540 142402 28552
rect 222194 28540 222200 28552
rect 142396 28512 222200 28540
rect 142396 28500 142402 28512
rect 222194 28500 222200 28512
rect 222252 28500 222258 28552
rect 143810 28432 143816 28484
rect 143868 28472 143874 28484
rect 242894 28472 242900 28484
rect 143868 28444 242900 28472
rect 143868 28432 143874 28444
rect 242894 28432 242900 28444
rect 242952 28432 242958 28484
rect 145098 28364 145104 28416
rect 145156 28404 145162 28416
rect 258074 28404 258080 28416
rect 145156 28376 258080 28404
rect 145156 28364 145162 28376
rect 258074 28364 258080 28376
rect 258132 28364 258138 28416
rect 161750 28296 161756 28348
rect 161808 28336 161814 28348
rect 463694 28336 463700 28348
rect 161808 28308 463700 28336
rect 161808 28296 161814 28308
rect 463694 28296 463700 28308
rect 463752 28296 463758 28348
rect 165890 28228 165896 28280
rect 165948 28268 165954 28280
rect 524414 28268 524420 28280
rect 165948 28240 524420 28268
rect 165948 28228 165954 28240
rect 524414 28228 524420 28240
rect 524472 28228 524478 28280
rect 141050 27276 141056 27328
rect 141108 27316 141114 27328
rect 201586 27316 201592 27328
rect 141108 27288 201592 27316
rect 141108 27276 141114 27288
rect 201586 27276 201592 27288
rect 201644 27276 201650 27328
rect 140958 27208 140964 27260
rect 141016 27248 141022 27260
rect 204254 27248 204260 27260
rect 141016 27220 204260 27248
rect 141016 27208 141022 27220
rect 204254 27208 204260 27220
rect 204312 27208 204318 27260
rect 145006 27140 145012 27192
rect 145064 27180 145070 27192
rect 253934 27180 253940 27192
rect 145064 27152 253940 27180
rect 145064 27140 145070 27152
rect 253934 27140 253940 27152
rect 253992 27140 253998 27192
rect 146662 27072 146668 27124
rect 146720 27112 146726 27124
rect 271874 27112 271880 27124
rect 146720 27084 271880 27112
rect 146720 27072 146726 27084
rect 271874 27072 271880 27084
rect 271932 27072 271938 27124
rect 153746 27004 153752 27056
rect 153804 27044 153810 27056
rect 357434 27044 357440 27056
rect 153804 27016 357440 27044
rect 153804 27004 153810 27016
rect 357434 27004 357440 27016
rect 357492 27004 357498 27056
rect 160554 26936 160560 26988
rect 160612 26976 160618 26988
rect 447134 26976 447140 26988
rect 160612 26948 447140 26976
rect 160612 26936 160618 26948
rect 447134 26936 447140 26948
rect 447192 26936 447198 26988
rect 161658 26868 161664 26920
rect 161716 26908 161722 26920
rect 470594 26908 470600 26920
rect 161716 26880 470600 26908
rect 161716 26868 161722 26880
rect 470594 26868 470600 26880
rect 470652 26868 470658 26920
rect 140406 25984 140412 26036
rect 140464 26024 140470 26036
rect 176746 26024 176752 26036
rect 140464 25996 176752 26024
rect 140464 25984 140470 25996
rect 176746 25984 176752 25996
rect 176804 25984 176810 26036
rect 139486 25916 139492 25968
rect 139544 25956 139550 25968
rect 179414 25956 179420 25968
rect 139544 25928 179420 25956
rect 139544 25916 139550 25928
rect 179414 25916 179420 25928
rect 179472 25916 179478 25968
rect 139670 25848 139676 25900
rect 139728 25888 139734 25900
rect 183554 25888 183560 25900
rect 139728 25860 183560 25888
rect 139728 25848 139734 25860
rect 183554 25848 183560 25860
rect 183612 25848 183618 25900
rect 139578 25780 139584 25832
rect 139636 25820 139642 25832
rect 186314 25820 186320 25832
rect 139636 25792 186320 25820
rect 139636 25780 139642 25792
rect 186314 25780 186320 25792
rect 186372 25780 186378 25832
rect 146570 25712 146576 25764
rect 146628 25752 146634 25764
rect 278774 25752 278780 25764
rect 146628 25724 278780 25752
rect 146628 25712 146634 25724
rect 278774 25712 278780 25724
rect 278832 25712 278838 25764
rect 152182 25644 152188 25696
rect 152240 25684 152246 25696
rect 346394 25684 346400 25696
rect 152240 25656 346400 25684
rect 152240 25644 152246 25656
rect 346394 25644 346400 25656
rect 346452 25644 346458 25696
rect 164602 25576 164608 25628
rect 164660 25616 164666 25628
rect 499574 25616 499580 25628
rect 164660 25588 499580 25616
rect 164660 25576 164666 25588
rect 499574 25576 499580 25588
rect 499632 25576 499638 25628
rect 164694 25508 164700 25560
rect 164752 25548 164758 25560
rect 503714 25548 503720 25560
rect 164752 25520 503720 25548
rect 164752 25508 164758 25520
rect 503714 25508 503720 25520
rect 503772 25508 503778 25560
rect 139394 24488 139400 24540
rect 139452 24528 139458 24540
rect 187694 24528 187700 24540
rect 139452 24500 187700 24528
rect 139452 24488 139458 24500
rect 187694 24488 187700 24500
rect 187752 24488 187758 24540
rect 150802 24420 150808 24472
rect 150860 24460 150866 24472
rect 324406 24460 324412 24472
rect 150860 24432 324412 24460
rect 150860 24420 150866 24432
rect 324406 24420 324412 24432
rect 324464 24420 324470 24472
rect 171686 24352 171692 24404
rect 171744 24392 171750 24404
rect 440234 24392 440240 24404
rect 171744 24364 440240 24392
rect 171744 24352 171750 24364
rect 440234 24352 440240 24364
rect 440292 24352 440298 24404
rect 168926 24284 168932 24336
rect 168984 24324 168990 24336
rect 552014 24324 552020 24336
rect 168984 24296 552020 24324
rect 168984 24284 168990 24296
rect 552014 24284 552020 24296
rect 552072 24284 552078 24336
rect 168834 24216 168840 24268
rect 168892 24256 168898 24268
rect 556154 24256 556160 24268
rect 168892 24228 556160 24256
rect 168892 24216 168898 24228
rect 556154 24216 556160 24228
rect 556212 24216 556218 24268
rect 168742 24148 168748 24200
rect 168800 24188 168806 24200
rect 563054 24188 563060 24200
rect 168800 24160 563060 24188
rect 168800 24148 168806 24160
rect 563054 24148 563060 24160
rect 563112 24148 563118 24200
rect 169938 24080 169944 24132
rect 169996 24120 170002 24132
rect 572806 24120 572812 24132
rect 169996 24092 572812 24120
rect 169996 24080 170002 24092
rect 572806 24080 572812 24092
rect 572864 24080 572870 24132
rect 3510 23196 3516 23248
rect 3568 23236 3574 23248
rect 174354 23236 174360 23248
rect 3568 23208 174360 23236
rect 3568 23196 3574 23208
rect 174354 23196 174360 23208
rect 174412 23196 174418 23248
rect 150710 23128 150716 23180
rect 150768 23168 150774 23180
rect 329834 23168 329840 23180
rect 150768 23140 329840 23168
rect 150768 23128 150774 23140
rect 329834 23128 329840 23140
rect 329892 23128 329898 23180
rect 157702 23060 157708 23112
rect 157760 23100 157766 23112
rect 415486 23100 415492 23112
rect 157760 23072 415492 23100
rect 157760 23060 157766 23072
rect 415486 23060 415492 23072
rect 415544 23060 415550 23112
rect 167362 22992 167368 23044
rect 167420 23032 167426 23044
rect 534074 23032 534080 23044
rect 167420 23004 534080 23032
rect 167420 22992 167426 23004
rect 534074 22992 534080 23004
rect 534132 22992 534138 23044
rect 167270 22924 167276 22976
rect 167328 22964 167334 22976
rect 538214 22964 538220 22976
rect 167328 22936 538220 22964
rect 167328 22924 167334 22936
rect 538214 22924 538220 22936
rect 538272 22924 538278 22976
rect 167178 22856 167184 22908
rect 167236 22896 167242 22908
rect 540974 22896 540980 22908
rect 167236 22868 540980 22896
rect 167236 22856 167242 22868
rect 540974 22856 540980 22868
rect 541032 22856 541038 22908
rect 52454 22788 52460 22840
rect 52512 22828 52518 22840
rect 128722 22828 128728 22840
rect 52512 22800 128728 22828
rect 52512 22788 52518 22800
rect 128722 22788 128728 22800
rect 128780 22788 128786 22840
rect 169846 22788 169852 22840
rect 169904 22828 169910 22840
rect 569954 22828 569960 22840
rect 169904 22800 569960 22828
rect 169904 22788 169910 22800
rect 569954 22788 569960 22800
rect 570012 22788 570018 22840
rect 118418 22720 118424 22772
rect 118476 22760 118482 22772
rect 580166 22760 580172 22772
rect 118476 22732 580172 22760
rect 118476 22720 118482 22732
rect 580166 22720 580172 22732
rect 580224 22720 580230 22772
rect 158346 21768 158352 21820
rect 158404 21808 158410 21820
rect 361574 21808 361580 21820
rect 158404 21780 361580 21808
rect 158404 21768 158410 21780
rect 361574 21768 361580 21780
rect 361632 21768 361638 21820
rect 173434 21700 173440 21752
rect 173492 21740 173498 21752
rect 432046 21740 432052 21752
rect 173492 21712 432052 21740
rect 173492 21700 173498 21712
rect 432046 21700 432052 21712
rect 432104 21700 432110 21752
rect 158990 21632 158996 21684
rect 159048 21672 159054 21684
rect 429194 21672 429200 21684
rect 159048 21644 429200 21672
rect 159048 21632 159054 21644
rect 429194 21632 429200 21644
rect 429252 21632 429258 21684
rect 159082 21564 159088 21616
rect 159140 21604 159146 21616
rect 436094 21604 436100 21616
rect 159140 21576 436100 21604
rect 159140 21564 159146 21576
rect 436094 21564 436100 21576
rect 436152 21564 436158 21616
rect 165706 21496 165712 21548
rect 165764 21536 165770 21548
rect 520274 21536 520280 21548
rect 165764 21508 520280 21536
rect 165764 21496 165770 21508
rect 520274 21496 520280 21508
rect 520332 21496 520338 21548
rect 165798 21428 165804 21480
rect 165856 21468 165862 21480
rect 523126 21468 523132 21480
rect 165856 21440 523132 21468
rect 165856 21428 165862 21440
rect 523126 21428 523132 21440
rect 523184 21428 523190 21480
rect 45554 21360 45560 21412
rect 45612 21400 45618 21412
rect 120810 21400 120816 21412
rect 45612 21372 120816 21400
rect 45612 21360 45618 21372
rect 120810 21360 120816 21372
rect 120868 21360 120874 21412
rect 165614 21360 165620 21412
rect 165672 21400 165678 21412
rect 527174 21400 527180 21412
rect 165672 21372 527180 21400
rect 165672 21360 165678 21372
rect 527174 21360 527180 21372
rect 527232 21360 527238 21412
rect 135990 20612 135996 20664
rect 136048 20652 136054 20664
rect 142246 20652 142252 20664
rect 136048 20624 142252 20652
rect 136048 20612 136054 20624
rect 142246 20612 142252 20624
rect 142304 20612 142310 20664
rect 144914 20340 144920 20392
rect 144972 20380 144978 20392
rect 255314 20380 255320 20392
rect 144972 20352 255320 20380
rect 144972 20340 144978 20352
rect 255314 20340 255320 20352
rect 255372 20340 255378 20392
rect 146478 20272 146484 20324
rect 146536 20312 146542 20324
rect 269114 20312 269120 20324
rect 146536 20284 269120 20312
rect 146536 20272 146542 20284
rect 269114 20272 269120 20284
rect 269172 20272 269178 20324
rect 143718 20204 143724 20256
rect 143776 20244 143782 20256
rect 241514 20244 241520 20256
rect 143776 20216 241520 20244
rect 143776 20204 143782 20216
rect 241514 20204 241520 20216
rect 241572 20204 241578 20256
rect 242158 20204 242164 20256
rect 242216 20244 242222 20256
rect 449894 20244 449900 20256
rect 242216 20216 449900 20244
rect 242216 20204 242222 20216
rect 449894 20204 449900 20216
rect 449952 20204 449958 20256
rect 173342 20136 173348 20188
rect 173400 20176 173406 20188
rect 418154 20176 418160 20188
rect 173400 20148 418160 20176
rect 173400 20136 173406 20148
rect 418154 20136 418160 20148
rect 418212 20136 418218 20188
rect 163130 20068 163136 20120
rect 163188 20108 163194 20120
rect 484394 20108 484400 20120
rect 163188 20080 484400 20108
rect 163188 20068 163194 20080
rect 484394 20068 484400 20080
rect 484452 20068 484458 20120
rect 106274 20000 106280 20052
rect 106332 20040 106338 20052
rect 133046 20040 133052 20052
rect 106332 20012 133052 20040
rect 106332 20000 106338 20012
rect 133046 20000 133052 20012
rect 133104 20000 133110 20052
rect 163222 20000 163228 20052
rect 163280 20040 163286 20052
rect 488534 20040 488540 20052
rect 163280 20012 488540 20040
rect 163280 20000 163286 20012
rect 488534 20000 488540 20012
rect 488592 20000 488598 20052
rect 70394 19932 70400 19984
rect 70452 19972 70458 19984
rect 130286 19972 130292 19984
rect 70452 19944 130292 19972
rect 70452 19932 70458 19944
rect 130286 19932 130292 19944
rect 130344 19932 130350 19984
rect 164510 19932 164516 19984
rect 164568 19972 164574 19984
rect 498286 19972 498292 19984
rect 164568 19944 498292 19972
rect 164568 19932 164574 19944
rect 498286 19932 498292 19944
rect 498344 19932 498350 19984
rect 150618 18912 150624 18964
rect 150676 18952 150682 18964
rect 322934 18952 322940 18964
rect 150676 18924 322940 18952
rect 150676 18912 150682 18924
rect 322934 18912 322940 18924
rect 322992 18912 322998 18964
rect 172422 18844 172428 18896
rect 172480 18884 172486 18896
rect 411254 18884 411260 18896
rect 172480 18856 411260 18884
rect 172480 18844 172486 18856
rect 411254 18844 411260 18856
rect 411312 18844 411318 18896
rect 161566 18776 161572 18828
rect 161624 18816 161630 18828
rect 465166 18816 465172 18828
rect 161624 18788 465172 18816
rect 161624 18776 161630 18788
rect 465166 18776 465172 18788
rect 465224 18776 465230 18828
rect 168466 18708 168472 18760
rect 168524 18748 168530 18760
rect 553394 18748 553400 18760
rect 168524 18720 553400 18748
rect 168524 18708 168530 18720
rect 553394 18708 553400 18720
rect 553452 18708 553458 18760
rect 168558 18640 168564 18692
rect 168616 18680 168622 18692
rect 556246 18680 556252 18692
rect 168616 18652 556252 18680
rect 168616 18640 168622 18652
rect 556246 18640 556252 18652
rect 556304 18640 556310 18692
rect 4154 18572 4160 18624
rect 4212 18612 4218 18624
rect 126146 18612 126152 18624
rect 4212 18584 126152 18612
rect 4212 18572 4218 18584
rect 126146 18572 126152 18584
rect 126204 18572 126210 18624
rect 168650 18572 168656 18624
rect 168708 18612 168714 18624
rect 560294 18612 560300 18624
rect 168708 18584 560300 18612
rect 168708 18572 168714 18584
rect 560294 18572 560300 18584
rect 560352 18572 560358 18624
rect 140866 17620 140872 17672
rect 140924 17660 140930 17672
rect 205634 17660 205640 17672
rect 140924 17632 205640 17660
rect 140924 17620 140930 17632
rect 205634 17620 205640 17632
rect 205692 17620 205698 17672
rect 158898 17552 158904 17604
rect 158956 17592 158962 17604
rect 433334 17592 433340 17604
rect 158956 17564 433340 17592
rect 158956 17552 158962 17564
rect 433334 17552 433340 17564
rect 433392 17552 433398 17604
rect 158806 17484 158812 17536
rect 158864 17524 158870 17536
rect 440326 17524 440332 17536
rect 158864 17496 440332 17524
rect 158864 17484 158870 17496
rect 440326 17484 440332 17496
rect 440384 17484 440390 17536
rect 160278 17416 160284 17468
rect 160336 17456 160342 17468
rect 448606 17456 448612 17468
rect 160336 17428 448612 17456
rect 160336 17416 160342 17428
rect 448606 17416 448612 17428
rect 448664 17416 448670 17468
rect 160462 17348 160468 17400
rect 160520 17388 160526 17400
rect 451274 17388 451280 17400
rect 160520 17360 451280 17388
rect 160520 17348 160526 17360
rect 451274 17348 451280 17360
rect 451332 17348 451338 17400
rect 160186 17280 160192 17332
rect 160244 17320 160250 17332
rect 452654 17320 452660 17332
rect 160244 17292 452660 17320
rect 160244 17280 160250 17292
rect 452654 17280 452660 17292
rect 452712 17280 452718 17332
rect 38654 17212 38660 17264
rect 38712 17252 38718 17264
rect 120718 17252 120724 17264
rect 38712 17224 120724 17252
rect 38712 17212 38718 17224
rect 120718 17212 120724 17224
rect 120776 17212 120782 17264
rect 160370 17212 160376 17264
rect 160428 17252 160434 17264
rect 455414 17252 455420 17264
rect 160428 17224 455420 17252
rect 160428 17212 160434 17224
rect 455414 17212 455420 17224
rect 455472 17212 455478 17264
rect 147858 16124 147864 16176
rect 147916 16164 147922 16176
rect 294874 16164 294880 16176
rect 147916 16136 294880 16164
rect 147916 16124 147922 16136
rect 294874 16124 294880 16136
rect 294932 16124 294938 16176
rect 154758 16056 154764 16108
rect 154816 16096 154822 16108
rect 378410 16096 378416 16108
rect 154816 16068 378416 16096
rect 154816 16056 154822 16068
rect 378410 16056 378416 16068
rect 378468 16056 378474 16108
rect 156414 15988 156420 16040
rect 156472 16028 156478 16040
rect 395338 16028 395344 16040
rect 156472 16000 395344 16028
rect 156472 15988 156478 16000
rect 395338 15988 395344 16000
rect 395396 15988 395402 16040
rect 157610 15920 157616 15972
rect 157668 15960 157674 15972
rect 420178 15960 420184 15972
rect 157668 15932 420184 15960
rect 157668 15920 157674 15932
rect 420178 15920 420184 15932
rect 420236 15920 420242 15972
rect 14274 15852 14280 15904
rect 14332 15892 14338 15904
rect 125042 15892 125048 15904
rect 14332 15864 125048 15892
rect 14332 15852 14338 15864
rect 125042 15852 125048 15864
rect 125100 15852 125106 15904
rect 164418 15852 164424 15904
rect 164476 15892 164482 15904
rect 509602 15892 509608 15904
rect 164476 15864 509608 15892
rect 164476 15852 164482 15864
rect 509602 15852 509608 15864
rect 509660 15852 509666 15904
rect 143626 14696 143632 14748
rect 143684 14736 143690 14748
rect 237650 14736 237656 14748
rect 143684 14708 237656 14736
rect 143684 14696 143690 14708
rect 237650 14696 237656 14708
rect 237708 14696 237714 14748
rect 152090 14628 152096 14680
rect 152148 14668 152154 14680
rect 342898 14668 342904 14680
rect 152148 14640 342904 14668
rect 152148 14628 152154 14640
rect 342898 14628 342904 14640
rect 342956 14628 342962 14680
rect 154666 14560 154672 14612
rect 154724 14600 154730 14612
rect 384298 14600 384304 14612
rect 154724 14572 384304 14600
rect 154724 14560 154730 14572
rect 384298 14560 384304 14572
rect 384356 14560 384362 14612
rect 172330 14492 172336 14544
rect 172388 14532 172394 14544
rect 404354 14532 404360 14544
rect 172388 14504 404360 14532
rect 172388 14492 172394 14504
rect 404354 14492 404360 14504
rect 404412 14492 404418 14544
rect 31938 14424 31944 14476
rect 31996 14464 32002 14476
rect 122190 14464 122196 14476
rect 31996 14436 122196 14464
rect 31996 14424 32002 14436
rect 122190 14424 122196 14436
rect 122248 14424 122254 14476
rect 156322 14424 156328 14476
rect 156380 14464 156386 14476
rect 390646 14464 390652 14476
rect 156380 14436 390652 14464
rect 156380 14424 156386 14436
rect 390646 14424 390652 14436
rect 390704 14424 390710 14476
rect 147766 13540 147772 13592
rect 147824 13580 147830 13592
rect 291378 13580 291384 13592
rect 147824 13552 291384 13580
rect 147824 13540 147830 13552
rect 291378 13540 291384 13552
rect 291436 13540 291442 13592
rect 151998 13472 152004 13524
rect 152056 13512 152062 13524
rect 339494 13512 339500 13524
rect 152056 13484 339500 13512
rect 152056 13472 152062 13484
rect 339494 13472 339500 13484
rect 339552 13472 339558 13524
rect 153654 13404 153660 13456
rect 153712 13444 153718 13456
rect 365714 13444 365720 13456
rect 153712 13416 365720 13444
rect 153712 13404 153718 13416
rect 365714 13404 365720 13416
rect 365772 13404 365778 13456
rect 154574 13336 154580 13388
rect 154632 13376 154638 13388
rect 381170 13376 381176 13388
rect 154632 13348 381176 13376
rect 154632 13336 154638 13348
rect 381170 13336 381176 13348
rect 381228 13336 381234 13388
rect 156230 13268 156236 13320
rect 156288 13308 156294 13320
rect 392578 13308 392584 13320
rect 156288 13280 392584 13308
rect 156288 13268 156294 13280
rect 392578 13268 392584 13280
rect 392636 13268 392642 13320
rect 156138 13200 156144 13252
rect 156196 13240 156202 13252
rect 400858 13240 400864 13252
rect 156196 13212 400864 13240
rect 156196 13200 156202 13212
rect 400858 13200 400864 13212
rect 400916 13200 400922 13252
rect 157518 13132 157524 13184
rect 157576 13172 157582 13184
rect 410794 13172 410800 13184
rect 157576 13144 410800 13172
rect 157576 13132 157582 13144
rect 410794 13132 410800 13144
rect 410852 13132 410858 13184
rect 164326 13064 164332 13116
rect 164384 13104 164390 13116
rect 506566 13104 506572 13116
rect 164384 13076 506572 13104
rect 164384 13064 164390 13076
rect 506566 13064 506572 13076
rect 506624 13064 506630 13116
rect 151906 11908 151912 11960
rect 151964 11948 151970 11960
rect 349246 11948 349252 11960
rect 151964 11920 349252 11948
rect 151964 11908 151970 11920
rect 349246 11908 349252 11920
rect 349304 11908 349310 11960
rect 153562 11840 153568 11892
rect 153620 11880 153626 11892
rect 361114 11880 361120 11892
rect 153620 11852 361120 11880
rect 153620 11840 153626 11852
rect 361114 11840 361120 11852
rect 361172 11840 361178 11892
rect 153470 11772 153476 11824
rect 153528 11812 153534 11824
rect 363506 11812 363512 11824
rect 153528 11784 363512 11812
rect 153528 11772 153534 11784
rect 363506 11772 363512 11784
rect 363564 11772 363570 11824
rect 117314 11704 117320 11756
rect 117372 11744 117378 11756
rect 134150 11744 134156 11756
rect 117372 11716 134156 11744
rect 117372 11704 117378 11716
rect 134150 11704 134156 11716
rect 134208 11704 134214 11756
rect 153378 11704 153384 11756
rect 153436 11744 153442 11756
rect 364610 11744 364616 11756
rect 153436 11716 364616 11744
rect 153436 11704 153442 11716
rect 364610 11704 364616 11716
rect 364668 11704 364674 11756
rect 176654 11636 176660 11688
rect 176712 11676 176718 11688
rect 177850 11676 177856 11688
rect 176712 11648 177856 11676
rect 176712 11636 176718 11648
rect 177850 11636 177856 11648
rect 177908 11636 177914 11688
rect 201494 11636 201500 11688
rect 201552 11676 201558 11688
rect 202690 11676 202696 11688
rect 201552 11648 202696 11676
rect 201552 11636 201558 11648
rect 202690 11636 202696 11648
rect 202748 11636 202754 11688
rect 234614 11636 234620 11688
rect 234672 11676 234678 11688
rect 235810 11676 235816 11688
rect 234672 11648 235816 11676
rect 234672 11636 234678 11648
rect 235810 11636 235816 11648
rect 235868 11636 235874 11688
rect 259454 11636 259460 11688
rect 259512 11676 259518 11688
rect 260650 11676 260656 11688
rect 259512 11648 260656 11676
rect 259512 11636 259518 11648
rect 260650 11636 260656 11648
rect 260708 11636 260714 11688
rect 149238 10684 149244 10736
rect 149296 10724 149302 10736
rect 314654 10724 314660 10736
rect 149296 10696 314660 10724
rect 149296 10684 149302 10696
rect 314654 10684 314660 10696
rect 314712 10684 314718 10736
rect 99834 10616 99840 10668
rect 99892 10656 99898 10668
rect 132954 10656 132960 10668
rect 99892 10628 132960 10656
rect 99892 10616 99898 10628
rect 132954 10616 132960 10628
rect 133012 10616 133018 10668
rect 150526 10616 150532 10668
rect 150584 10656 150590 10668
rect 327994 10656 328000 10668
rect 150584 10628 328000 10656
rect 150584 10616 150590 10628
rect 327994 10616 328000 10628
rect 328052 10616 328058 10668
rect 81618 10548 81624 10600
rect 81676 10588 81682 10600
rect 131758 10588 131764 10600
rect 81676 10560 131764 10588
rect 81676 10548 81682 10560
rect 131758 10548 131764 10560
rect 131816 10548 131822 10600
rect 151814 10548 151820 10600
rect 151872 10588 151878 10600
rect 345290 10588 345296 10600
rect 151872 10560 345296 10588
rect 151872 10548 151878 10560
rect 345290 10548 345296 10560
rect 345348 10548 345354 10600
rect 78122 10480 78128 10532
rect 78180 10520 78186 10532
rect 128446 10520 128452 10532
rect 78180 10492 128452 10520
rect 78180 10480 78186 10492
rect 128446 10480 128452 10492
rect 128504 10480 128510 10532
rect 172238 10480 172244 10532
rect 172296 10520 172302 10532
rect 397730 10520 397736 10532
rect 172296 10492 397736 10520
rect 172296 10480 172302 10492
rect 397730 10480 397736 10492
rect 397788 10480 397794 10532
rect 67634 10412 67640 10464
rect 67692 10452 67698 10464
rect 130194 10452 130200 10464
rect 67692 10424 130200 10452
rect 67692 10412 67698 10424
rect 130194 10412 130200 10424
rect 130252 10412 130258 10464
rect 158714 10412 158720 10464
rect 158772 10452 158778 10464
rect 428458 10452 428464 10464
rect 158772 10424 428464 10452
rect 158772 10412 158778 10424
rect 428458 10412 428464 10424
rect 428516 10412 428522 10464
rect 64322 10344 64328 10396
rect 64380 10384 64386 10396
rect 126330 10384 126336 10396
rect 64380 10356 126336 10384
rect 64380 10344 64386 10356
rect 126330 10344 126336 10356
rect 126388 10344 126394 10396
rect 164234 10344 164240 10396
rect 164292 10384 164298 10396
rect 502978 10384 502984 10396
rect 164292 10356 502984 10384
rect 164292 10344 164298 10356
rect 502978 10344 502984 10356
rect 503036 10344 503042 10396
rect 25314 10276 25320 10328
rect 25372 10316 25378 10328
rect 57238 10316 57244 10328
rect 25372 10288 57244 10316
rect 25372 10276 25378 10288
rect 57238 10276 57244 10288
rect 57296 10276 57302 10328
rect 60826 10276 60832 10328
rect 60884 10316 60890 10328
rect 129090 10316 129096 10328
rect 60884 10288 129096 10316
rect 60884 10276 60890 10288
rect 129090 10276 129096 10288
rect 129148 10276 129154 10328
rect 167086 10276 167092 10328
rect 167144 10316 167150 10328
rect 539686 10316 539692 10328
rect 167144 10288 539692 10316
rect 167144 10276 167150 10288
rect 539686 10276 539692 10288
rect 539744 10276 539750 10328
rect 116394 9256 116400 9308
rect 116452 9296 116458 9308
rect 134702 9296 134708 9308
rect 116452 9268 134708 9296
rect 116452 9256 116458 9268
rect 134702 9256 134708 9268
rect 134760 9256 134766 9308
rect 53742 9188 53748 9240
rect 53800 9228 53806 9240
rect 128630 9228 128636 9240
rect 53800 9200 128636 9228
rect 53800 9188 53806 9200
rect 128630 9188 128636 9200
rect 128688 9188 128694 9240
rect 138382 9188 138388 9240
rect 138440 9228 138446 9240
rect 144914 9228 144920 9240
rect 138440 9200 144920 9228
rect 138440 9188 138446 9200
rect 144914 9188 144920 9200
rect 144972 9188 144978 9240
rect 149054 9188 149060 9240
rect 149112 9228 149118 9240
rect 311434 9228 311440 9240
rect 149112 9200 311440 9228
rect 149112 9188 149118 9200
rect 311434 9188 311440 9200
rect 311492 9188 311498 9240
rect 50154 9120 50160 9172
rect 50212 9160 50218 9172
rect 127618 9160 127624 9172
rect 50212 9132 127624 9160
rect 50212 9120 50218 9132
rect 127618 9120 127624 9132
rect 127676 9120 127682 9172
rect 149146 9120 149152 9172
rect 149204 9160 149210 9172
rect 313826 9160 313832 9172
rect 149204 9132 313832 9160
rect 149204 9120 149210 9132
rect 313826 9120 313832 9132
rect 313884 9120 313890 9172
rect 34790 9052 34796 9104
rect 34848 9092 34854 9104
rect 127342 9092 127348 9104
rect 34848 9064 127348 9092
rect 34848 9052 34854 9064
rect 127342 9052 127348 9064
rect 127400 9052 127406 9104
rect 153286 9052 153292 9104
rect 153344 9092 153350 9104
rect 365806 9092 365812 9104
rect 153344 9064 365812 9092
rect 153344 9052 153350 9064
rect 365806 9052 365812 9064
rect 365864 9052 365870 9104
rect 9950 8984 9956 9036
rect 10008 9024 10014 9036
rect 126054 9024 126060 9036
rect 10008 8996 126060 9024
rect 10008 8984 10014 8996
rect 126054 8984 126060 8996
rect 126112 8984 126118 9036
rect 157426 8984 157432 9036
rect 157484 9024 157490 9036
rect 417878 9024 417884 9036
rect 157484 8996 417884 9024
rect 157484 8984 157490 8996
rect 417878 8984 417884 8996
rect 417936 8984 417942 9036
rect 566 8916 572 8968
rect 624 8956 630 8968
rect 124214 8956 124220 8968
rect 624 8928 124220 8956
rect 624 8916 630 8928
rect 124214 8916 124220 8928
rect 124272 8916 124278 8968
rect 163038 8916 163044 8968
rect 163096 8956 163102 8968
rect 492306 8956 492312 8968
rect 163096 8928 492312 8956
rect 163096 8916 163102 8928
rect 492306 8916 492312 8928
rect 492364 8916 492370 8968
rect 105722 8032 105728 8084
rect 105780 8072 105786 8084
rect 132770 8072 132776 8084
rect 105780 8044 132776 8072
rect 105780 8032 105786 8044
rect 132770 8032 132776 8044
rect 132828 8032 132834 8084
rect 104526 7964 104532 8016
rect 104584 8004 104590 8016
rect 132678 8004 132684 8016
rect 104584 7976 132684 8004
rect 104584 7964 104590 7976
rect 132678 7964 132684 7976
rect 132736 7964 132742 8016
rect 98638 7896 98644 7948
rect 98696 7936 98702 7948
rect 132862 7936 132868 7948
rect 98696 7908 132868 7936
rect 98696 7896 98702 7908
rect 132862 7896 132868 7908
rect 132920 7896 132926 7948
rect 84470 7828 84476 7880
rect 84528 7868 84534 7880
rect 131482 7868 131488 7880
rect 84528 7840 131488 7868
rect 84528 7828 84534 7840
rect 131482 7828 131488 7840
rect 131540 7828 131546 7880
rect 80882 7760 80888 7812
rect 80940 7800 80946 7812
rect 131666 7800 131672 7812
rect 80940 7772 131672 7800
rect 80940 7760 80946 7772
rect 131666 7760 131672 7772
rect 131724 7760 131730 7812
rect 143534 7760 143540 7812
rect 143592 7800 143598 7812
rect 242986 7800 242992 7812
rect 143592 7772 242992 7800
rect 143592 7760 143598 7772
rect 242986 7760 242992 7772
rect 243044 7760 243050 7812
rect 77386 7692 77392 7744
rect 77444 7732 77450 7744
rect 131574 7732 131580 7744
rect 77444 7704 131580 7732
rect 77444 7692 77450 7704
rect 131574 7692 131580 7704
rect 131632 7692 131638 7744
rect 146386 7692 146392 7744
rect 146444 7732 146450 7744
rect 278314 7732 278320 7744
rect 146444 7704 278320 7732
rect 146444 7692 146450 7704
rect 278314 7692 278320 7704
rect 278372 7692 278378 7744
rect 6454 7624 6460 7676
rect 6512 7664 6518 7676
rect 22738 7664 22744 7676
rect 6512 7636 22744 7664
rect 6512 7624 6518 7636
rect 22738 7624 22744 7636
rect 22796 7624 22802 7676
rect 27706 7624 27712 7676
rect 27764 7664 27770 7676
rect 127250 7664 127256 7676
rect 27764 7636 127256 7664
rect 27764 7624 27770 7636
rect 127250 7624 127256 7636
rect 127308 7624 127314 7676
rect 147674 7624 147680 7676
rect 147732 7664 147738 7676
rect 293678 7664 293684 7676
rect 147732 7636 293684 7664
rect 147732 7624 147738 7636
rect 293678 7624 293684 7636
rect 293736 7624 293742 7676
rect 18230 7556 18236 7608
rect 18288 7596 18294 7608
rect 125962 7596 125968 7608
rect 18288 7568 125968 7596
rect 18288 7556 18294 7568
rect 125962 7556 125968 7568
rect 126020 7556 126026 7608
rect 161474 7556 161480 7608
rect 161532 7596 161538 7608
rect 473446 7596 473452 7608
rect 161532 7568 473452 7596
rect 161532 7556 161538 7568
rect 473446 7556 473452 7568
rect 473504 7556 473510 7608
rect 555418 6808 555424 6860
rect 555476 6848 555482 6860
rect 580166 6848 580172 6860
rect 555476 6820 580172 6848
rect 555476 6808 555482 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 140774 6604 140780 6656
rect 140832 6644 140838 6656
rect 203886 6644 203892 6656
rect 140832 6616 203892 6644
rect 140832 6604 140838 6616
rect 203886 6604 203892 6616
rect 203944 6604 203950 6656
rect 142154 6536 142160 6588
rect 142212 6576 142218 6588
rect 225138 6576 225144 6588
rect 142212 6548 225144 6576
rect 142212 6536 142218 6548
rect 225138 6536 225144 6548
rect 225196 6536 225202 6588
rect 66714 6468 66720 6520
rect 66772 6508 66778 6520
rect 130102 6508 130108 6520
rect 66772 6480 130108 6508
rect 66772 6468 66778 6480
rect 130102 6468 130108 6480
rect 130160 6468 130166 6520
rect 146294 6468 146300 6520
rect 146352 6508 146358 6520
rect 276014 6508 276020 6520
rect 146352 6480 276020 6508
rect 146352 6468 146358 6480
rect 276014 6468 276020 6480
rect 276072 6468 276078 6520
rect 391198 6468 391204 6520
rect 391256 6508 391262 6520
rect 582190 6508 582196 6520
rect 391256 6480 582196 6508
rect 391256 6468 391262 6480
rect 582190 6468 582196 6480
rect 582248 6468 582254 6520
rect 63218 6400 63224 6452
rect 63276 6440 63282 6452
rect 130010 6440 130016 6452
rect 63276 6412 130016 6440
rect 63276 6400 63282 6412
rect 130010 6400 130016 6412
rect 130068 6400 130074 6452
rect 155954 6400 155960 6452
rect 156012 6440 156018 6452
rect 394234 6440 394240 6452
rect 156012 6412 394240 6440
rect 156012 6400 156018 6412
rect 394234 6400 394240 6412
rect 394292 6400 394298 6452
rect 48958 6332 48964 6384
rect 49016 6372 49022 6384
rect 128538 6372 128544 6384
rect 49016 6344 128544 6372
rect 49016 6332 49022 6344
rect 128538 6332 128544 6344
rect 128596 6332 128602 6384
rect 156046 6332 156052 6384
rect 156104 6372 156110 6384
rect 400122 6372 400128 6384
rect 156104 6344 400128 6372
rect 156104 6332 156110 6344
rect 400122 6332 400128 6344
rect 400180 6332 400186 6384
rect 44266 6264 44272 6316
rect 44324 6304 44330 6316
rect 129274 6304 129280 6316
rect 44324 6276 129280 6304
rect 44324 6264 44330 6276
rect 129274 6264 129280 6276
rect 129332 6264 129338 6316
rect 160094 6264 160100 6316
rect 160152 6304 160158 6316
rect 446214 6304 446220 6316
rect 160152 6276 446220 6304
rect 160152 6264 160158 6276
rect 446214 6264 446220 6276
rect 446272 6264 446278 6316
rect 33594 6196 33600 6248
rect 33652 6236 33658 6248
rect 127158 6236 127164 6248
rect 33652 6208 127164 6236
rect 33652 6196 33658 6208
rect 127158 6196 127164 6208
rect 127216 6196 127222 6248
rect 162946 6196 162952 6248
rect 163004 6236 163010 6248
rect 493502 6236 493508 6248
rect 163004 6208 493508 6236
rect 163004 6196 163010 6208
rect 493502 6196 493508 6208
rect 493560 6196 493566 6248
rect 24210 6128 24216 6180
rect 24268 6168 24274 6180
rect 122098 6168 122104 6180
rect 24268 6140 122104 6168
rect 24268 6128 24274 6140
rect 122098 6128 122104 6140
rect 122156 6128 122162 6180
rect 168374 6128 168380 6180
rect 168432 6168 168438 6180
rect 562042 6168 562048 6180
rect 168432 6140 562048 6168
rect 168432 6128 168438 6140
rect 562042 6128 562048 6140
rect 562100 6128 562106 6180
rect 101030 5380 101036 5432
rect 101088 5420 101094 5432
rect 133138 5420 133144 5432
rect 101088 5392 133144 5420
rect 101088 5380 101094 5392
rect 133138 5380 133144 5392
rect 133196 5380 133202 5432
rect 97442 5312 97448 5364
rect 97500 5352 97506 5364
rect 133322 5352 133328 5364
rect 97500 5324 133328 5352
rect 97500 5312 97506 5324
rect 133322 5312 133328 5324
rect 133380 5312 133386 5364
rect 136726 5312 136732 5364
rect 136784 5352 136790 5364
rect 150618 5352 150624 5364
rect 136784 5324 150624 5352
rect 136784 5312 136790 5324
rect 150618 5312 150624 5324
rect 150676 5312 150682 5364
rect 85666 5244 85672 5296
rect 85724 5284 85730 5296
rect 131390 5284 131396 5296
rect 85724 5256 131396 5284
rect 85724 5244 85730 5256
rect 131390 5244 131396 5256
rect 131448 5244 131454 5296
rect 138290 5244 138296 5296
rect 138348 5284 138354 5296
rect 171962 5284 171968 5296
rect 138348 5256 171968 5284
rect 138348 5244 138354 5256
rect 171962 5244 171968 5256
rect 172020 5244 172026 5296
rect 15930 5176 15936 5228
rect 15988 5216 15994 5228
rect 46198 5216 46204 5228
rect 15988 5188 46204 5216
rect 15988 5176 15994 5188
rect 46198 5176 46204 5188
rect 46256 5176 46262 5228
rect 59630 5176 59636 5228
rect 59688 5216 59694 5228
rect 129918 5216 129924 5228
rect 59688 5188 129924 5216
rect 59688 5176 59694 5188
rect 129918 5176 129924 5188
rect 129976 5176 129982 5228
rect 151538 5176 151544 5228
rect 151596 5216 151602 5228
rect 329190 5216 329196 5228
rect 151596 5188 329196 5216
rect 151596 5176 151602 5188
rect 329190 5176 329196 5188
rect 329248 5176 329254 5228
rect 30098 5108 30104 5160
rect 30156 5148 30162 5160
rect 127526 5148 127532 5160
rect 30156 5120 127532 5148
rect 30156 5108 30162 5120
rect 127526 5108 127532 5120
rect 127584 5108 127590 5160
rect 136910 5108 136916 5160
rect 136968 5148 136974 5160
rect 148318 5148 148324 5160
rect 136968 5120 148324 5148
rect 136968 5108 136974 5120
rect 148318 5108 148324 5120
rect 148376 5108 148382 5160
rect 153194 5108 153200 5160
rect 153252 5148 153258 5160
rect 358722 5148 358728 5160
rect 153252 5120 358728 5148
rect 153252 5108 153258 5120
rect 358722 5108 358728 5120
rect 358780 5108 358786 5160
rect 28902 5040 28908 5092
rect 28960 5080 28966 5092
rect 127802 5080 127808 5092
rect 28960 5052 127808 5080
rect 28960 5040 28966 5052
rect 127802 5040 127808 5052
rect 127860 5040 127866 5092
rect 137002 5040 137008 5092
rect 137060 5080 137066 5092
rect 151814 5080 151820 5092
rect 137060 5052 151820 5080
rect 137060 5040 137066 5052
rect 151814 5040 151820 5052
rect 151872 5040 151878 5092
rect 157334 5040 157340 5092
rect 157392 5080 157398 5092
rect 414290 5080 414296 5092
rect 157392 5052 414296 5080
rect 157392 5040 157398 5052
rect 414290 5040 414296 5052
rect 414348 5040 414354 5092
rect 19426 4972 19432 5024
rect 19484 5012 19490 5024
rect 124858 5012 124864 5024
rect 19484 4984 124864 5012
rect 19484 4972 19490 4984
rect 124858 4972 124864 4984
rect 124916 4972 124922 5024
rect 138106 4972 138112 5024
rect 138164 5012 138170 5024
rect 167178 5012 167184 5024
rect 138164 4984 167184 5012
rect 138164 4972 138170 4984
rect 167178 4972 167184 4984
rect 167236 4972 167242 5024
rect 170674 4972 170680 5024
rect 170732 5012 170738 5024
rect 480530 5012 480536 5024
rect 170732 4984 480536 5012
rect 170732 4972 170738 4984
rect 480530 4972 480536 4984
rect 480588 4972 480594 5024
rect 13538 4904 13544 4956
rect 13596 4944 13602 4956
rect 126514 4944 126520 4956
rect 13596 4916 126520 4944
rect 13596 4904 13602 4916
rect 126514 4904 126520 4916
rect 126572 4904 126578 4956
rect 137094 4904 137100 4956
rect 137152 4944 137158 4956
rect 154206 4944 154212 4956
rect 137152 4916 154212 4944
rect 137152 4904 137158 4916
rect 154206 4904 154212 4916
rect 154264 4904 154270 4956
rect 162854 4904 162860 4956
rect 162912 4944 162918 4956
rect 491110 4944 491116 4956
rect 162912 4916 491116 4944
rect 162912 4904 162918 4916
rect 491110 4904 491116 4916
rect 491168 4904 491174 4956
rect 11146 4836 11152 4888
rect 11204 4876 11210 4888
rect 125870 4876 125876 4888
rect 11204 4848 125876 4876
rect 11204 4836 11210 4848
rect 125870 4836 125876 4848
rect 125928 4836 125934 4888
rect 157794 4876 157800 4888
rect 137986 4848 157800 4876
rect 8754 4768 8760 4820
rect 8812 4808 8818 4820
rect 125778 4808 125784 4820
rect 8812 4780 125784 4808
rect 8812 4768 8818 4780
rect 125778 4768 125784 4780
rect 125836 4768 125842 4820
rect 136818 4700 136824 4752
rect 136876 4740 136882 4752
rect 137986 4740 138014 4848
rect 157794 4836 157800 4848
rect 157852 4836 157858 4888
rect 168190 4836 168196 4888
rect 168248 4876 168254 4888
rect 545482 4876 545488 4888
rect 168248 4848 545488 4876
rect 168248 4836 168254 4848
rect 545482 4836 545488 4848
rect 545540 4836 545546 4888
rect 138198 4768 138204 4820
rect 138256 4808 138262 4820
rect 162486 4808 162492 4820
rect 138256 4780 162492 4808
rect 138256 4768 138262 4780
rect 162486 4768 162492 4780
rect 162544 4768 162550 4820
rect 169754 4768 169760 4820
rect 169812 4808 169818 4820
rect 576302 4808 576308 4820
rect 169812 4780 576308 4808
rect 169812 4768 169818 4780
rect 576302 4768 576308 4780
rect 576360 4768 576366 4820
rect 136876 4712 138014 4740
rect 136876 4700 136882 4712
rect 135990 4156 135996 4208
rect 136048 4196 136054 4208
rect 141234 4196 141240 4208
rect 136048 4168 141240 4196
rect 136048 4156 136054 4168
rect 141234 4156 141240 4168
rect 141292 4156 141298 4208
rect 119890 4088 119896 4140
rect 119948 4128 119954 4140
rect 124950 4128 124956 4140
rect 119948 4100 124956 4128
rect 119948 4088 119954 4100
rect 124950 4088 124956 4100
rect 125008 4088 125014 4140
rect 125870 4088 125876 4140
rect 125928 4128 125934 4140
rect 134518 4128 134524 4140
rect 125928 4100 134524 4128
rect 125928 4088 125934 4100
rect 134518 4088 134524 4100
rect 134576 4088 134582 4140
rect 137738 4088 137744 4140
rect 137796 4128 137802 4140
rect 144730 4128 144736 4140
rect 137796 4100 144736 4128
rect 137796 4088 137802 4100
rect 144730 4088 144736 4100
rect 144788 4088 144794 4140
rect 138934 4020 138940 4072
rect 138992 4060 138998 4072
rect 143534 4060 143540 4072
rect 138992 4032 143540 4060
rect 138992 4020 138998 4032
rect 143534 4020 143540 4032
rect 143592 4020 143598 4072
rect 12342 3952 12348 4004
rect 12400 3992 12406 4004
rect 126422 3992 126428 4004
rect 12400 3964 126428 3992
rect 12400 3952 12406 3964
rect 126422 3952 126428 3964
rect 126480 3952 126486 4004
rect 138658 3952 138664 4004
rect 138716 3992 138722 4004
rect 145926 3992 145932 4004
rect 138716 3964 145932 3992
rect 138716 3952 138722 3964
rect 145926 3952 145932 3964
rect 145984 3952 145990 4004
rect 144454 3884 144460 3936
rect 144512 3924 144518 3936
rect 153010 3924 153016 3936
rect 144512 3896 153016 3924
rect 144512 3884 144518 3896
rect 153010 3884 153016 3896
rect 153068 3884 153074 3936
rect 86862 3816 86868 3868
rect 86920 3856 86926 3868
rect 131850 3856 131856 3868
rect 86920 3828 131856 3856
rect 86920 3816 86926 3828
rect 131850 3816 131856 3828
rect 131908 3816 131914 3868
rect 135714 3816 135720 3868
rect 135772 3856 135778 3868
rect 140038 3856 140044 3868
rect 135772 3828 140044 3856
rect 135772 3816 135778 3828
rect 140038 3816 140044 3828
rect 140096 3816 140102 3868
rect 140130 3816 140136 3868
rect 140188 3856 140194 3868
rect 149514 3856 149520 3868
rect 140188 3828 149520 3856
rect 140188 3816 140194 3828
rect 149514 3816 149520 3828
rect 149572 3816 149578 3868
rect 211798 3816 211804 3868
rect 211856 3856 211862 3868
rect 211856 3828 219434 3856
rect 211856 3816 211862 3828
rect 83274 3748 83280 3800
rect 83332 3788 83338 3800
rect 83332 3760 131436 3788
rect 83332 3748 83338 3760
rect 79686 3680 79692 3732
rect 79744 3720 79750 3732
rect 131298 3720 131304 3732
rect 79744 3692 131304 3720
rect 79744 3680 79750 3692
rect 131298 3680 131304 3692
rect 131356 3680 131362 3732
rect 131408 3720 131436 3760
rect 131758 3748 131764 3800
rect 131816 3788 131822 3800
rect 135806 3788 135812 3800
rect 131816 3760 135812 3788
rect 131816 3748 131822 3760
rect 135806 3748 135812 3760
rect 135864 3748 135870 3800
rect 142982 3748 142988 3800
rect 143040 3788 143046 3800
rect 155402 3788 155408 3800
rect 143040 3760 155408 3788
rect 143040 3748 143046 3760
rect 155402 3748 155408 3760
rect 155460 3748 155466 3800
rect 172054 3748 172060 3800
rect 172112 3788 172118 3800
rect 212166 3788 212172 3800
rect 172112 3760 212172 3788
rect 172112 3748 172118 3760
rect 212166 3748 212172 3760
rect 212224 3748 212230 3800
rect 219406 3788 219434 3828
rect 242894 3816 242900 3868
rect 242952 3856 242958 3868
rect 244090 3856 244096 3868
rect 242952 3828 244096 3856
rect 242952 3816 242958 3828
rect 244090 3816 244096 3828
rect 244148 3816 244154 3868
rect 251174 3816 251180 3868
rect 251232 3856 251238 3868
rect 252370 3856 252376 3868
rect 251232 3828 252376 3856
rect 251232 3816 251238 3828
rect 252370 3816 252376 3828
rect 252428 3816 252434 3868
rect 284294 3816 284300 3868
rect 284352 3856 284358 3868
rect 285030 3856 285036 3868
rect 284352 3828 285036 3856
rect 284352 3816 284358 3828
rect 285030 3816 285036 3828
rect 285088 3816 285094 3868
rect 344554 3788 344560 3800
rect 219406 3760 344560 3788
rect 344554 3748 344560 3760
rect 344612 3748 344618 3800
rect 132034 3720 132040 3732
rect 131408 3692 132040 3720
rect 132034 3680 132040 3692
rect 132092 3680 132098 3732
rect 135438 3680 135444 3732
rect 135496 3720 135502 3732
rect 137646 3720 137652 3732
rect 135496 3692 137652 3720
rect 135496 3680 135502 3692
rect 137646 3680 137652 3692
rect 137704 3680 137710 3732
rect 144914 3680 144920 3732
rect 144972 3720 144978 3732
rect 144972 3692 147674 3720
rect 144972 3680 144978 3692
rect 72602 3612 72608 3664
rect 72660 3652 72666 3664
rect 126238 3652 126244 3664
rect 72660 3624 126244 3652
rect 72660 3612 72666 3624
rect 126238 3612 126244 3624
rect 126296 3612 126302 3664
rect 130654 3652 130660 3664
rect 126716 3624 130660 3652
rect 69106 3544 69112 3596
rect 69164 3584 69170 3596
rect 126716 3584 126744 3624
rect 130654 3612 130660 3624
rect 130712 3612 130718 3664
rect 132954 3612 132960 3664
rect 133012 3652 133018 3664
rect 135530 3652 135536 3664
rect 133012 3624 135536 3652
rect 133012 3612 133018 3624
rect 135530 3612 135536 3624
rect 135588 3612 135594 3664
rect 135622 3612 135628 3664
rect 135680 3652 135686 3664
rect 138842 3652 138848 3664
rect 135680 3624 138848 3652
rect 135680 3612 135686 3624
rect 138842 3612 138848 3624
rect 138900 3612 138906 3664
rect 139946 3612 139952 3664
rect 140004 3652 140010 3664
rect 147646 3652 147674 3692
rect 149974 3680 149980 3732
rect 150032 3720 150038 3732
rect 163682 3720 163688 3732
rect 150032 3692 163688 3720
rect 150032 3680 150038 3692
rect 163682 3680 163688 3692
rect 163740 3680 163746 3732
rect 171778 3680 171784 3732
rect 171836 3720 171842 3732
rect 445018 3720 445024 3732
rect 171836 3692 445024 3720
rect 171836 3680 171842 3692
rect 445018 3680 445024 3692
rect 445076 3680 445082 3732
rect 169570 3652 169576 3664
rect 140004 3624 147352 3652
rect 147646 3624 169576 3652
rect 140004 3612 140010 3624
rect 69164 3556 126744 3584
rect 69164 3544 69170 3556
rect 126974 3544 126980 3596
rect 127032 3584 127038 3596
rect 130378 3584 130384 3596
rect 127032 3556 130384 3584
rect 127032 3544 127038 3556
rect 130378 3544 130384 3556
rect 130436 3544 130442 3596
rect 135346 3544 135352 3596
rect 135404 3584 135410 3596
rect 136450 3584 136456 3596
rect 135404 3556 136456 3584
rect 135404 3544 135410 3556
rect 136450 3544 136456 3556
rect 136508 3544 136514 3596
rect 142798 3544 142804 3596
rect 142856 3584 142862 3596
rect 147324 3584 147352 3624
rect 169570 3612 169576 3624
rect 169628 3612 169634 3664
rect 171870 3612 171876 3664
rect 171928 3652 171934 3664
rect 465166 3652 465172 3664
rect 171928 3624 465172 3652
rect 171928 3612 171934 3624
rect 465166 3612 465172 3624
rect 465224 3612 465230 3664
rect 166074 3584 166080 3596
rect 142856 3556 147260 3584
rect 147324 3556 166080 3584
rect 142856 3544 142862 3556
rect 23014 3476 23020 3528
rect 23072 3516 23078 3528
rect 88150 3516 88156 3528
rect 23072 3488 88156 3516
rect 23072 3476 23078 3488
rect 88150 3476 88156 3488
rect 88208 3476 88214 3528
rect 93854 3476 93860 3528
rect 93912 3516 93918 3528
rect 94774 3516 94780 3528
rect 93912 3488 94780 3516
rect 93912 3476 93918 3488
rect 94774 3476 94780 3488
rect 94832 3476 94838 3528
rect 110414 3476 110420 3528
rect 110472 3516 110478 3528
rect 111610 3516 111616 3528
rect 110472 3488 111616 3516
rect 110472 3476 110478 3488
rect 111610 3476 111616 3488
rect 111668 3476 111674 3528
rect 124674 3476 124680 3528
rect 124732 3516 124738 3528
rect 134610 3516 134616 3528
rect 124732 3488 134616 3516
rect 124732 3476 124738 3488
rect 134610 3476 134616 3488
rect 134668 3476 134674 3528
rect 135162 3476 135168 3528
rect 135220 3516 135226 3528
rect 147122 3516 147128 3528
rect 135220 3488 147128 3516
rect 135220 3476 135226 3488
rect 147122 3476 147128 3488
rect 147180 3476 147186 3528
rect 147232 3516 147260 3556
rect 166074 3544 166080 3556
rect 166132 3544 166138 3596
rect 172146 3544 172152 3596
rect 172204 3584 172210 3596
rect 468662 3584 468668 3596
rect 172204 3556 468668 3584
rect 172204 3544 172210 3556
rect 468662 3544 468668 3556
rect 468720 3544 468726 3596
rect 475746 3584 475752 3596
rect 470566 3556 475752 3584
rect 147232 3488 163636 3516
rect 35894 3408 35900 3460
rect 35952 3448 35958 3460
rect 36814 3448 36820 3460
rect 35952 3420 36820 3448
rect 35952 3408 35958 3420
rect 36814 3408 36820 3420
rect 36872 3408 36878 3460
rect 60734 3408 60740 3460
rect 60792 3448 60798 3460
rect 61654 3448 61660 3460
rect 60792 3420 61660 3448
rect 60792 3408 60798 3420
rect 61654 3408 61660 3420
rect 61712 3408 61718 3460
rect 139026 3408 139032 3460
rect 139084 3448 139090 3460
rect 139084 3420 161474 3448
rect 139084 3408 139090 3420
rect 161446 3312 161474 3420
rect 163608 3380 163636 3488
rect 163774 3476 163780 3528
rect 163832 3516 163838 3528
rect 164878 3516 164884 3528
rect 163832 3488 164884 3516
rect 163832 3476 163838 3488
rect 164878 3476 164884 3488
rect 164936 3476 164942 3528
rect 172238 3476 172244 3528
rect 172296 3516 172302 3528
rect 470566 3516 470594 3556
rect 475746 3544 475752 3556
rect 475804 3544 475810 3596
rect 172296 3488 470594 3516
rect 172296 3476 172302 3488
rect 471238 3476 471244 3528
rect 471296 3516 471302 3528
rect 472250 3516 472256 3528
rect 471296 3488 472256 3516
rect 471296 3476 471302 3488
rect 472250 3476 472256 3488
rect 472308 3476 472314 3528
rect 506474 3476 506480 3528
rect 506532 3516 506538 3528
rect 507302 3516 507308 3528
rect 506532 3488 507308 3516
rect 506532 3476 506538 3488
rect 507302 3476 507308 3488
rect 507360 3476 507366 3528
rect 539594 3476 539600 3528
rect 539652 3516 539658 3528
rect 540422 3516 540428 3528
rect 539652 3488 540428 3516
rect 539652 3476 539658 3488
rect 540422 3476 540428 3488
rect 540480 3476 540486 3528
rect 173250 3408 173256 3460
rect 173308 3448 173314 3460
rect 512454 3448 512460 3460
rect 173308 3420 512460 3448
rect 173308 3408 173314 3420
rect 512454 3408 512460 3420
rect 512512 3408 512518 3460
rect 170766 3380 170772 3392
rect 163608 3352 170772 3380
rect 170766 3340 170772 3352
rect 170824 3340 170830 3392
rect 307754 3340 307760 3392
rect 307812 3380 307818 3392
rect 309042 3380 309048 3392
rect 307812 3352 309048 3380
rect 307812 3340 307818 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 316034 3340 316040 3392
rect 316092 3380 316098 3392
rect 317322 3380 317328 3392
rect 316092 3352 317328 3380
rect 316092 3340 316098 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 324406 3340 324412 3392
rect 324464 3380 324470 3392
rect 325602 3380 325608 3392
rect 324464 3352 325608 3380
rect 324464 3340 324470 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 340966 3340 340972 3392
rect 341024 3380 341030 3392
rect 342162 3380 342168 3392
rect 341024 3352 342168 3380
rect 341024 3340 341030 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 365714 3340 365720 3392
rect 365772 3380 365778 3392
rect 367002 3380 367008 3392
rect 365772 3352 367008 3380
rect 365772 3340 365778 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382366 3340 382372 3392
rect 382424 3380 382430 3392
rect 383562 3380 383568 3392
rect 382424 3352 383568 3380
rect 382424 3340 382430 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 390646 3340 390652 3392
rect 390704 3380 390710 3392
rect 391842 3380 391848 3392
rect 390704 3352 391848 3380
rect 390704 3340 390710 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 407114 3340 407120 3392
rect 407172 3380 407178 3392
rect 408402 3380 408408 3392
rect 407172 3352 408408 3380
rect 407172 3340 407178 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 415394 3340 415400 3392
rect 415452 3380 415458 3392
rect 416682 3380 416688 3392
rect 415452 3352 416688 3380
rect 415452 3340 415458 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 432046 3340 432052 3392
rect 432104 3380 432110 3392
rect 433242 3380 433248 3392
rect 432104 3352 433248 3380
rect 432104 3340 432110 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 440326 3340 440332 3392
rect 440384 3380 440390 3392
rect 441522 3380 441528 3392
rect 440384 3352 441528 3380
rect 440384 3340 440390 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 456794 3340 456800 3392
rect 456852 3380 456858 3392
rect 458082 3380 458088 3392
rect 456852 3352 458088 3380
rect 456852 3340 456858 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 168374 3312 168380 3324
rect 161446 3284 168380 3312
rect 168374 3272 168380 3284
rect 168432 3272 168438 3324
rect 152826 3136 152832 3188
rect 152884 3176 152890 3188
rect 156598 3176 156604 3188
rect 152884 3148 156604 3176
rect 152884 3136 152890 3148
rect 156598 3136 156604 3148
rect 156656 3136 156662 3188
rect 478138 3136 478144 3188
rect 478196 3176 478202 3188
rect 479334 3176 479340 3188
rect 478196 3148 479340 3176
rect 478196 3136 478202 3148
rect 479334 3136 479340 3148
rect 479392 3136 479398 3188
rect 173158 3068 173164 3120
rect 173216 3108 173222 3120
rect 179046 3108 179052 3120
rect 173216 3080 179052 3108
rect 173216 3068 173222 3080
rect 179046 3068 179052 3080
rect 179104 3068 179110 3120
rect 349154 1368 349160 1420
rect 349212 1408 349218 1420
rect 350442 1408 350448 1420
rect 349212 1380 350448 1408
rect 349212 1368 349218 1380
rect 350442 1368 350448 1380
rect 350500 1368 350506 1420
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 410524 700476 410576 700528
rect 429844 700476 429896 700528
rect 399484 700408 399536 700460
rect 446128 700408 446180 700460
rect 409144 700340 409196 700392
rect 494796 700340 494848 700392
rect 24308 700272 24360 700324
rect 33784 700272 33836 700324
rect 407764 700272 407816 700324
rect 559656 700272 559708 700324
rect 196624 699660 196676 699712
rect 202788 699660 202840 699712
rect 229744 699660 229796 699712
rect 235172 699660 235224 699712
rect 364984 699660 365036 699712
rect 369124 699660 369176 699712
rect 300124 697688 300176 697740
rect 307024 697688 307076 697740
rect 260104 697280 260156 697332
rect 267648 697280 267700 697332
rect 152832 696940 152884 696992
rect 154120 696940 154172 696992
rect 504364 696940 504416 696992
rect 580172 696940 580224 696992
rect 150440 692792 150492 692844
rect 152832 692792 152884 692844
rect 185584 692044 185636 692096
rect 196624 692044 196676 692096
rect 210424 690616 210476 690668
rect 229744 690616 229796 690668
rect 180064 689256 180116 689308
rect 185584 689256 185636 689308
rect 369124 688576 369176 688628
rect 374644 688576 374696 688628
rect 347780 688440 347832 688492
rect 351920 688440 351972 688492
rect 146944 687148 146996 687200
rect 150348 687216 150400 687268
rect 307024 684428 307076 684480
rect 310244 684428 310296 684480
rect 351920 683748 351972 683800
rect 362224 683748 362276 683800
rect 374644 682252 374696 682304
rect 380256 682252 380308 682304
rect 362224 680960 362276 681012
rect 371240 680960 371292 681012
rect 217324 680348 217376 680400
rect 218060 680348 218112 680400
rect 310244 678716 310296 678768
rect 315304 678716 315356 678768
rect 253572 678444 253624 678496
rect 260104 678444 260156 678496
rect 144920 678240 144972 678292
rect 146944 678240 146996 678292
rect 135996 676812 136048 676864
rect 144920 676812 144972 676864
rect 371240 675452 371292 675504
rect 380164 675452 380216 675504
rect 380256 675452 380308 675504
rect 396448 675452 396500 675504
rect 278412 674772 278464 674824
rect 282828 674772 282880 674824
rect 331220 674772 331272 674824
rect 334624 674772 334676 674824
rect 133880 674432 133932 674484
rect 135996 674432 136048 674484
rect 250444 674024 250496 674076
rect 253572 674024 253624 674076
rect 2780 670692 2832 670744
rect 6184 670692 6236 670744
rect 544384 670692 544436 670744
rect 580172 670692 580224 670744
rect 276664 669060 276716 669112
rect 278412 669060 278464 669112
rect 131764 667496 131816 667548
rect 133880 667496 133932 667548
rect 202144 667156 202196 667208
rect 210424 667156 210476 667208
rect 177304 666408 177356 666460
rect 180064 666408 180116 666460
rect 247684 663756 247736 663808
rect 250444 663756 250496 663808
rect 334624 663008 334676 663060
rect 358084 663008 358136 663060
rect 127624 662396 127676 662448
rect 131764 662396 131816 662448
rect 174544 662396 174596 662448
rect 177304 662396 177356 662448
rect 273904 661036 273956 661088
rect 276664 661036 276716 661088
rect 214564 658792 214616 658844
rect 217324 658792 217376 658844
rect 315304 653352 315356 653404
rect 319812 653352 319864 653404
rect 171692 651380 171744 651432
rect 174544 651380 174596 651432
rect 195244 650700 195296 650752
rect 202144 650700 202196 650752
rect 269764 649952 269816 650004
rect 273904 650020 273956 650072
rect 358084 649952 358136 650004
rect 366364 649952 366416 650004
rect 163504 649272 163556 649324
rect 171692 649272 171744 649324
rect 380164 649272 380216 649324
rect 387064 649272 387116 649324
rect 319812 648864 319864 648916
rect 324964 648864 325016 648916
rect 124864 648524 124916 648576
rect 127624 648592 127676 648644
rect 265624 647912 265676 647964
rect 269764 647912 269816 647964
rect 366364 647164 366416 647216
rect 371884 647164 371936 647216
rect 244924 645804 244976 645856
rect 247684 645804 247736 645856
rect 324964 640228 325016 640280
rect 327724 640228 327776 640280
rect 156604 638460 156656 638512
rect 163504 638460 163556 638512
rect 371884 635468 371936 635520
rect 388904 635468 388956 635520
rect 327724 632476 327776 632528
rect 329932 632476 329984 632528
rect 388904 631660 388956 631712
rect 395344 631660 395396 631712
rect 329932 629892 329984 629944
rect 339500 629892 339552 629944
rect 339500 626492 339552 626544
rect 344008 626492 344060 626544
rect 186964 623024 187016 623076
rect 195244 623024 195296 623076
rect 152464 622412 152516 622464
rect 156604 622412 156656 622464
rect 344008 620236 344060 620288
rect 353300 620236 353352 620288
rect 3516 618264 3568 618316
rect 15844 618264 15896 618316
rect 353300 617516 353352 617568
rect 395436 617516 395488 617568
rect 406384 616836 406436 616888
rect 579712 616836 579764 616888
rect 184204 612756 184256 612808
rect 186964 612756 187016 612808
rect 211804 609696 211856 609748
rect 214564 609696 214616 609748
rect 138664 603712 138716 603764
rect 152464 603712 152516 603764
rect 178040 603712 178092 603764
rect 184204 603712 184256 603764
rect 121460 603032 121512 603084
rect 124864 603100 124916 603152
rect 171784 600312 171836 600364
rect 178040 600312 178092 600364
rect 119988 599564 120040 599616
rect 121460 599564 121512 599616
rect 263600 598748 263652 598800
rect 265624 598748 265676 598800
rect 117688 597184 117740 597236
rect 119988 597184 120040 597236
rect 249064 595416 249116 595468
rect 263600 595416 263652 595468
rect 210424 592016 210476 592068
rect 211804 592016 211856 592068
rect 115204 590588 115256 590640
rect 117688 590588 117740 590640
rect 241612 581136 241664 581188
rect 244924 581136 244976 581188
rect 112444 580932 112496 580984
rect 115204 580932 115256 580984
rect 135904 580660 135956 580712
rect 138664 580660 138716 580712
rect 157984 580252 158036 580304
rect 171784 580252 171836 580304
rect 3332 579640 3384 579692
rect 19984 579640 20036 579692
rect 238760 577600 238812 577652
rect 241612 577600 241664 577652
rect 236644 574064 236696 574116
rect 238760 574064 238812 574116
rect 126244 571956 126296 572008
rect 135904 571956 135956 572008
rect 3056 565836 3108 565888
rect 43444 565836 43496 565888
rect 405004 563048 405056 563100
rect 580172 563048 580224 563100
rect 233240 562096 233292 562148
rect 236644 562096 236696 562148
rect 209044 558152 209096 558204
rect 233240 558152 233292 558204
rect 207664 554412 207716 554464
rect 210424 554412 210476 554464
rect 149704 545708 149756 545760
rect 157984 545708 158036 545760
rect 206284 543736 206336 543788
rect 207664 543736 207716 543788
rect 204904 536800 204956 536852
rect 209044 536800 209096 536852
rect 2964 527144 3016 527196
rect 20076 527144 20128 527196
rect 108948 525716 109000 525768
rect 112444 525784 112496 525836
rect 123484 525784 123536 525836
rect 126244 525784 126296 525836
rect 106924 522520 106976 522572
rect 108948 522520 109000 522572
rect 2780 514768 2832 514820
rect 4804 514768 4856 514820
rect 105544 514768 105596 514820
rect 106924 514768 106976 514820
rect 115204 514020 115256 514072
rect 123484 514020 123536 514072
rect 203524 511912 203576 511964
rect 206284 511912 206336 511964
rect 403624 510620 403676 510672
rect 580172 510620 580224 510672
rect 201868 507832 201920 507884
rect 204904 507832 204956 507884
rect 88984 504364 89036 504416
rect 115204 504364 115256 504416
rect 189724 500216 189776 500268
rect 201868 500216 201920 500268
rect 236644 497428 236696 497480
rect 249064 497428 249116 497480
rect 138020 496068 138072 496120
rect 149704 496068 149756 496120
rect 80704 491920 80756 491972
rect 88984 491920 89036 491972
rect 128544 490560 128596 490612
rect 138020 490560 138072 490612
rect 125692 487500 125744 487552
rect 128544 487500 128596 487552
rect 120724 485052 120776 485104
rect 125692 485052 125744 485104
rect 77944 478864 77996 478916
rect 80704 478864 80756 478916
rect 235264 474648 235316 474700
rect 236644 474648 236696 474700
rect 232504 466420 232556 466472
rect 235264 466420 235316 466472
rect 115572 466080 115624 466132
rect 120724 466080 120776 466132
rect 3240 462544 3292 462596
rect 8944 462544 8996 462596
rect 109684 462340 109736 462392
rect 115572 462340 115624 462392
rect 64144 457444 64196 457496
rect 77944 457444 77996 457496
rect 400864 456764 400916 456816
rect 580172 456764 580224 456816
rect 226432 446360 226484 446412
rect 232504 446360 232556 446412
rect 201592 445816 201644 445868
rect 203524 445816 203576 445868
rect 199384 445340 199436 445392
rect 201592 445340 201644 445392
rect 48412 445000 48464 445052
rect 64144 445000 64196 445052
rect 104164 442892 104216 442944
rect 105544 442892 105596 442944
rect 225604 442416 225656 442468
rect 226432 442416 226484 442468
rect 46664 442280 46716 442332
rect 48412 442280 48464 442332
rect 184204 438880 184256 438932
rect 189724 438880 189776 438932
rect 196624 437384 196676 437436
rect 199384 437452 199436 437504
rect 45008 436840 45060 436892
rect 46664 436840 46716 436892
rect 174544 435344 174596 435396
rect 184204 435344 184256 435396
rect 396724 430584 396776 430636
rect 579988 430584 580040 430636
rect 169024 429836 169076 429888
rect 174544 429836 174596 429888
rect 193864 426844 193916 426896
rect 196624 426844 196676 426896
rect 106924 423580 106976 423632
rect 109684 423580 109736 423632
rect 3148 422900 3200 422952
rect 6276 422900 6328 422952
rect 3148 409844 3200 409896
rect 10324 409844 10376 409896
rect 166264 407532 166316 407584
rect 169024 407532 169076 407584
rect 224224 407328 224276 407380
rect 225604 407328 225656 407380
rect 191104 404268 191156 404320
rect 193864 404336 193916 404388
rect 418804 404336 418856 404388
rect 580080 404336 580132 404388
rect 69664 396720 69716 396772
rect 136640 396720 136692 396772
rect 223028 395972 223080 396024
rect 224224 395972 224276 396024
rect 95884 392572 95936 392624
rect 106924 392572 106976 392624
rect 163504 391960 163556 392012
rect 166264 391960 166316 392012
rect 209044 387064 209096 387116
rect 223028 387064 223080 387116
rect 68284 384956 68336 385008
rect 69664 384956 69716 385008
rect 186964 384956 187016 385008
rect 191104 385024 191156 385076
rect 78588 382916 78640 382968
rect 95884 382916 95936 382968
rect 205640 382236 205692 382288
rect 209044 382236 209096 382288
rect 102784 381488 102836 381540
rect 163504 381488 163556 381540
rect 64236 380128 64288 380180
rect 78588 380128 78640 380180
rect 102140 379176 102192 379228
rect 104164 379176 104216 379228
rect 396816 378156 396868 378208
rect 580080 378156 580132 378208
rect 202144 378088 202196 378140
rect 205640 378088 205692 378140
rect 101404 374960 101456 375012
rect 102140 374960 102192 375012
rect 198004 372512 198056 372564
rect 202144 372580 202196 372632
rect 3240 371220 3292 371272
rect 24124 371220 24176 371272
rect 95884 369860 95936 369912
rect 102784 369860 102836 369912
rect 398104 364352 398156 364404
rect 579804 364352 579856 364404
rect 100024 362924 100076 362976
rect 101404 362924 101456 362976
rect 65432 358776 65484 358828
rect 68284 358776 68336 358828
rect 64144 358096 64196 358148
rect 65432 358096 65484 358148
rect 3240 357552 3292 357604
rect 6368 357552 6420 357604
rect 60188 356464 60240 356516
rect 64236 356464 64288 356516
rect 49608 353948 49660 354000
rect 60188 353948 60240 354000
rect 93124 352384 93176 352436
rect 95884 352384 95936 352436
rect 417424 351908 417476 351960
rect 580080 351908 580132 351960
rect 46204 350548 46256 350600
rect 49608 350548 49660 350600
rect 185584 350548 185636 350600
rect 186964 350548 187016 350600
rect 195244 346332 195296 346384
rect 198004 346332 198056 346384
rect 45376 342932 45428 342984
rect 46204 342932 46256 342984
rect 184204 338716 184256 338768
rect 185584 338716 185636 338768
rect 94412 332120 94464 332172
rect 100024 332120 100076 332172
rect 62856 331848 62908 331900
rect 88340 331848 88392 331900
rect 91744 329400 91796 329452
rect 94412 329400 94464 329452
rect 182824 329128 182876 329180
rect 184204 329128 184256 329180
rect 194048 328040 194100 328092
rect 195244 328040 195296 328092
rect 397000 324300 397052 324352
rect 580080 324300 580132 324352
rect 183376 322192 183428 322244
rect 194048 322192 194100 322244
rect 181444 320152 181496 320204
rect 183376 320152 183428 320204
rect 62764 319404 62816 319456
rect 64144 319404 64196 319456
rect 3240 318792 3292 318844
rect 24216 318792 24268 318844
rect 61476 318384 61528 318436
rect 62856 318384 62908 318436
rect 84844 315256 84896 315308
rect 104900 315256 104952 315308
rect 179512 314644 179564 314696
rect 181444 314644 181496 314696
rect 398196 311856 398248 311908
rect 580080 311856 580132 311908
rect 60004 311176 60056 311228
rect 61476 311176 61528 311228
rect 178684 309544 178736 309596
rect 179512 309544 179564 309596
rect 176660 305192 176712 305244
rect 178684 305192 178736 305244
rect 170128 304240 170180 304292
rect 176660 304240 176712 304292
rect 180064 302064 180116 302116
rect 182824 302064 182876 302116
rect 169024 300228 169076 300280
rect 170128 300228 170180 300280
rect 60832 299412 60884 299464
rect 62764 299412 62816 299464
rect 414664 298120 414716 298172
rect 580080 298120 580132 298172
rect 90364 298052 90416 298104
rect 93124 298052 93176 298104
rect 167644 295332 167696 295384
rect 169024 295332 169076 295384
rect 60096 293972 60148 294024
rect 60832 293972 60884 294024
rect 2780 292816 2832 292868
rect 4896 292816 4948 292868
rect 58624 291116 58676 291168
rect 60004 291116 60056 291168
rect 175648 290980 175700 291032
rect 180064 290980 180116 291032
rect 169024 289076 169076 289128
rect 175648 289076 175700 289128
rect 57244 287648 57296 287700
rect 71780 287648 71832 287700
rect 56508 284248 56560 284300
rect 58624 284316 58676 284368
rect 82084 284248 82136 284300
rect 84844 284316 84896 284368
rect 57980 282888 58032 282940
rect 60096 282888 60148 282940
rect 54300 281120 54352 281172
rect 56508 281120 56560 281172
rect 60004 280780 60056 280832
rect 169760 280780 169812 280832
rect 53288 278808 53340 278860
rect 54300 278808 54352 278860
rect 54484 278808 54536 278860
rect 57888 278808 57940 278860
rect 162860 278672 162912 278724
rect 167644 278740 167696 278792
rect 53840 277312 53892 277364
rect 57244 277380 57296 277432
rect 55864 276632 55916 276684
rect 82084 276632 82136 276684
rect 53104 274660 53156 274712
rect 53840 274660 53892 274712
rect 159364 274660 159416 274712
rect 162860 274660 162912 274712
rect 166264 273164 166316 273216
rect 169024 273232 169076 273284
rect 51816 272076 51868 272128
rect 53288 272076 53340 272128
rect 396908 271872 396960 271924
rect 579804 271872 579856 271924
rect 86960 270648 87012 270700
rect 90364 270648 90416 270700
rect 77944 268336 77996 268388
rect 86960 268336 87012 268388
rect 56600 268064 56652 268116
rect 60004 268064 60056 268116
rect 3056 266364 3108 266416
rect 40684 266364 40736 266416
rect 53196 266364 53248 266416
rect 54484 266364 54536 266416
rect 54576 266364 54628 266416
rect 55864 266364 55916 266416
rect 51724 264868 51776 264920
rect 56508 264936 56560 264988
rect 164240 264936 164292 264988
rect 166264 264936 166316 264988
rect 49700 263576 49752 263628
rect 51816 263576 51868 263628
rect 53288 263576 53340 263628
rect 54576 263576 54628 263628
rect 156604 261944 156656 261996
rect 159364 261944 159416 261996
rect 162124 260040 162176 260092
rect 164240 260040 164292 260092
rect 46940 258952 46992 259004
rect 49700 258952 49752 259004
rect 398288 258068 398340 258120
rect 579988 258068 580040 258120
rect 50436 256640 50488 256692
rect 53288 256708 53340 256760
rect 154028 256708 154080 256760
rect 156604 256708 156656 256760
rect 45560 255280 45612 255332
rect 46940 255280 46992 255332
rect 151084 255280 151136 255332
rect 154028 255280 154080 255332
rect 3148 253920 3200 253972
rect 22744 253920 22796 253972
rect 46204 253852 46256 253904
rect 53196 253988 53248 254040
rect 47584 253920 47636 253972
rect 50436 253920 50488 253972
rect 51816 252560 51868 252612
rect 53104 252560 53156 252612
rect 50344 250792 50396 250844
rect 51816 250792 51868 250844
rect 75184 249704 75236 249756
rect 77944 249704 77996 249756
rect 89168 249704 89220 249756
rect 91744 249704 91796 249756
rect 160100 245896 160152 245948
rect 162124 245896 162176 245948
rect 45836 245624 45888 245676
rect 47584 245624 47636 245676
rect 49700 245624 49752 245676
rect 51724 245624 51776 245676
rect 145196 245624 145248 245676
rect 151084 245624 151136 245676
rect 45192 245556 45244 245608
rect 46204 245556 46256 245608
rect 81440 244876 81492 244928
rect 89168 244876 89220 244928
rect 413284 244264 413336 244316
rect 579988 244264 580040 244316
rect 75092 242972 75144 243024
rect 81440 242972 81492 243024
rect 45744 242836 45796 242888
rect 49700 242904 49752 242956
rect 142988 241816 143040 241868
rect 145196 241816 145248 241868
rect 45100 240932 45152 240984
rect 75092 240932 75144 240984
rect 44916 240864 44968 240916
rect 75184 240864 75236 240916
rect 45376 240796 45428 240848
rect 142988 240796 143040 240848
rect 46848 240728 46900 240780
rect 160100 240728 160152 240780
rect 45652 240388 45704 240440
rect 50344 240388 50396 240440
rect 2780 240184 2832 240236
rect 4988 240184 5040 240236
rect 395344 239980 395396 240032
rect 396632 239980 396684 240032
rect 395436 239776 395488 239828
rect 44824 239708 44876 239760
rect 46848 239708 46900 239760
rect 45468 238756 45520 238808
rect 45836 238756 45888 238808
rect 396540 238688 396592 238740
rect 45744 233044 45796 233096
rect 45652 232976 45704 233028
rect 45468 232908 45520 232960
rect 45836 232908 45888 232960
rect 62764 232364 62816 232416
rect 80704 232364 80756 232416
rect 395436 232364 395488 232416
rect 396540 232364 396592 232416
rect 45376 231956 45428 232008
rect 46572 231956 46624 232008
rect 45100 231888 45152 231940
rect 45284 231820 45336 231872
rect 46848 231820 46900 231872
rect 393964 231820 394016 231872
rect 580080 231820 580132 231872
rect 49148 231752 49200 231804
rect 44824 231684 44876 231736
rect 49792 231684 49844 231736
rect 45836 231140 45888 231192
rect 142160 231140 142212 231192
rect 3332 231072 3384 231124
rect 180800 231072 180852 231124
rect 385684 231072 385736 231124
rect 396632 231072 396684 231124
rect 45192 231004 45244 231056
rect 64880 231004 64932 231056
rect 46572 230460 46624 230512
rect 49700 230392 49752 230444
rect 395344 230392 395396 230444
rect 396448 230392 396500 230444
rect 49792 230120 49844 230172
rect 55128 230120 55180 230172
rect 166264 229712 166316 229764
rect 176660 229712 176712 229764
rect 45008 229032 45060 229084
rect 47032 229032 47084 229084
rect 157984 228420 158036 228472
rect 266544 228420 266596 228472
rect 297364 228420 297416 228472
rect 327080 228420 327132 228472
rect 236644 228352 236696 228404
rect 386512 228352 386564 228404
rect 142160 228284 142212 228336
rect 143540 228284 143592 228336
rect 391204 227672 391256 227724
rect 395436 227740 395488 227792
rect 49700 226312 49752 226364
rect 44916 226244 44968 226296
rect 50436 226244 50488 226296
rect 64880 226312 64932 226364
rect 69572 226312 69624 226364
rect 56232 226244 56284 226296
rect 47032 225700 47084 225752
rect 53840 225700 53892 225752
rect 46940 224952 46992 225004
rect 50344 224884 50396 224936
rect 389824 223048 389876 223100
rect 394332 223048 394384 223100
rect 55220 222912 55272 222964
rect 57336 222912 57388 222964
rect 53840 222844 53892 222896
rect 69664 222844 69716 222896
rect 49148 222164 49200 222216
rect 55128 222096 55180 222148
rect 56232 222096 56284 222148
rect 57244 222096 57296 222148
rect 378048 220804 378100 220856
rect 385684 220804 385736 220856
rect 69664 220056 69716 220108
rect 79324 220056 79376 220108
rect 143540 220056 143592 220108
rect 158628 220056 158680 220108
rect 69664 218628 69716 218680
rect 71872 218628 71924 218680
rect 119436 218016 119488 218068
rect 580080 218016 580132 218068
rect 57336 217268 57388 217320
rect 67548 217268 67600 217320
rect 62764 215908 62816 215960
rect 70400 215908 70452 215960
rect 367744 215908 367796 215960
rect 378048 215908 378100 215960
rect 67548 215568 67600 215620
rect 69020 215568 69072 215620
rect 50436 215092 50488 215144
rect 54484 215092 54536 215144
rect 71872 214548 71924 214600
rect 73988 214548 74040 214600
rect 80704 214548 80756 214600
rect 91744 214548 91796 214600
rect 55220 214072 55272 214124
rect 57336 214072 57388 214124
rect 3332 213936 3384 213988
rect 180984 213936 181036 213988
rect 50344 213868 50396 213920
rect 53104 213868 53156 213920
rect 158720 213868 158772 213920
rect 160100 213868 160152 213920
rect 69020 213528 69072 213580
rect 71044 213528 71096 213580
rect 70400 212984 70452 213036
rect 73804 212984 73856 213036
rect 389916 212168 389968 212220
rect 391204 212168 391256 212220
rect 160100 211148 160152 211200
rect 57244 211080 57296 211132
rect 58624 211080 58676 211132
rect 162860 211080 162912 211132
rect 378784 210400 378836 210452
rect 395344 210400 395396 210452
rect 73988 209720 74040 209772
rect 75460 209720 75512 209772
rect 53104 209448 53156 209500
rect 54576 209448 54628 209500
rect 162860 209108 162912 209160
rect 164240 209108 164292 209160
rect 79324 209040 79376 209092
rect 91100 209040 91152 209092
rect 71044 208904 71096 208956
rect 73896 208904 73948 208956
rect 57336 208360 57388 208412
rect 63500 208292 63552 208344
rect 75460 208292 75512 208344
rect 77576 208292 77628 208344
rect 91744 208292 91796 208344
rect 95148 208292 95200 208344
rect 164240 206660 164292 206712
rect 166356 206660 166408 206712
rect 91100 206252 91152 206304
rect 104716 206252 104768 206304
rect 356704 206252 356756 206304
rect 367744 206252 367796 206304
rect 189724 205640 189776 205692
rect 580080 205640 580132 205692
rect 95148 204892 95200 204944
rect 106648 204892 106700 204944
rect 77576 204824 77628 204876
rect 80060 204824 80112 204876
rect 63500 204212 63552 204264
rect 65524 204212 65576 204264
rect 58624 202784 58676 202836
rect 63500 202784 63552 202836
rect 80060 202784 80112 202836
rect 81808 202784 81860 202836
rect 104716 202784 104768 202836
rect 108672 202784 108724 202836
rect 106648 202716 106700 202768
rect 110236 202716 110288 202768
rect 2964 201492 3016 201544
rect 22836 201492 22888 201544
rect 45560 201424 45612 201476
rect 47584 201424 47636 201476
rect 73804 199384 73856 199436
rect 81440 199384 81492 199436
rect 81808 199384 81860 199436
rect 88984 199384 89036 199436
rect 155960 199384 156012 199436
rect 296720 199384 296772 199436
rect 63500 197956 63552 198008
rect 69572 197956 69624 198008
rect 110236 197956 110288 198008
rect 117320 197956 117372 198008
rect 148968 197956 149020 198008
rect 207020 197956 207072 198008
rect 108672 197480 108724 197532
rect 111064 197480 111116 197532
rect 154488 197412 154540 197464
rect 155960 197412 156012 197464
rect 54576 197276 54628 197328
rect 56508 197276 56560 197328
rect 73896 197276 73948 197328
rect 76288 197276 76340 197328
rect 152740 197276 152792 197328
rect 157984 197276 158036 197328
rect 147956 196732 148008 196784
rect 166264 196732 166316 196784
rect 160836 196664 160888 196716
rect 236644 196664 236696 196716
rect 81440 196596 81492 196648
rect 88340 196596 88392 196648
rect 151176 196596 151228 196648
rect 236000 196596 236052 196648
rect 69572 196120 69624 196172
rect 71780 196120 71832 196172
rect 56600 195916 56652 195968
rect 138112 195916 138164 195968
rect 157524 195916 157576 195968
rect 356060 195916 356112 195968
rect 76288 195848 76340 195900
rect 77944 195848 77996 195900
rect 86960 195848 87012 195900
rect 139400 195848 139452 195900
rect 157432 195848 157484 195900
rect 297364 195848 297416 195900
rect 115940 194556 115992 194608
rect 140780 194556 140832 194608
rect 117320 194352 117372 194404
rect 120724 194352 120776 194404
rect 88340 193536 88392 193588
rect 91744 193536 91796 193588
rect 71780 193128 71832 193180
rect 74264 193128 74316 193180
rect 166356 193128 166408 193180
rect 168472 193128 168524 193180
rect 180064 191836 180116 191888
rect 580080 191836 580132 191888
rect 88984 190612 89036 190664
rect 93860 190612 93912 190664
rect 140964 190952 141016 191004
rect 140780 190476 140832 190528
rect 144460 190476 144512 190528
rect 140780 190340 140832 190392
rect 145012 190272 145064 190324
rect 140872 190204 140924 190256
rect 120724 189252 120776 189304
rect 123668 189252 123720 189304
rect 144644 188912 144696 188964
rect 145012 188912 145064 188964
rect 93860 187892 93912 187944
rect 95884 187892 95936 187944
rect 3332 187688 3384 187740
rect 116584 187688 116636 187740
rect 166172 187620 166224 187672
rect 399484 187620 399536 187672
rect 54484 186940 54536 186992
rect 68284 186940 68336 186992
rect 371240 186940 371292 186992
rect 389824 186940 389876 186992
rect 56600 186396 56652 186448
rect 58624 186396 58676 186448
rect 387800 186328 387852 186380
rect 389916 186328 389968 186380
rect 74264 186260 74316 186312
rect 76564 186260 76616 186312
rect 111064 186260 111116 186312
rect 113824 186260 113876 186312
rect 168472 184832 168524 184884
rect 170404 184832 170456 184884
rect 369124 183880 369176 183932
rect 371240 183880 371292 183932
rect 385040 183472 385092 183524
rect 387800 183540 387852 183592
rect 123668 182112 123720 182164
rect 126520 182112 126572 182164
rect 144644 181500 144696 181552
rect 145196 181500 145248 181552
rect 3240 181432 3292 181484
rect 46204 181432 46256 181484
rect 121460 180072 121512 180124
rect 136364 180072 136416 180124
rect 384304 179392 384356 179444
rect 385040 179392 385092 179444
rect 158812 179324 158864 179376
rect 165160 179324 165212 179376
rect 580816 179324 580868 179376
rect 113824 178916 113876 178968
rect 117964 178916 118016 178968
rect 136364 178780 136416 178832
rect 136732 178780 136784 178832
rect 124864 178712 124916 178764
rect 136456 178712 136508 178764
rect 126520 178644 126572 178696
rect 153936 178644 153988 178696
rect 135996 177760 136048 177812
rect 136640 177760 136692 177812
rect 124220 177284 124272 177336
rect 136456 177284 136508 177336
rect 68284 176604 68336 176656
rect 76656 176604 76708 176656
rect 149244 176604 149296 176656
rect 126980 176060 127032 176112
rect 135996 176060 136048 176112
rect 141792 176060 141844 176112
rect 154396 176400 154448 176452
rect 125600 175924 125652 175976
rect 136364 175992 136416 176044
rect 160468 175924 160520 175976
rect 159180 175856 159232 175908
rect 163596 175856 163648 175908
rect 159088 175788 159140 175840
rect 162492 175788 162544 175840
rect 141608 175652 141660 175704
rect 149336 175652 149388 175704
rect 144460 175516 144512 175568
rect 148692 175516 148744 175568
rect 95884 175244 95936 175296
rect 58624 175176 58676 175228
rect 60648 175176 60700 175228
rect 77944 175176 77996 175228
rect 79416 175176 79468 175228
rect 100024 175176 100076 175228
rect 128360 175176 128412 175228
rect 136456 175176 136508 175228
rect 144092 174904 144144 174956
rect 142068 174836 142120 174888
rect 350540 174564 350592 174616
rect 356704 174564 356756 174616
rect 161480 174496 161532 174548
rect 133880 173884 133932 173936
rect 137284 173884 137336 173936
rect 165436 172932 165488 172984
rect 60648 172524 60700 172576
rect 131120 172524 131172 172576
rect 136640 172524 136692 172576
rect 63500 172456 63552 172508
rect 65524 172456 65576 172508
rect 66260 172456 66312 172508
rect 76564 172456 76616 172508
rect 79324 172456 79376 172508
rect 160468 172456 160520 172508
rect 162124 172456 162176 172508
rect 376116 172456 376168 172508
rect 378784 172524 378836 172576
rect 348424 172320 348476 172372
rect 350540 172320 350592 172372
rect 135260 171912 135312 171964
rect 138664 171912 138716 171964
rect 145472 171844 145524 171896
rect 157984 171844 158036 171896
rect 47584 171776 47636 171828
rect 61660 171776 61712 171828
rect 118700 171776 118752 171828
rect 580172 171776 580224 171828
rect 91744 171164 91796 171216
rect 94504 171164 94556 171216
rect 132500 171096 132552 171148
rect 136732 171096 136784 171148
rect 138020 171096 138072 171148
rect 140780 171096 140832 171148
rect 376024 170348 376076 170400
rect 384304 170348 384356 170400
rect 152372 170280 152424 170332
rect 156512 170280 156564 170332
rect 149336 170008 149388 170060
rect 150440 170008 150492 170060
rect 63500 169532 63552 169584
rect 65616 169532 65668 169584
rect 66260 169532 66312 169584
rect 69664 169532 69716 169584
rect 61660 168716 61712 168768
rect 63500 168716 63552 168768
rect 63500 166268 63552 166320
rect 75184 166268 75236 166320
rect 142436 166268 142488 166320
rect 142620 166268 142672 166320
rect 100024 165588 100076 165640
rect 188344 165588 188396 165640
rect 580172 165588 580224 165640
rect 102784 165520 102836 165572
rect 76656 164160 76708 164212
rect 81808 164160 81860 164212
rect 94504 164160 94556 164212
rect 97264 164160 97316 164212
rect 40684 163548 40736 163600
rect 182364 163548 182416 163600
rect 24216 163480 24268 163532
rect 182916 163480 182968 163532
rect 3332 162868 3384 162920
rect 179512 162868 179564 162920
rect 65616 162800 65668 162852
rect 71044 162800 71096 162852
rect 374000 162800 374052 162852
rect 376116 162800 376168 162852
rect 81808 161236 81860 161288
rect 85488 161236 85540 161288
rect 162124 160692 162176 160744
rect 179420 160692 179472 160744
rect 75184 157972 75236 158024
rect 86132 157972 86184 158024
rect 366732 157700 366784 157752
rect 373908 157700 373960 157752
rect 375012 157360 375064 157412
rect 376024 157360 376076 157412
rect 359464 156680 359516 156732
rect 369124 156680 369176 156732
rect 353944 156612 353996 156664
rect 366732 156612 366784 156664
rect 85488 155864 85540 155916
rect 90364 155864 90416 155916
rect 86132 154504 86184 154556
rect 91744 154504 91796 154556
rect 170404 153892 170456 153944
rect 172520 153892 172572 153944
rect 71044 153824 71096 153876
rect 100024 153824 100076 153876
rect 373356 153212 373408 153264
rect 375012 153212 375064 153264
rect 154488 152464 154540 152516
rect 169760 152464 169812 152516
rect 97264 152260 97316 152312
rect 103612 152260 103664 152312
rect 180156 151784 180208 151836
rect 580172 151784 580224 151836
rect 102784 151376 102836 151428
rect 104532 151376 104584 151428
rect 172520 150492 172572 150544
rect 176568 150492 176620 150544
rect 103612 149540 103664 149592
rect 109684 149540 109736 149592
rect 3332 149064 3384 149116
rect 24216 149064 24268 149116
rect 104532 148860 104584 148912
rect 106280 148860 106332 148912
rect 339868 146956 339920 147008
rect 353944 146956 353996 147008
rect 118792 146888 118844 146940
rect 580080 146888 580132 146940
rect 176660 146208 176712 146260
rect 178684 146208 178736 146260
rect 371884 146208 371936 146260
rect 373356 146208 373408 146260
rect 157984 145596 158036 145648
rect 164976 145596 165028 145648
rect 119068 145528 119120 145580
rect 477500 145528 477552 145580
rect 69664 144848 69716 144900
rect 71044 144848 71096 144900
rect 336004 144304 336056 144356
rect 339868 144304 339920 144356
rect 343640 144236 343692 144288
rect 348424 144236 348476 144288
rect 118976 144168 119028 144220
rect 580264 144168 580316 144220
rect 79416 143488 79468 143540
rect 80704 143488 80756 143540
rect 164976 143488 165028 143540
rect 168380 143488 168432 143540
rect 24124 143012 24176 143064
rect 182732 143012 182784 143064
rect 20076 142944 20128 142996
rect 182824 142944 182876 142996
rect 6276 142876 6328 142928
rect 182272 142876 182324 142928
rect 118332 142808 118384 142860
rect 398104 142808 398156 142860
rect 106280 142128 106332 142180
rect 330944 142128 330996 142180
rect 336004 142128 336056 142180
rect 109776 142060 109828 142112
rect 40040 141652 40092 141704
rect 181076 141652 181128 141704
rect 19984 141584 20036 141636
rect 182640 141584 182692 141636
rect 326344 141584 326396 141636
rect 343640 141584 343692 141636
rect 118516 141516 118568 141568
rect 398288 141516 398340 141568
rect 118424 141448 118476 141500
rect 398196 141448 398248 141500
rect 119160 141380 119212 141432
rect 580448 141380 580500 141432
rect 369860 140768 369912 140820
rect 371884 140768 371936 140820
rect 140688 140700 140740 140752
rect 142252 140700 142304 140752
rect 90364 140564 90416 140616
rect 94504 140564 94556 140616
rect 150532 140496 150584 140548
rect 154580 140496 154632 140548
rect 163688 140428 163740 140480
rect 174636 140428 174688 140480
rect 164516 140360 164568 140412
rect 176200 140360 176252 140412
rect 144460 140292 144512 140344
rect 160560 140292 160612 140344
rect 163504 140292 163556 140344
rect 178040 140292 178092 140344
rect 142528 140224 142580 140276
rect 173072 140224 173124 140276
rect 119344 140156 119396 140208
rect 412640 140156 412692 140208
rect 120724 140088 120776 140140
rect 542360 140088 542412 140140
rect 118884 140020 118936 140072
rect 580908 140020 580960 140072
rect 178684 139952 178736 140004
rect 179696 139952 179748 140004
rect 123668 139748 123720 139800
rect 124864 139748 124916 139800
rect 146484 139748 146536 139800
rect 148048 139748 148100 139800
rect 153476 139748 153528 139800
rect 158996 139748 159048 139800
rect 137744 139680 137796 139732
rect 139584 139680 139636 139732
rect 147496 139680 147548 139732
rect 149612 139680 149664 139732
rect 152464 139680 152516 139732
rect 157432 139680 157484 139732
rect 149520 139612 149572 139664
rect 152740 139612 152792 139664
rect 120632 138932 120684 138984
rect 158444 138932 158496 138984
rect 100024 138864 100076 138916
rect 182456 138864 182508 138916
rect 3608 138796 3660 138848
rect 179604 138796 179656 138848
rect 3424 138728 3476 138780
rect 182548 138728 182600 138780
rect 320180 138728 320232 138780
rect 330944 138728 330996 138780
rect 119252 138660 119304 138712
rect 580632 138660 580684 138712
rect 117872 137980 117924 138032
rect 580172 137980 580224 138032
rect 179696 137912 179748 137964
rect 181168 137912 181220 137964
rect 366364 137300 366416 137352
rect 369860 137300 369912 137352
rect 46204 137232 46256 137284
rect 117320 137232 117372 137284
rect 119528 137232 119580 137284
rect 359464 137232 359516 137284
rect 318248 136960 318300 137012
rect 320180 136960 320232 137012
rect 3424 136688 3476 136740
rect 116676 136688 116728 136740
rect 19984 136620 20036 136672
rect 182180 136620 182232 136672
rect 94504 136484 94556 136536
rect 100116 136484 100168 136536
rect 306748 135872 306800 135924
rect 318248 135872 318300 135924
rect 91744 134580 91796 134632
rect 94228 134580 94280 134632
rect 3424 133900 3476 133952
rect 117320 133900 117372 133952
rect 305000 133900 305052 133952
rect 306748 133900 306800 133952
rect 3608 132472 3660 132524
rect 117320 132472 117372 132524
rect 71044 131996 71096 132048
rect 72516 131996 72568 132048
rect 100116 131928 100168 131980
rect 105544 131928 105596 131980
rect 94228 131180 94280 131232
rect 99380 131180 99432 131232
rect 3332 131112 3384 131164
rect 117320 131112 117372 131164
rect 361948 129888 362000 129940
rect 366364 129888 366416 129940
rect 24216 129684 24268 129736
rect 117320 129684 117372 129736
rect 300768 128324 300820 128376
rect 305000 128324 305052 128376
rect 22836 128256 22888 128308
rect 117320 128256 117372 128308
rect 22744 126896 22796 126948
rect 117320 126896 117372 126948
rect 99380 126828 99432 126880
rect 106188 126828 106240 126880
rect 314660 126216 314712 126268
rect 326344 126216 326396 126268
rect 184204 125604 184256 125656
rect 580080 125604 580132 125656
rect 72516 125536 72568 125588
rect 73896 125536 73948 125588
rect 6368 124108 6420 124160
rect 117320 124108 117372 124160
rect 118608 124108 118660 124160
rect 119528 124108 119580 124160
rect 312176 123904 312228 123956
rect 314660 123904 314712 123956
rect 360936 123632 360988 123684
rect 361948 123632 362000 123684
rect 106188 123428 106240 123480
rect 115296 123428 115348 123480
rect 295248 123428 295300 123480
rect 300768 123428 300820 123480
rect 10324 122748 10376 122800
rect 117320 122748 117372 122800
rect 73896 122680 73948 122732
rect 75460 122680 75512 122732
rect 109776 121932 109828 121984
rect 111800 121932 111852 121984
rect 8944 121388 8996 121440
rect 117320 121388 117372 121440
rect 80704 120640 80756 120692
rect 82820 120640 82872 120692
rect 4804 120028 4856 120080
rect 117320 120028 117372 120080
rect 105544 119076 105596 119128
rect 109776 119076 109828 119128
rect 43444 118600 43496 118652
rect 117320 118600 117372 118652
rect 82820 118532 82872 118584
rect 86224 118532 86276 118584
rect 79324 118260 79376 118312
rect 81072 118260 81124 118312
rect 307024 117512 307076 117564
rect 312176 117512 312228 117564
rect 358820 117512 358872 117564
rect 360936 117512 360988 117564
rect 292580 117376 292632 117428
rect 295248 117376 295300 117428
rect 15844 117240 15896 117292
rect 117320 117240 117372 117292
rect 111800 117172 111852 117224
rect 115204 117172 115256 117224
rect 6184 115880 6236 115932
rect 117320 115880 117372 115932
rect 354680 115880 354732 115932
rect 358820 115880 358872 115932
rect 81072 115812 81124 115864
rect 82728 115812 82780 115864
rect 118148 114792 118200 114844
rect 119436 114792 119488 114844
rect 75460 114520 75512 114572
rect 81348 114452 81400 114504
rect 291108 114248 291160 114300
rect 292580 114248 292632 114300
rect 33784 113092 33836 113144
rect 117320 113092 117372 113144
rect 86224 112412 86276 112464
rect 87420 112412 87472 112464
rect 180248 111800 180300 111852
rect 580172 111800 580224 111852
rect 3240 111732 3292 111784
rect 19984 111732 20036 111784
rect 115296 111732 115348 111784
rect 117320 111732 117372 111784
rect 303620 111052 303672 111104
rect 307024 111052 307076 111104
rect 81348 110440 81400 110492
rect 117320 110372 117372 110424
rect 87420 109692 87472 109744
rect 97908 109692 97960 109744
rect 97908 108944 97960 108996
rect 117320 108944 117372 108996
rect 183468 108944 183520 108996
rect 354588 108944 354640 108996
rect 82820 107584 82872 107636
rect 117320 107584 117372 107636
rect 183468 107584 183520 107636
rect 291108 107652 291160 107704
rect 109684 107516 109736 107568
rect 112444 107516 112496 107568
rect 183468 106224 183520 106276
rect 410524 106224 410576 106276
rect 291844 105544 291896 105596
rect 303620 105544 303672 105596
rect 183468 104796 183520 104848
rect 409144 104796 409196 104848
rect 183468 103436 183520 103488
rect 407764 103436 407816 103488
rect 183468 102076 183520 102128
rect 544384 102076 544436 102128
rect 109776 102008 109828 102060
rect 115848 102008 115900 102060
rect 182824 100648 182876 100700
rect 406384 100648 406436 100700
rect 180340 99356 180392 99408
rect 580172 99356 580224 99408
rect 182824 99288 182876 99340
rect 405004 99288 405056 99340
rect 117964 98676 118016 98728
rect 120908 98676 120960 98728
rect 115204 97928 115256 97980
rect 116768 97928 116820 97980
rect 183468 97928 183520 97980
rect 403624 97928 403676 97980
rect 115848 95140 115900 95192
rect 120816 95140 120868 95192
rect 183468 95140 183520 95192
rect 400864 95140 400916 95192
rect 183468 93780 183520 93832
rect 418804 93780 418856 93832
rect 183468 92420 183520 92472
rect 417424 92420 417476 92472
rect 183468 90992 183520 91044
rect 414664 90992 414716 91044
rect 182272 89632 182324 89684
rect 413284 89632 413336 89684
rect 116768 88952 116820 89004
rect 117964 88952 118016 89004
rect 183468 88136 183520 88188
rect 189724 88136 189776 88188
rect 284944 87592 284996 87644
rect 291844 87592 291896 87644
rect 183468 86844 183520 86896
rect 188344 86844 188396 86896
rect 182272 85552 182324 85604
rect 580172 85552 580224 85604
rect 182180 85484 182232 85536
rect 184204 85484 184256 85536
rect 120908 85008 120960 85060
rect 120908 84804 120960 84856
rect 3148 84192 3200 84244
rect 120724 84192 120776 84244
rect 117964 81404 118016 81456
rect 120816 81336 120868 81388
rect 183468 80044 183520 80096
rect 555424 80044 555476 80096
rect 178960 79296 179012 79348
rect 580540 79296 580592 79348
rect 120632 78616 120684 78668
rect 124772 78616 124824 78668
rect 124956 78548 125008 78600
rect 4896 78480 4948 78532
rect 4068 78344 4120 78396
rect 3884 78208 3936 78260
rect 118792 78208 118844 78260
rect 122104 78072 122156 78124
rect 124864 78004 124916 78056
rect 112444 77936 112496 77988
rect 124772 77936 124824 77988
rect 125324 77868 125376 77920
rect 125830 77868 125882 77920
rect 121644 77800 121696 77852
rect 126106 77800 126158 77852
rect 126198 77800 126250 77852
rect 126382 77800 126434 77852
rect 126152 77664 126204 77716
rect 126336 77664 126388 77716
rect 126658 77664 126710 77716
rect 119804 77596 119856 77648
rect 125048 77460 125100 77512
rect 125876 77392 125928 77444
rect 126934 77868 126986 77920
rect 127026 77868 127078 77920
rect 127118 77868 127170 77920
rect 127210 77868 127262 77920
rect 127072 77732 127124 77784
rect 126980 77664 127032 77716
rect 127486 77868 127538 77920
rect 127670 77868 127722 77920
rect 127762 77868 127814 77920
rect 127854 77868 127906 77920
rect 127946 77868 127998 77920
rect 128130 77868 128182 77920
rect 128222 77868 128274 77920
rect 128314 77868 128366 77920
rect 127302 77800 127354 77852
rect 127394 77800 127446 77852
rect 127808 77732 127860 77784
rect 127900 77732 127952 77784
rect 127624 77664 127676 77716
rect 127992 77664 128044 77716
rect 128084 77664 128136 77716
rect 127256 77596 127308 77648
rect 127440 77596 127492 77648
rect 128314 77664 128366 77716
rect 127348 77392 127400 77444
rect 127716 77460 127768 77512
rect 128498 77868 128550 77920
rect 128590 77868 128642 77920
rect 128682 77868 128734 77920
rect 129142 77868 129194 77920
rect 129326 77868 129378 77920
rect 129418 77868 129470 77920
rect 129510 77868 129562 77920
rect 129602 77868 129654 77920
rect 129234 77800 129286 77852
rect 128544 77528 128596 77580
rect 128636 77528 128688 77580
rect 129096 77664 129148 77716
rect 129464 77732 129516 77784
rect 129372 77664 129424 77716
rect 129556 77664 129608 77716
rect 129188 77596 129240 77648
rect 129970 77868 130022 77920
rect 130154 77868 130206 77920
rect 130246 77868 130298 77920
rect 129924 77732 129976 77784
rect 130200 77664 130252 77716
rect 130016 77528 130068 77580
rect 128820 77460 128872 77512
rect 129280 77392 129332 77444
rect 130614 77868 130666 77920
rect 130706 77868 130758 77920
rect 130798 77868 130850 77920
rect 130982 77868 131034 77920
rect 131166 77868 131218 77920
rect 131258 77868 131310 77920
rect 131442 77868 131494 77920
rect 131534 77868 131586 77920
rect 131810 77868 131862 77920
rect 131902 77868 131954 77920
rect 130660 77732 130712 77784
rect 130752 77732 130804 77784
rect 131212 77732 131264 77784
rect 130844 77596 130896 77648
rect 130936 77596 130988 77648
rect 131120 77596 131172 77648
rect 131580 77596 131632 77648
rect 131672 77528 131724 77580
rect 131764 77460 131816 77512
rect 132178 77868 132230 77920
rect 132270 77868 132322 77920
rect 132454 77868 132506 77920
rect 132638 77868 132690 77920
rect 132730 77868 132782 77920
rect 133098 77868 133150 77920
rect 133374 77868 133426 77920
rect 133466 77868 133518 77920
rect 133558 77868 133610 77920
rect 133742 77868 133794 77920
rect 133926 77868 133978 77920
rect 134018 77868 134070 77920
rect 134110 77868 134162 77920
rect 134202 77868 134254 77920
rect 134478 77868 134530 77920
rect 134570 77868 134622 77920
rect 132316 77664 132368 77716
rect 132592 77732 132644 77784
rect 132822 77732 132874 77784
rect 132224 77596 132276 77648
rect 132684 77596 132736 77648
rect 132408 77528 132460 77580
rect 133236 77596 133288 77648
rect 133052 77528 133104 77580
rect 133144 77528 133196 77580
rect 133420 77460 133472 77512
rect 133880 77732 133932 77784
rect 133696 77528 133748 77580
rect 134064 77596 134116 77648
rect 134432 77732 134484 77784
rect 134340 77528 134392 77580
rect 133972 77460 134024 77512
rect 134846 77868 134898 77920
rect 134938 77868 134990 77920
rect 135030 77868 135082 77920
rect 135214 77868 135266 77920
rect 135306 77868 135358 77920
rect 135490 77868 135542 77920
rect 135582 77868 135634 77920
rect 135674 77868 135726 77920
rect 135858 77868 135910 77920
rect 135950 77868 136002 77920
rect 134800 77664 134852 77716
rect 134892 77664 134944 77716
rect 134984 77664 135036 77716
rect 135260 77664 135312 77716
rect 135352 77596 135404 77648
rect 135444 77596 135496 77648
rect 134708 77528 134760 77580
rect 135628 77664 135680 77716
rect 136134 77800 136186 77852
rect 136088 77664 136140 77716
rect 135904 77596 135956 77648
rect 136272 77596 136324 77648
rect 135996 77528 136048 77580
rect 136502 77868 136554 77920
rect 136778 77868 136830 77920
rect 136594 77800 136646 77852
rect 136732 77664 136784 77716
rect 136640 77596 136692 77648
rect 137330 77868 137382 77920
rect 137514 77868 137566 77920
rect 137606 77868 137658 77920
rect 137054 77800 137106 77852
rect 136548 77528 136600 77580
rect 136916 77528 136968 77580
rect 137468 77664 137520 77716
rect 137790 77868 137842 77920
rect 137882 77868 137934 77920
rect 137974 77868 138026 77920
rect 138158 77868 138210 77920
rect 138250 77868 138302 77920
rect 138342 77868 138394 77920
rect 138526 77868 138578 77920
rect 138618 77868 138670 77920
rect 138802 77868 138854 77920
rect 138986 77868 139038 77920
rect 137836 77732 137888 77784
rect 137928 77664 137980 77716
rect 137652 77528 137704 77580
rect 138296 77732 138348 77784
rect 138204 77664 138256 77716
rect 138112 77528 138164 77580
rect 135536 77460 135588 77512
rect 131856 77392 131908 77444
rect 133512 77392 133564 77444
rect 138848 77596 138900 77648
rect 138940 77596 138992 77648
rect 138756 77528 138808 77580
rect 139170 77868 139222 77920
rect 139354 77868 139406 77920
rect 139446 77868 139498 77920
rect 139538 77868 139590 77920
rect 139630 77868 139682 77920
rect 139722 77868 139774 77920
rect 140182 77868 140234 77920
rect 140366 77868 140418 77920
rect 140734 77868 140786 77920
rect 140826 77868 140878 77920
rect 139032 77460 139084 77512
rect 139492 77664 139544 77716
rect 139308 77596 139360 77648
rect 139400 77596 139452 77648
rect 140550 77800 140602 77852
rect 140228 77596 140280 77648
rect 140412 77596 140464 77648
rect 139952 77528 140004 77580
rect 139768 77460 139820 77512
rect 139860 77460 139912 77512
rect 140780 77664 140832 77716
rect 140688 77596 140740 77648
rect 126704 77324 126756 77376
rect 118792 77188 118844 77240
rect 130568 77324 130620 77376
rect 130752 77324 130804 77376
rect 134156 77256 134208 77308
rect 138664 77392 138716 77444
rect 138572 77324 138624 77376
rect 139584 77324 139636 77376
rect 141010 77868 141062 77920
rect 141102 77868 141154 77920
rect 141194 77868 141246 77920
rect 141286 77868 141338 77920
rect 141562 77868 141614 77920
rect 141654 77868 141706 77920
rect 141838 77868 141890 77920
rect 141930 77868 141982 77920
rect 141148 77596 141200 77648
rect 141332 77460 141384 77512
rect 141240 77392 141292 77444
rect 141148 77324 141200 77376
rect 138572 77188 138624 77240
rect 140964 77188 141016 77240
rect 141608 77732 141660 77784
rect 141884 77664 141936 77716
rect 141792 77596 141844 77648
rect 142206 77868 142258 77920
rect 142298 77868 142350 77920
rect 142482 77868 142534 77920
rect 142574 77868 142626 77920
rect 142666 77868 142718 77920
rect 142758 77868 142810 77920
rect 142252 77664 142304 77716
rect 142436 77596 142488 77648
rect 143034 77800 143086 77852
rect 142620 77664 142672 77716
rect 142712 77596 142764 77648
rect 142344 77528 142396 77580
rect 142896 77528 142948 77580
rect 142160 77460 142212 77512
rect 142344 77392 142396 77444
rect 142620 77324 142672 77376
rect 143310 77868 143362 77920
rect 143494 77800 143546 77852
rect 143862 77868 143914 77920
rect 143954 77868 144006 77920
rect 144046 77868 144098 77920
rect 144414 77868 144466 77920
rect 144506 77868 144558 77920
rect 143632 77528 143684 77580
rect 144138 77800 144190 77852
rect 144092 77664 144144 77716
rect 144000 77460 144052 77512
rect 143264 77392 143316 77444
rect 143448 77392 143500 77444
rect 143908 77392 143960 77444
rect 144184 77528 144236 77580
rect 143540 77256 143592 77308
rect 144460 77664 144512 77716
rect 144552 77596 144604 77648
rect 180340 78684 180392 78736
rect 174544 78616 174596 78668
rect 145150 77800 145202 77852
rect 145242 77800 145294 77852
rect 145426 77868 145478 77920
rect 145518 77868 145570 77920
rect 145610 77868 145662 77920
rect 145334 77732 145386 77784
rect 145196 77528 145248 77580
rect 145426 77664 145478 77716
rect 145380 77528 145432 77580
rect 145610 77732 145662 77784
rect 145794 77868 145846 77920
rect 146070 77868 146122 77920
rect 145656 77460 145708 77512
rect 145288 77392 145340 77444
rect 145472 77392 145524 77444
rect 144920 77256 144972 77308
rect 145472 77256 145524 77308
rect 145840 77528 145892 77580
rect 145840 77392 145892 77444
rect 146714 77868 146766 77920
rect 147174 77868 147226 77920
rect 147266 77868 147318 77920
rect 147358 77868 147410 77920
rect 147450 77868 147502 77920
rect 147542 77868 147594 77920
rect 147634 77868 147686 77920
rect 147726 77868 147778 77920
rect 148002 77868 148054 77920
rect 148278 77868 148330 77920
rect 148370 77868 148422 77920
rect 148462 77868 148514 77920
rect 148554 77868 148606 77920
rect 148738 77868 148790 77920
rect 148830 77868 148882 77920
rect 148922 77868 148974 77920
rect 149014 77868 149066 77920
rect 149198 77868 149250 77920
rect 149290 77868 149342 77920
rect 149382 77868 149434 77920
rect 149474 77868 149526 77920
rect 146346 77800 146398 77852
rect 146438 77800 146490 77852
rect 146990 77732 147042 77784
rect 146852 77596 146904 77648
rect 146944 77528 146996 77580
rect 146392 77460 146444 77512
rect 146668 77460 146720 77512
rect 147220 77732 147272 77784
rect 147312 77664 147364 77716
rect 147404 77664 147456 77716
rect 147680 77732 147732 77784
rect 147496 77596 147548 77648
rect 148324 77732 148376 77784
rect 148324 77596 148376 77648
rect 147956 77528 148008 77580
rect 146300 77392 146352 77444
rect 148232 77392 148284 77444
rect 148784 77664 148836 77716
rect 148876 77664 148928 77716
rect 148968 77664 149020 77716
rect 148692 77528 148744 77580
rect 148508 77324 148560 77376
rect 149244 77732 149296 77784
rect 149336 77664 149388 77716
rect 149428 77664 149480 77716
rect 149750 77868 149802 77920
rect 149842 77868 149894 77920
rect 149934 77868 149986 77920
rect 150118 77868 150170 77920
rect 150302 77868 150354 77920
rect 150394 77868 150446 77920
rect 150486 77868 150538 77920
rect 150578 77868 150630 77920
rect 149658 77732 149710 77784
rect 149796 77732 149848 77784
rect 149888 77732 149940 77784
rect 149704 77596 149756 77648
rect 150164 77596 150216 77648
rect 149980 77528 150032 77580
rect 150348 77732 150400 77784
rect 149612 77460 149664 77512
rect 149336 77324 149388 77376
rect 150532 77664 150584 77716
rect 151038 77868 151090 77920
rect 151130 77868 151182 77920
rect 151314 77868 151366 77920
rect 151498 77868 151550 77920
rect 151774 77868 151826 77920
rect 151866 77868 151918 77920
rect 150992 77664 151044 77716
rect 151176 77596 151228 77648
rect 151728 77732 151780 77784
rect 151820 77664 151872 77716
rect 151360 77528 151412 77580
rect 152142 77868 152194 77920
rect 152418 77868 152470 77920
rect 152510 77868 152562 77920
rect 152694 77868 152746 77920
rect 152878 77868 152930 77920
rect 152970 77868 153022 77920
rect 153062 77868 153114 77920
rect 153246 77868 153298 77920
rect 152188 77596 152240 77648
rect 152280 77528 152332 77580
rect 152004 77460 152056 77512
rect 152464 77664 152516 77716
rect 152556 77596 152608 77648
rect 152832 77664 152884 77716
rect 152924 77664 152976 77716
rect 152648 77528 152700 77580
rect 153200 77528 153252 77580
rect 153890 77868 153942 77920
rect 153798 77800 153850 77852
rect 153752 77664 153804 77716
rect 154166 77800 154218 77852
rect 154258 77800 154310 77852
rect 154120 77664 154172 77716
rect 153936 77596 153988 77648
rect 153384 77460 153436 77512
rect 154396 77460 154448 77512
rect 154810 77868 154862 77920
rect 154948 77596 155000 77648
rect 149060 77256 149112 77308
rect 152372 77256 152424 77308
rect 154672 77324 154724 77376
rect 154856 77324 154908 77376
rect 155270 77868 155322 77920
rect 155362 77868 155414 77920
rect 155454 77868 155506 77920
rect 155730 77868 155782 77920
rect 155822 77868 155874 77920
rect 155224 77528 155276 77580
rect 155408 77664 155460 77716
rect 155868 77732 155920 77784
rect 155592 77596 155644 77648
rect 156098 77868 156150 77920
rect 156374 77868 156426 77920
rect 156466 77868 156518 77920
rect 156558 77868 156610 77920
rect 156420 77732 156472 77784
rect 156236 77596 156288 77648
rect 156512 77596 156564 77648
rect 156742 77868 156794 77920
rect 156834 77868 156886 77920
rect 157294 77868 157346 77920
rect 156788 77732 156840 77784
rect 157478 77868 157530 77920
rect 157570 77868 157622 77920
rect 157662 77868 157714 77920
rect 157846 77868 157898 77920
rect 157938 77868 157990 77920
rect 158214 77868 158266 77920
rect 158306 77868 158358 77920
rect 157340 77664 157392 77716
rect 157156 77596 157208 77648
rect 157524 77732 157576 77784
rect 157708 77732 157760 77784
rect 157708 77596 157760 77648
rect 157800 77596 157852 77648
rect 158260 77664 158312 77716
rect 156604 77528 156656 77580
rect 156880 77528 156932 77580
rect 156972 77528 157024 77580
rect 157248 77528 157300 77580
rect 156972 77392 157024 77444
rect 158076 77460 158128 77512
rect 158444 77460 158496 77512
rect 158858 77868 158910 77920
rect 158950 77868 159002 77920
rect 159042 77868 159094 77920
rect 159134 77868 159186 77920
rect 159594 77868 159646 77920
rect 159778 77868 159830 77920
rect 159870 77868 159922 77920
rect 159962 77868 160014 77920
rect 160054 77868 160106 77920
rect 160146 77868 160198 77920
rect 159318 77800 159370 77852
rect 159410 77800 159462 77852
rect 158812 77596 158864 77648
rect 158996 77596 159048 77648
rect 159088 77596 159140 77648
rect 158904 77528 158956 77580
rect 159180 77528 159232 77580
rect 159272 77460 159324 77512
rect 159640 77596 159692 77648
rect 159916 77596 159968 77648
rect 160008 77596 160060 77648
rect 160100 77596 160152 77648
rect 160330 77868 160382 77920
rect 159364 77324 159416 77376
rect 156696 77256 156748 77308
rect 158444 77256 158496 77308
rect 160284 77528 160336 77580
rect 160514 77868 160566 77920
rect 160606 77800 160658 77852
rect 160560 77596 160612 77648
rect 160882 77868 160934 77920
rect 160974 77868 161026 77920
rect 160928 77664 160980 77716
rect 160744 77596 160796 77648
rect 160652 77528 160704 77580
rect 161020 77528 161072 77580
rect 161618 77868 161670 77920
rect 161710 77868 161762 77920
rect 161802 77868 161854 77920
rect 161250 77800 161302 77852
rect 161342 77800 161394 77852
rect 161434 77800 161486 77852
rect 161296 77664 161348 77716
rect 161388 77664 161440 77716
rect 161986 77868 162038 77920
rect 162170 77868 162222 77920
rect 162078 77800 162130 77852
rect 161756 77528 161808 77580
rect 161204 77460 161256 77512
rect 161664 77460 161716 77512
rect 162032 77664 162084 77716
rect 162124 77664 162176 77716
rect 162446 77868 162498 77920
rect 162630 77868 162682 77920
rect 162308 77596 162360 77648
rect 161940 77528 161992 77580
rect 162216 77392 162268 77444
rect 162814 77868 162866 77920
rect 162906 77868 162958 77920
rect 162998 77868 163050 77920
rect 162492 77460 162544 77512
rect 162584 77392 162636 77444
rect 162860 77596 162912 77648
rect 162768 77528 162820 77580
rect 163366 77868 163418 77920
rect 163550 77868 163602 77920
rect 163642 77868 163694 77920
rect 163734 77868 163786 77920
rect 163826 77868 163878 77920
rect 163918 77868 163970 77920
rect 163412 77732 163464 77784
rect 163504 77596 163556 77648
rect 163964 77732 164016 77784
rect 163688 77664 163740 77716
rect 163780 77664 163832 77716
rect 175924 78412 175976 78464
rect 164286 77868 164338 77920
rect 164470 77868 164522 77920
rect 164562 77868 164614 77920
rect 164930 77868 164982 77920
rect 165022 77868 165074 77920
rect 165114 77868 165166 77920
rect 165206 77868 165258 77920
rect 163872 77596 163924 77648
rect 163596 77528 163648 77580
rect 162952 77460 163004 77512
rect 164332 77596 164384 77648
rect 164148 77528 164200 77580
rect 164516 77664 164568 77716
rect 165574 77800 165626 77852
rect 165068 77664 165120 77716
rect 165160 77664 165212 77716
rect 164424 77460 164476 77512
rect 165252 77596 165304 77648
rect 164884 77528 164936 77580
rect 164976 77528 165028 77580
rect 165942 77868 165994 77920
rect 165896 77732 165948 77784
rect 166126 77868 166178 77920
rect 166218 77868 166270 77920
rect 166494 77868 166546 77920
rect 166586 77868 166638 77920
rect 166678 77868 166730 77920
rect 166080 77596 166132 77648
rect 164700 77460 164752 77512
rect 166540 77664 166592 77716
rect 166632 77664 166684 77716
rect 166816 77596 166868 77648
rect 166356 77460 166408 77512
rect 166908 77460 166960 77512
rect 167690 77868 167742 77920
rect 167782 77868 167834 77920
rect 168150 77868 168202 77920
rect 168334 77868 168386 77920
rect 168426 77868 168478 77920
rect 168978 77868 169030 77920
rect 168104 77732 168156 77784
rect 167736 77664 167788 77716
rect 168288 77596 168340 77648
rect 168886 77800 168938 77852
rect 168932 77596 168984 77648
rect 169622 77868 169674 77920
rect 169990 77868 170042 77920
rect 169714 77800 169766 77852
rect 174636 78276 174688 78328
rect 170358 77868 170410 77920
rect 170726 77868 170778 77920
rect 174728 78208 174780 78260
rect 174820 78140 174872 78192
rect 180064 78072 180116 78124
rect 393964 78004 394016 78056
rect 171186 77868 171238 77920
rect 171278 77868 171330 77920
rect 171370 77868 171422 77920
rect 171738 77868 171790 77920
rect 171094 77800 171146 77852
rect 170312 77732 170364 77784
rect 170680 77732 170732 77784
rect 169576 77664 169628 77716
rect 169668 77664 169720 77716
rect 169990 77664 170042 77716
rect 171922 77868 171974 77920
rect 172014 77868 172066 77920
rect 173026 77868 173078 77920
rect 170404 77596 170456 77648
rect 171692 77596 171744 77648
rect 171784 77596 171836 77648
rect 171508 77528 171560 77580
rect 174636 77936 174688 77988
rect 173670 77868 173722 77920
rect 173762 77868 173814 77920
rect 174544 77868 174596 77920
rect 580356 77936 580408 77988
rect 176108 77800 176160 77852
rect 396908 77800 396960 77852
rect 171968 77664 172020 77716
rect 172106 77664 172158 77716
rect 175832 77664 175884 77716
rect 175924 77664 175976 77716
rect 231860 77664 231912 77716
rect 172244 77596 172296 77648
rect 172060 77528 172112 77580
rect 173624 77596 173676 77648
rect 200120 77596 200172 77648
rect 168564 77460 168616 77512
rect 175832 77528 175884 77580
rect 175924 77528 175976 77580
rect 284300 77528 284352 77580
rect 252560 77460 252612 77512
rect 167552 77392 167604 77444
rect 172060 77392 172112 77444
rect 172244 77392 172296 77444
rect 302240 77392 302292 77444
rect 165436 77324 165488 77376
rect 165804 77324 165856 77376
rect 320180 77324 320232 77376
rect 161572 77256 161624 77308
rect 462412 77256 462464 77308
rect 147588 77188 147640 77240
rect 149152 77188 149204 77240
rect 162952 77188 163004 77240
rect 163596 77188 163648 77240
rect 170312 77188 170364 77240
rect 171692 77188 171744 77240
rect 116584 77120 116636 77172
rect 171968 77120 172020 77172
rect 180248 77120 180300 77172
rect 116676 77052 116728 77104
rect 173992 77052 174044 77104
rect 120724 76984 120776 77036
rect 174176 76984 174228 77036
rect 142252 76916 142304 76968
rect 213920 76916 213972 76968
rect 144276 76848 144328 76900
rect 144552 76848 144604 76900
rect 146944 76848 146996 76900
rect 4988 76576 5040 76628
rect 124772 76712 124824 76764
rect 130936 76712 130988 76764
rect 147588 76780 147640 76832
rect 152004 76780 152056 76832
rect 155316 76780 155368 76832
rect 162676 76780 162728 76832
rect 158628 76712 158680 76764
rect 267740 76848 267792 76900
rect 165528 76780 165580 76832
rect 306380 76780 306432 76832
rect 154672 76644 154724 76696
rect 155316 76644 155368 76696
rect 155684 76644 155736 76696
rect 156144 76644 156196 76696
rect 157524 76644 157576 76696
rect 158720 76644 158772 76696
rect 121368 76440 121420 76492
rect 126980 76440 127032 76492
rect 125784 76304 125836 76356
rect 126152 76304 126204 76356
rect 127256 76304 127308 76356
rect 127624 76304 127676 76356
rect 129832 76304 129884 76356
rect 130108 76304 130160 76356
rect 130292 76304 130344 76356
rect 130752 76304 130804 76356
rect 130016 76236 130068 76288
rect 130476 76236 130528 76288
rect 127624 76168 127676 76220
rect 129096 76168 129148 76220
rect 126060 76100 126112 76152
rect 126244 76100 126296 76152
rect 146300 76440 146352 76492
rect 152372 76576 152424 76628
rect 161204 76576 161256 76628
rect 162216 76644 162268 76696
rect 167000 76712 167052 76764
rect 168656 76712 168708 76764
rect 170772 76712 170824 76764
rect 171140 76712 171192 76764
rect 175924 76712 175976 76764
rect 178408 76712 178460 76764
rect 431960 76712 432012 76764
rect 426440 76644 426492 76696
rect 156144 76508 156196 76560
rect 156788 76508 156840 76560
rect 160100 76508 160152 76560
rect 171048 76576 171100 76628
rect 171324 76576 171376 76628
rect 176108 76576 176160 76628
rect 176200 76576 176252 76628
rect 462320 76576 462372 76628
rect 164332 76508 164384 76560
rect 168748 76508 168800 76560
rect 170404 76508 170456 76560
rect 557540 76508 557592 76560
rect 156420 76372 156472 76424
rect 156788 76372 156840 76424
rect 146300 76304 146352 76356
rect 146852 76304 146904 76356
rect 161572 76304 161624 76356
rect 161940 76304 161992 76356
rect 156052 76236 156104 76288
rect 156420 76236 156472 76288
rect 164240 76440 164292 76492
rect 165344 76440 165396 76492
rect 167276 76440 167328 76492
rect 168104 76440 168156 76492
rect 168656 76440 168708 76492
rect 169392 76440 169444 76492
rect 171968 76440 172020 76492
rect 173900 76440 173952 76492
rect 163044 76372 163096 76424
rect 172060 76372 172112 76424
rect 172336 76372 172388 76424
rect 175832 76372 175884 76424
rect 162952 76304 163004 76356
rect 172244 76304 172296 76356
rect 174360 76236 174412 76288
rect 146576 76168 146628 76220
rect 147312 76168 147364 76220
rect 159548 76168 159600 76220
rect 159916 76168 159968 76220
rect 161940 76168 161992 76220
rect 165804 76168 165856 76220
rect 171140 76168 171192 76220
rect 172704 76168 172756 76220
rect 146392 76100 146444 76152
rect 146760 76100 146812 76152
rect 147680 76100 147732 76152
rect 150164 76100 150216 76152
rect 153108 76100 153160 76152
rect 158536 76100 158588 76152
rect 160468 76100 160520 76152
rect 167552 76100 167604 76152
rect 168012 76100 168064 76152
rect 169392 76100 169444 76152
rect 146576 76032 146628 76084
rect 159180 76032 159232 76084
rect 159916 76032 159968 76084
rect 160100 76032 160152 76084
rect 195980 76032 196032 76084
rect 148600 75964 148652 76016
rect 155592 75964 155644 76016
rect 157432 75964 157484 76016
rect 158352 75964 158404 76016
rect 161572 75964 161624 76016
rect 161756 75964 161808 76016
rect 165804 75964 165856 76016
rect 249800 75964 249852 76016
rect 121092 75828 121144 75880
rect 129188 75896 129240 75948
rect 152832 75896 152884 75948
rect 154120 75896 154172 75948
rect 157156 75896 157208 75948
rect 157524 75896 157576 75948
rect 159180 75896 159232 75948
rect 159364 75896 159416 75948
rect 162124 75896 162176 75948
rect 288440 75896 288492 75948
rect 153476 75828 153528 75880
rect 153936 75828 153988 75880
rect 154672 75828 154724 75880
rect 155132 75828 155184 75880
rect 155960 75828 156012 75880
rect 156328 75828 156380 75880
rect 156696 75828 156748 75880
rect 161940 75828 161992 75880
rect 125232 75760 125284 75812
rect 133512 75760 133564 75812
rect 141148 75760 141200 75812
rect 164884 75828 164936 75880
rect 163872 75760 163924 75812
rect 164056 75760 164108 75812
rect 128544 75692 128596 75744
rect 129372 75692 129424 75744
rect 139400 75692 139452 75744
rect 143632 75624 143684 75676
rect 144092 75624 144144 75676
rect 145012 75624 145064 75676
rect 165804 75692 165856 75744
rect 167920 75692 167972 75744
rect 168104 75692 168156 75744
rect 169024 75760 169076 75812
rect 169668 75760 169720 75812
rect 172612 75760 172664 75812
rect 284944 75760 284996 75812
rect 173164 75692 173216 75744
rect 164516 75624 164568 75676
rect 165528 75624 165580 75676
rect 167460 75624 167512 75676
rect 167736 75624 167788 75676
rect 169024 75624 169076 75676
rect 169484 75624 169536 75676
rect 169944 75624 169996 75676
rect 170128 75624 170180 75676
rect 145196 75556 145248 75608
rect 150440 75556 150492 75608
rect 150716 75556 150768 75608
rect 151084 75556 151136 75608
rect 153476 75556 153528 75608
rect 153752 75556 153804 75608
rect 153844 75556 153896 75608
rect 155132 75556 155184 75608
rect 155776 75556 155828 75608
rect 157340 75556 157392 75608
rect 157892 75556 157944 75608
rect 158444 75556 158496 75608
rect 159364 75556 159416 75608
rect 160284 75556 160336 75608
rect 160468 75556 160520 75608
rect 160652 75556 160704 75608
rect 242164 75556 242216 75608
rect 149152 75488 149204 75540
rect 149888 75488 149940 75540
rect 150532 75488 150584 75540
rect 150900 75488 150952 75540
rect 152924 75488 152976 75540
rect 154948 75488 155000 75540
rect 155684 75420 155736 75472
rect 156420 75420 156472 75472
rect 156604 75420 156656 75472
rect 156880 75420 156932 75472
rect 157432 75488 157484 75540
rect 157984 75488 158036 75540
rect 158720 75488 158772 75540
rect 162400 75488 162452 75540
rect 110420 75352 110472 75404
rect 133972 75352 134024 75404
rect 140412 75352 140464 75404
rect 148600 75352 148652 75404
rect 153292 75352 153344 75404
rect 153752 75352 153804 75404
rect 57244 75284 57296 75336
rect 127440 75284 127492 75336
rect 128728 75284 128780 75336
rect 129556 75284 129608 75336
rect 130108 75284 130160 75336
rect 130660 75284 130712 75336
rect 143724 75284 143776 75336
rect 144000 75284 144052 75336
rect 157616 75284 157668 75336
rect 157892 75284 157944 75336
rect 160284 75420 160336 75472
rect 160560 75420 160612 75472
rect 161296 75420 161348 75472
rect 162952 75420 163004 75472
rect 163964 75420 164016 75472
rect 164148 75420 164200 75472
rect 164608 75420 164660 75472
rect 174728 75488 174780 75540
rect 391204 75488 391256 75540
rect 471244 75420 471296 75472
rect 158536 75352 158588 75404
rect 161940 75352 161992 75404
rect 164240 75352 164292 75404
rect 164792 75352 164844 75404
rect 165436 75352 165488 75404
rect 478144 75352 478196 75404
rect 160560 75284 160612 75336
rect 161664 75284 161716 75336
rect 162216 75284 162268 75336
rect 163136 75284 163188 75336
rect 483020 75284 483072 75336
rect 46204 75216 46256 75268
rect 119804 75216 119856 75268
rect 129188 75216 129240 75268
rect 130200 75216 130252 75268
rect 139216 75216 139268 75268
rect 140412 75216 140464 75268
rect 140872 75216 140924 75268
rect 153108 75216 153160 75268
rect 154396 75216 154448 75268
rect 162400 75216 162452 75268
rect 162768 75216 162820 75268
rect 163964 75216 164016 75268
rect 168748 75216 168800 75268
rect 498200 75216 498252 75268
rect 22744 75148 22796 75200
rect 123760 75148 123812 75200
rect 135076 75148 135128 75200
rect 137744 75148 137796 75200
rect 152740 75148 152792 75200
rect 153844 75148 153896 75200
rect 154028 75148 154080 75200
rect 156696 75148 156748 75200
rect 126796 75080 126848 75132
rect 127440 75080 127492 75132
rect 128176 75080 128228 75132
rect 129372 75080 129424 75132
rect 133880 75080 133932 75132
rect 133972 75080 134024 75132
rect 136088 75080 136140 75132
rect 145012 75080 145064 75132
rect 145380 75080 145432 75132
rect 149612 75080 149664 75132
rect 149796 75080 149848 75132
rect 151820 75080 151872 75132
rect 154488 75080 154540 75132
rect 155224 75080 155276 75132
rect 157248 75080 157300 75132
rect 157616 75148 157668 75200
rect 158076 75148 158128 75200
rect 160376 75148 160428 75200
rect 160652 75148 160704 75200
rect 161112 75148 161164 75200
rect 164424 75080 164476 75132
rect 164884 75080 164936 75132
rect 165068 75080 165120 75132
rect 169392 75148 169444 75200
rect 532700 75148 532752 75200
rect 170404 75080 170456 75132
rect 125324 75012 125376 75064
rect 132960 75012 133012 75064
rect 133512 75012 133564 75064
rect 135536 75012 135588 75064
rect 135720 75012 135772 75064
rect 136548 75012 136600 75064
rect 123484 74944 123536 74996
rect 134892 74944 134944 74996
rect 135076 74944 135128 74996
rect 137008 75012 137060 75064
rect 147680 75012 147732 75064
rect 148140 75012 148192 75064
rect 150440 75012 150492 75064
rect 150992 75012 151044 75064
rect 158260 75012 158312 75064
rect 136732 74944 136784 74996
rect 137744 74944 137796 74996
rect 138664 74944 138716 74996
rect 139032 74944 139084 74996
rect 143816 74944 143868 74996
rect 144092 74944 144144 74996
rect 147956 74944 148008 74996
rect 155224 74944 155276 74996
rect 158904 74944 158956 74996
rect 159272 74944 159324 74996
rect 163228 74944 163280 74996
rect 163504 74944 163556 74996
rect 167552 75012 167604 75064
rect 173440 75012 173492 75064
rect 173348 74944 173400 74996
rect 127164 74876 127216 74928
rect 128084 74876 128136 74928
rect 128452 74876 128504 74928
rect 131488 74876 131540 74928
rect 135536 74876 135588 74928
rect 135904 74876 135956 74928
rect 138112 74876 138164 74928
rect 138756 74876 138808 74928
rect 139860 74876 139912 74928
rect 140044 74876 140096 74928
rect 144920 74876 144972 74928
rect 145472 74876 145524 74928
rect 147864 74876 147916 74928
rect 148140 74876 148192 74928
rect 125140 74808 125192 74860
rect 132316 74808 132368 74860
rect 134064 74808 134116 74860
rect 134524 74808 134576 74860
rect 135444 74808 135496 74860
rect 136180 74808 136232 74860
rect 136640 74808 136692 74860
rect 137008 74808 137060 74860
rect 140780 74808 140832 74860
rect 141424 74808 141476 74860
rect 145288 74808 145340 74860
rect 145748 74808 145800 74860
rect 129740 74740 129792 74792
rect 135628 74740 135680 74792
rect 135904 74740 135956 74792
rect 136456 74740 136508 74792
rect 145472 74740 145524 74792
rect 146024 74740 146076 74792
rect 160100 74876 160152 74928
rect 160560 74876 160612 74928
rect 161388 74876 161440 74928
rect 167552 74876 167604 74928
rect 167828 74876 167880 74928
rect 170128 74876 170180 74928
rect 170956 74876 171008 74928
rect 171784 74876 171836 74928
rect 183008 74876 183060 74928
rect 155224 74808 155276 74860
rect 162124 74808 162176 74860
rect 162860 74808 162912 74860
rect 163504 74808 163556 74860
rect 164424 74808 164476 74860
rect 172244 74808 172296 74860
rect 120724 74672 120776 74724
rect 128636 74672 128688 74724
rect 135260 74672 135312 74724
rect 136272 74672 136324 74724
rect 140872 74672 140924 74724
rect 158812 74740 158864 74792
rect 159548 74740 159600 74792
rect 160376 74740 160428 74792
rect 161020 74740 161072 74792
rect 165252 74740 165304 74792
rect 170496 74740 170548 74792
rect 171876 74740 171928 74792
rect 580724 74740 580776 74792
rect 154580 74672 154632 74724
rect 155224 74672 155276 74724
rect 164424 74672 164476 74724
rect 165160 74672 165212 74724
rect 165804 74672 165856 74724
rect 166264 74672 166316 74724
rect 170404 74672 170456 74724
rect 215944 74672 215996 74724
rect 124956 74468 125008 74520
rect 134800 74604 134852 74656
rect 135628 74604 135680 74656
rect 136364 74604 136416 74656
rect 162860 74604 162912 74656
rect 163688 74604 163740 74656
rect 165620 74604 165672 74656
rect 171508 74604 171560 74656
rect 131212 74536 131264 74588
rect 131856 74536 131908 74588
rect 168564 74536 168616 74588
rect 170772 74536 170824 74588
rect 122840 74400 122892 74452
rect 126796 74400 126848 74452
rect 171140 74468 171192 74520
rect 130292 74400 130344 74452
rect 131028 74400 131080 74452
rect 131120 74400 131172 74452
rect 167000 74400 167052 74452
rect 121000 74196 121052 74248
rect 128084 74332 128136 74384
rect 168288 74400 168340 74452
rect 169392 74400 169444 74452
rect 172980 74400 173032 74452
rect 168564 74332 168616 74384
rect 168932 74332 168984 74384
rect 169760 74332 169812 74384
rect 170404 74332 170456 74384
rect 102140 74128 102192 74180
rect 131856 74196 131908 74248
rect 132224 74196 132276 74248
rect 93860 74060 93912 74112
rect 128636 74060 128688 74112
rect 86960 73992 87012 74044
rect 131948 74128 132000 74180
rect 133052 74264 133104 74316
rect 133788 74264 133840 74316
rect 137100 74264 137152 74316
rect 137468 74264 137520 74316
rect 143816 74264 143868 74316
rect 144460 74264 144512 74316
rect 147680 74264 147732 74316
rect 148416 74264 148468 74316
rect 153108 74264 153160 74316
rect 197360 74264 197412 74316
rect 132776 74196 132828 74248
rect 133696 74196 133748 74248
rect 133972 74196 134024 74248
rect 134432 74196 134484 74248
rect 134616 74196 134668 74248
rect 135168 74196 135220 74248
rect 142252 74196 142304 74248
rect 142712 74196 142764 74248
rect 147496 74196 147548 74248
rect 226340 74196 226392 74248
rect 133420 74128 133472 74180
rect 139952 74128 140004 74180
rect 140320 74128 140372 74180
rect 144552 74128 144604 74180
rect 240140 74128 240192 74180
rect 131396 74060 131448 74112
rect 132408 74060 132460 74112
rect 132684 74060 132736 74112
rect 133604 74060 133656 74112
rect 138296 74060 138348 74112
rect 138664 74060 138716 74112
rect 142344 74060 142396 74112
rect 142712 74060 142764 74112
rect 145932 74060 145984 74112
rect 260840 74060 260892 74112
rect 131488 73992 131540 74044
rect 132132 73992 132184 74044
rect 138572 73992 138624 74044
rect 138848 73992 138900 74044
rect 139400 73992 139452 74044
rect 140228 73992 140280 74044
rect 160192 73992 160244 74044
rect 160836 73992 160888 74044
rect 69020 73924 69072 73976
rect 124772 73924 124824 73976
rect 134524 73924 134576 73976
rect 135352 73924 135404 73976
rect 136824 73924 136876 73976
rect 137836 73924 137888 73976
rect 146392 73924 146444 73976
rect 146668 73924 146720 73976
rect 44180 73856 44232 73908
rect 30380 73788 30432 73840
rect 122196 73856 122248 73908
rect 127532 73856 127584 73908
rect 143080 73856 143132 73908
rect 147496 73856 147548 73908
rect 159088 73856 159140 73908
rect 159272 73856 159324 73908
rect 128360 73788 128412 73840
rect 127992 73720 128044 73772
rect 143724 73720 143776 73772
rect 144368 73720 144420 73772
rect 151912 73720 151964 73772
rect 152648 73720 152700 73772
rect 155592 73720 155644 73772
rect 296720 73992 296772 74044
rect 120908 73652 120960 73704
rect 127072 73652 127124 73704
rect 136732 73652 136784 73704
rect 138940 73652 138992 73704
rect 161940 73652 161992 73704
rect 162308 73652 162360 73704
rect 165712 73652 165764 73704
rect 166264 73652 166316 73704
rect 120816 73584 120868 73636
rect 128084 73584 128136 73636
rect 157248 73584 157300 73636
rect 382280 73924 382332 73976
rect 166908 73856 166960 73908
rect 390560 73856 390612 73908
rect 168380 73788 168432 73840
rect 168932 73788 168984 73840
rect 169760 73788 169812 73840
rect 170680 73788 170732 73840
rect 166724 73720 166776 73772
rect 171876 73720 171928 73772
rect 169668 73652 169720 73704
rect 558920 73788 558972 73840
rect 168288 73584 168340 73636
rect 172704 73584 172756 73636
rect 125876 73516 125928 73568
rect 126336 73516 126388 73568
rect 127072 73516 127124 73568
rect 131120 73516 131172 73568
rect 165620 73516 165672 73568
rect 166632 73516 166684 73568
rect 136732 73448 136784 73500
rect 137284 73448 137336 73500
rect 139584 73448 139636 73500
rect 140136 73448 140188 73500
rect 152832 73448 152884 73500
rect 161020 73448 161072 73500
rect 161296 73448 161348 73500
rect 172428 73448 172480 73500
rect 146576 73380 146628 73432
rect 147220 73380 147272 73432
rect 149244 73380 149296 73432
rect 152648 73380 152700 73432
rect 166172 73380 166224 73432
rect 166816 73380 166868 73432
rect 127532 73312 127584 73364
rect 127900 73312 127952 73364
rect 152188 73312 152240 73364
rect 152556 73312 152608 73364
rect 163044 73312 163096 73364
rect 163780 73312 163832 73364
rect 137376 73244 137428 73296
rect 144460 73244 144512 73296
rect 149244 73244 149296 73296
rect 150072 73244 150124 73296
rect 132592 73176 132644 73228
rect 132960 73176 133012 73228
rect 128360 73108 128412 73160
rect 133512 73108 133564 73160
rect 431960 73108 432012 73160
rect 580172 73108 580224 73160
rect 140964 73040 141016 73092
rect 141516 73040 141568 73092
rect 132960 72972 133012 73024
rect 133328 72972 133380 73024
rect 121460 72836 121512 72888
rect 134984 72836 135036 72888
rect 107660 72768 107712 72820
rect 129372 72768 129424 72820
rect 162676 72768 162728 72820
rect 172060 72768 172112 72820
rect 51080 72700 51132 72752
rect 129464 72700 129516 72752
rect 159916 72700 159968 72752
rect 431960 72700 432012 72752
rect 60740 72632 60792 72684
rect 130752 72632 130804 72684
rect 152924 72632 152976 72684
rect 158352 72632 158404 72684
rect 163872 72632 163924 72684
rect 438860 72632 438912 72684
rect 42800 72564 42852 72616
rect 128912 72564 128964 72616
rect 150716 72564 150768 72616
rect 151268 72564 151320 72616
rect 161204 72564 161256 72616
rect 454040 72564 454092 72616
rect 16580 72496 16632 72548
rect 6920 72428 6972 72480
rect 121644 72428 121696 72480
rect 126336 72496 126388 72548
rect 126612 72496 126664 72548
rect 154948 72496 155000 72548
rect 155500 72496 155552 72548
rect 164056 72496 164108 72548
rect 489920 72496 489972 72548
rect 126888 72428 126940 72480
rect 128636 72428 128688 72480
rect 129648 72428 129700 72480
rect 138756 72428 138808 72480
rect 124220 72360 124272 72412
rect 125416 72360 125468 72412
rect 167828 72428 167880 72480
rect 535460 72428 535512 72480
rect 168656 72360 168708 72412
rect 169116 72360 169168 72412
rect 174268 72360 174320 72412
rect 174636 72360 174688 72412
rect 163780 72292 163832 72344
rect 168380 72292 168432 72344
rect 169208 72292 169260 72344
rect 168748 72224 168800 72276
rect 169116 72224 169168 72276
rect 151452 72088 151504 72140
rect 154212 72088 154264 72140
rect 168748 72088 168800 72140
rect 169300 72088 169352 72140
rect 159088 71952 159140 72004
rect 159456 71952 159508 72004
rect 154672 71816 154724 71868
rect 155408 71816 155460 71868
rect 163964 71748 164016 71800
rect 170680 71748 170732 71800
rect 3516 71680 3568 71732
rect 171784 71680 171836 71732
rect 137652 71612 137704 71664
rect 142988 71612 143040 71664
rect 149612 71544 149664 71596
rect 150256 71544 150308 71596
rect 171048 71544 171100 71596
rect 171784 71544 171836 71596
rect 140688 71408 140740 71460
rect 184940 71408 184992 71460
rect 118700 71340 118752 71392
rect 134064 71340 134116 71392
rect 154120 71340 154172 71392
rect 211804 71340 211856 71392
rect 93952 71272 94004 71324
rect 132592 71272 132644 71324
rect 141792 71272 141844 71324
rect 209780 71272 209832 71324
rect 75920 71204 75972 71256
rect 131212 71204 131264 71256
rect 142896 71204 142948 71256
rect 216680 71204 216732 71256
rect 64880 71136 64932 71188
rect 130844 71136 130896 71188
rect 143080 71136 143132 71188
rect 223580 71136 223632 71188
rect 46940 71068 46992 71120
rect 127624 71068 127676 71120
rect 147864 71068 147916 71120
rect 148232 71068 148284 71120
rect 161388 71068 161440 71120
rect 375380 71068 375432 71120
rect 26240 71000 26292 71052
rect 126612 71000 126664 71052
rect 169116 71000 169168 71052
rect 564440 71000 564492 71052
rect 141148 70864 141200 70916
rect 141700 70864 141752 70916
rect 142344 70864 142396 70916
rect 142804 70864 142856 70916
rect 146852 70728 146904 70780
rect 147128 70728 147180 70780
rect 148232 70728 148284 70780
rect 148508 70728 148560 70780
rect 150992 70456 151044 70508
rect 151360 70456 151412 70508
rect 151820 70456 151872 70508
rect 152464 70456 152516 70508
rect 152648 69980 152700 70032
rect 305000 69980 305052 70032
rect 149888 69912 149940 69964
rect 311900 69912 311952 69964
rect 151176 69844 151228 69896
rect 325700 69844 325752 69896
rect 154488 69776 154540 69828
rect 332600 69776 332652 69828
rect 154028 69708 154080 69760
rect 340880 69708 340932 69760
rect 114560 69640 114612 69692
rect 133972 69640 134024 69692
rect 138664 69640 138716 69692
rect 149980 69640 150032 69692
rect 156788 69640 156840 69692
rect 382372 69640 382424 69692
rect 149060 69572 149112 69624
rect 149796 69572 149848 69624
rect 138572 68960 138624 69012
rect 142804 68960 142856 69012
rect 148968 68552 149020 68604
rect 190460 68552 190512 68604
rect 163596 68484 163648 68536
rect 487160 68484 487212 68536
rect 165528 68416 165580 68468
rect 500960 68416 501012 68468
rect 164976 68348 165028 68400
rect 505100 68348 505152 68400
rect 169024 68280 169076 68332
rect 564532 68280 564584 68332
rect 140044 67192 140096 67244
rect 182180 67192 182232 67244
rect 141516 67124 141568 67176
rect 209872 67124 209924 67176
rect 156696 67056 156748 67108
rect 396080 67056 396132 67108
rect 166356 66988 166408 67040
rect 523040 66988 523092 67040
rect 167736 66920 167788 66972
rect 536840 66920 536892 66972
rect 170772 66852 170824 66904
rect 550640 66852 550692 66904
rect 142712 65832 142764 65884
rect 218060 65832 218112 65884
rect 154212 65764 154264 65816
rect 332692 65764 332744 65816
rect 157984 65696 158036 65748
rect 408500 65696 408552 65748
rect 167644 65628 167696 65680
rect 539600 65628 539652 65680
rect 167552 65560 167604 65612
rect 543740 65560 543792 65612
rect 170404 65492 170456 65544
rect 568580 65492 568632 65544
rect 139952 64540 140004 64592
rect 189080 64540 189132 64592
rect 141424 64472 141476 64524
rect 207020 64472 207072 64524
rect 145656 64404 145708 64456
rect 256700 64404 256752 64456
rect 147128 64336 147180 64388
rect 270500 64336 270552 64388
rect 151084 64268 151136 64320
rect 324320 64268 324372 64320
rect 162216 64200 162268 64252
rect 368480 64200 368532 64252
rect 159364 64132 159416 64184
rect 437480 64132 437532 64184
rect 139860 63112 139912 63164
rect 185032 63112 185084 63164
rect 145564 63044 145616 63096
rect 259460 63044 259512 63096
rect 161020 62976 161072 63028
rect 347780 62976 347832 63028
rect 152372 62908 152424 62960
rect 340972 62908 341024 62960
rect 155316 62840 155368 62892
rect 376760 62840 376812 62892
rect 157892 62772 157944 62824
rect 412640 62772 412692 62824
rect 138480 62160 138532 62212
rect 140044 62160 140096 62212
rect 137284 62092 137336 62144
rect 138664 62092 138716 62144
rect 144184 61820 144236 61872
rect 234620 61820 234672 61872
rect 144276 61752 144328 61804
rect 238760 61752 238812 61804
rect 147036 61684 147088 61736
rect 274640 61684 274692 61736
rect 150992 61616 151044 61668
rect 331220 61616 331272 61668
rect 153936 61548 153988 61600
rect 358820 61548 358872 61600
rect 159272 61480 159324 61532
rect 430580 61480 430632 61532
rect 166264 61412 166316 61464
rect 516140 61412 516192 61464
rect 170312 61344 170364 61396
rect 572720 61344 572772 61396
rect 118516 60664 118568 60716
rect 580172 60664 580224 60716
rect 142620 60256 142672 60308
rect 220820 60256 220872 60308
rect 148324 60188 148376 60240
rect 292580 60188 292632 60240
rect 149704 60120 149756 60172
rect 309140 60120 309192 60172
rect 153844 60052 153896 60104
rect 356060 60052 356112 60104
rect 157800 59984 157852 60036
rect 415400 59984 415452 60036
rect 162308 58760 162360 58812
rect 354680 58760 354732 58812
rect 160652 58692 160704 58744
rect 448520 58692 448572 58744
rect 163504 58624 163556 58676
rect 481640 58624 481692 58676
rect 137192 57876 137244 57928
rect 140136 57876 140188 57928
rect 155224 57332 155276 57384
rect 374000 57332 374052 57384
rect 164884 57264 164936 57316
rect 507860 57264 507912 57316
rect 166172 57196 166224 57248
rect 525800 57196 525852 57248
rect 95240 55836 95292 55888
rect 125324 55836 125376 55888
rect 152280 55836 152332 55888
rect 338120 55836 338172 55888
rect 148232 54544 148284 54596
rect 295340 54544 295392 54596
rect 102232 54476 102284 54528
rect 125232 54476 125284 54528
rect 156604 54476 156656 54528
rect 401600 54476 401652 54528
rect 149612 53048 149664 53100
rect 316040 53048 316092 53100
rect 156512 50464 156564 50516
rect 398840 50464 398892 50516
rect 161940 50396 161992 50448
rect 469220 50396 469272 50448
rect 163412 50328 163464 50380
rect 481732 50328 481784 50380
rect 182824 46860 182876 46912
rect 580172 46860 580224 46912
rect 139768 46180 139820 46232
rect 180800 46180 180852 46232
rect 3516 45500 3568 45552
rect 174636 45500 174688 45552
rect 35992 44820 36044 44872
rect 127440 44820 127492 44872
rect 171508 42032 171560 42084
rect 514852 42032 514904 42084
rect 120080 40264 120132 40316
rect 123484 40264 123536 40316
rect 88340 36524 88392 36576
rect 125140 36524 125192 36576
rect 145472 35572 145524 35624
rect 262220 35572 262272 35624
rect 146944 35504 146996 35556
rect 273260 35504 273312 35556
rect 146852 35436 146904 35488
rect 276020 35436 276072 35488
rect 148140 35368 148192 35420
rect 287060 35368 287112 35420
rect 149520 35300 149572 35352
rect 307760 35300 307812 35352
rect 155040 35232 155092 35284
rect 379520 35232 379572 35284
rect 155132 35164 155184 35216
rect 386420 35164 386472 35216
rect 141240 34144 141292 34196
rect 198740 34144 198792 34196
rect 142528 34076 142580 34128
rect 219440 34076 219492 34128
rect 144092 34008 144144 34060
rect 234712 34008 234764 34060
rect 145380 33940 145432 33992
rect 251180 33940 251232 33992
rect 145288 33872 145340 33924
rect 259552 33872 259604 33924
rect 141332 33804 141384 33856
rect 201500 33804 201552 33856
rect 215944 33804 215996 33856
rect 456800 33804 456852 33856
rect 170220 33736 170272 33788
rect 574100 33736 574152 33788
rect 170128 33056 170180 33108
rect 580172 33056 580224 33108
rect 3516 32988 3568 33040
rect 180892 32988 180944 33040
rect 174544 32580 174596 32632
rect 425060 32580 425112 32632
rect 163320 32512 163372 32564
rect 485780 32512 485832 32564
rect 167460 32444 167512 32496
rect 542360 32444 542412 32496
rect 170036 32376 170088 32428
rect 571340 32376 571392 32428
rect 149336 31492 149388 31544
rect 303620 31492 303672 31544
rect 149428 31424 149480 31476
rect 307852 31424 307904 31476
rect 150900 31356 150952 31408
rect 321560 31356 321612 31408
rect 154948 31288 155000 31340
rect 385040 31288 385092 31340
rect 159180 31220 159232 31272
rect 434720 31220 434772 31272
rect 164792 31152 164844 31204
rect 506480 31152 506532 31204
rect 166080 31084 166132 31136
rect 517520 31084 517572 31136
rect 165988 31016 166040 31068
rect 521660 31016 521712 31068
rect 144000 30064 144052 30116
rect 233240 30064 233292 30116
rect 143908 29996 143960 30048
rect 236000 29996 236052 30048
rect 145196 29928 145248 29980
rect 251272 29928 251324 29980
rect 146760 29860 146812 29912
rect 267832 29860 267884 29912
rect 147956 29792 148008 29844
rect 285680 29792 285732 29844
rect 148048 29724 148100 29776
rect 289820 29724 289872 29776
rect 154856 29656 154908 29708
rect 374092 29656 374144 29708
rect 161848 29588 161900 29640
rect 466460 29588 466512 29640
rect 141148 28704 141200 28756
rect 208400 28704 208452 28756
rect 142436 28636 142488 28688
rect 215300 28636 215352 28688
rect 142252 28568 142304 28620
rect 218152 28568 218204 28620
rect 142344 28500 142396 28552
rect 222200 28500 222252 28552
rect 143816 28432 143868 28484
rect 242900 28432 242952 28484
rect 145104 28364 145156 28416
rect 258080 28364 258132 28416
rect 161756 28296 161808 28348
rect 463700 28296 463752 28348
rect 165896 28228 165948 28280
rect 524420 28228 524472 28280
rect 141056 27276 141108 27328
rect 201592 27276 201644 27328
rect 140964 27208 141016 27260
rect 204260 27208 204312 27260
rect 145012 27140 145064 27192
rect 253940 27140 253992 27192
rect 146668 27072 146720 27124
rect 271880 27072 271932 27124
rect 153752 27004 153804 27056
rect 357440 27004 357492 27056
rect 160560 26936 160612 26988
rect 447140 26936 447192 26988
rect 161664 26868 161716 26920
rect 470600 26868 470652 26920
rect 140412 25984 140464 26036
rect 176752 25984 176804 26036
rect 139492 25916 139544 25968
rect 179420 25916 179472 25968
rect 139676 25848 139728 25900
rect 183560 25848 183612 25900
rect 139584 25780 139636 25832
rect 186320 25780 186372 25832
rect 146576 25712 146628 25764
rect 278780 25712 278832 25764
rect 152188 25644 152240 25696
rect 346400 25644 346452 25696
rect 164608 25576 164660 25628
rect 499580 25576 499632 25628
rect 164700 25508 164752 25560
rect 503720 25508 503772 25560
rect 139400 24488 139452 24540
rect 187700 24488 187752 24540
rect 150808 24420 150860 24472
rect 324412 24420 324464 24472
rect 171692 24352 171744 24404
rect 440240 24352 440292 24404
rect 168932 24284 168984 24336
rect 552020 24284 552072 24336
rect 168840 24216 168892 24268
rect 556160 24216 556212 24268
rect 168748 24148 168800 24200
rect 563060 24148 563112 24200
rect 169944 24080 169996 24132
rect 572812 24080 572864 24132
rect 3516 23196 3568 23248
rect 174360 23196 174412 23248
rect 150716 23128 150768 23180
rect 329840 23128 329892 23180
rect 157708 23060 157760 23112
rect 415492 23060 415544 23112
rect 167368 22992 167420 23044
rect 534080 22992 534132 23044
rect 167276 22924 167328 22976
rect 538220 22924 538272 22976
rect 167184 22856 167236 22908
rect 540980 22856 541032 22908
rect 52460 22788 52512 22840
rect 128728 22788 128780 22840
rect 169852 22788 169904 22840
rect 569960 22788 570012 22840
rect 118424 22720 118476 22772
rect 580172 22720 580224 22772
rect 158352 21768 158404 21820
rect 361580 21768 361632 21820
rect 173440 21700 173492 21752
rect 432052 21700 432104 21752
rect 158996 21632 159048 21684
rect 429200 21632 429252 21684
rect 159088 21564 159140 21616
rect 436100 21564 436152 21616
rect 165712 21496 165764 21548
rect 520280 21496 520332 21548
rect 165804 21428 165856 21480
rect 523132 21428 523184 21480
rect 45560 21360 45612 21412
rect 120816 21360 120868 21412
rect 165620 21360 165672 21412
rect 527180 21360 527232 21412
rect 135996 20612 136048 20664
rect 142252 20612 142304 20664
rect 144920 20340 144972 20392
rect 255320 20340 255372 20392
rect 146484 20272 146536 20324
rect 269120 20272 269172 20324
rect 143724 20204 143776 20256
rect 241520 20204 241572 20256
rect 242164 20204 242216 20256
rect 449900 20204 449952 20256
rect 173348 20136 173400 20188
rect 418160 20136 418212 20188
rect 163136 20068 163188 20120
rect 484400 20068 484452 20120
rect 106280 20000 106332 20052
rect 133052 20000 133104 20052
rect 163228 20000 163280 20052
rect 488540 20000 488592 20052
rect 70400 19932 70452 19984
rect 130292 19932 130344 19984
rect 164516 19932 164568 19984
rect 498292 19932 498344 19984
rect 150624 18912 150676 18964
rect 322940 18912 322992 18964
rect 172428 18844 172480 18896
rect 411260 18844 411312 18896
rect 161572 18776 161624 18828
rect 465172 18776 465224 18828
rect 168472 18708 168524 18760
rect 553400 18708 553452 18760
rect 168564 18640 168616 18692
rect 556252 18640 556304 18692
rect 4160 18572 4212 18624
rect 126152 18572 126204 18624
rect 168656 18572 168708 18624
rect 560300 18572 560352 18624
rect 140872 17620 140924 17672
rect 205640 17620 205692 17672
rect 158904 17552 158956 17604
rect 433340 17552 433392 17604
rect 158812 17484 158864 17536
rect 440332 17484 440384 17536
rect 160284 17416 160336 17468
rect 448612 17416 448664 17468
rect 160468 17348 160520 17400
rect 451280 17348 451332 17400
rect 160192 17280 160244 17332
rect 452660 17280 452712 17332
rect 38660 17212 38712 17264
rect 120724 17212 120776 17264
rect 160376 17212 160428 17264
rect 455420 17212 455472 17264
rect 147864 16124 147916 16176
rect 294880 16124 294932 16176
rect 154764 16056 154816 16108
rect 378416 16056 378468 16108
rect 156420 15988 156472 16040
rect 395344 15988 395396 16040
rect 157616 15920 157668 15972
rect 420184 15920 420236 15972
rect 14280 15852 14332 15904
rect 125048 15852 125100 15904
rect 164424 15852 164476 15904
rect 509608 15852 509660 15904
rect 143632 14696 143684 14748
rect 237656 14696 237708 14748
rect 152096 14628 152148 14680
rect 342904 14628 342956 14680
rect 154672 14560 154724 14612
rect 384304 14560 384356 14612
rect 172336 14492 172388 14544
rect 404360 14492 404412 14544
rect 31944 14424 31996 14476
rect 122196 14424 122248 14476
rect 156328 14424 156380 14476
rect 390652 14424 390704 14476
rect 147772 13540 147824 13592
rect 291384 13540 291436 13592
rect 152004 13472 152056 13524
rect 339500 13472 339552 13524
rect 153660 13404 153712 13456
rect 365720 13404 365772 13456
rect 154580 13336 154632 13388
rect 381176 13336 381228 13388
rect 156236 13268 156288 13320
rect 392584 13268 392636 13320
rect 156144 13200 156196 13252
rect 400864 13200 400916 13252
rect 157524 13132 157576 13184
rect 410800 13132 410852 13184
rect 164332 13064 164384 13116
rect 506572 13064 506624 13116
rect 151912 11908 151964 11960
rect 349252 11908 349304 11960
rect 153568 11840 153620 11892
rect 361120 11840 361172 11892
rect 153476 11772 153528 11824
rect 363512 11772 363564 11824
rect 117320 11704 117372 11756
rect 134156 11704 134208 11756
rect 153384 11704 153436 11756
rect 364616 11704 364668 11756
rect 176660 11636 176712 11688
rect 177856 11636 177908 11688
rect 201500 11636 201552 11688
rect 202696 11636 202748 11688
rect 234620 11636 234672 11688
rect 235816 11636 235868 11688
rect 259460 11636 259512 11688
rect 260656 11636 260708 11688
rect 149244 10684 149296 10736
rect 314660 10684 314712 10736
rect 99840 10616 99892 10668
rect 132960 10616 133012 10668
rect 150532 10616 150584 10668
rect 328000 10616 328052 10668
rect 81624 10548 81676 10600
rect 131764 10548 131816 10600
rect 151820 10548 151872 10600
rect 345296 10548 345348 10600
rect 78128 10480 78180 10532
rect 128452 10480 128504 10532
rect 172244 10480 172296 10532
rect 397736 10480 397788 10532
rect 67640 10412 67692 10464
rect 130200 10412 130252 10464
rect 158720 10412 158772 10464
rect 428464 10412 428516 10464
rect 64328 10344 64380 10396
rect 126336 10344 126388 10396
rect 164240 10344 164292 10396
rect 502984 10344 503036 10396
rect 25320 10276 25372 10328
rect 57244 10276 57296 10328
rect 60832 10276 60884 10328
rect 129096 10276 129148 10328
rect 167092 10276 167144 10328
rect 539692 10276 539744 10328
rect 116400 9256 116452 9308
rect 134708 9256 134760 9308
rect 53748 9188 53800 9240
rect 128636 9188 128688 9240
rect 138388 9188 138440 9240
rect 144920 9188 144972 9240
rect 149060 9188 149112 9240
rect 311440 9188 311492 9240
rect 50160 9120 50212 9172
rect 127624 9120 127676 9172
rect 149152 9120 149204 9172
rect 313832 9120 313884 9172
rect 34796 9052 34848 9104
rect 127348 9052 127400 9104
rect 153292 9052 153344 9104
rect 365812 9052 365864 9104
rect 9956 8984 10008 9036
rect 126060 8984 126112 9036
rect 157432 8984 157484 9036
rect 417884 8984 417936 9036
rect 572 8916 624 8968
rect 124220 8916 124272 8968
rect 163044 8916 163096 8968
rect 492312 8916 492364 8968
rect 105728 8032 105780 8084
rect 132776 8032 132828 8084
rect 104532 7964 104584 8016
rect 132684 7964 132736 8016
rect 98644 7896 98696 7948
rect 132868 7896 132920 7948
rect 84476 7828 84528 7880
rect 131488 7828 131540 7880
rect 80888 7760 80940 7812
rect 131672 7760 131724 7812
rect 143540 7760 143592 7812
rect 242992 7760 243044 7812
rect 77392 7692 77444 7744
rect 131580 7692 131632 7744
rect 146392 7692 146444 7744
rect 278320 7692 278372 7744
rect 6460 7624 6512 7676
rect 22744 7624 22796 7676
rect 27712 7624 27764 7676
rect 127256 7624 127308 7676
rect 147680 7624 147732 7676
rect 293684 7624 293736 7676
rect 18236 7556 18288 7608
rect 125968 7556 126020 7608
rect 161480 7556 161532 7608
rect 473452 7556 473504 7608
rect 555424 6808 555476 6860
rect 580172 6808 580224 6860
rect 140780 6604 140832 6656
rect 203892 6604 203944 6656
rect 142160 6536 142212 6588
rect 225144 6536 225196 6588
rect 66720 6468 66772 6520
rect 130108 6468 130160 6520
rect 146300 6468 146352 6520
rect 276020 6468 276072 6520
rect 391204 6468 391256 6520
rect 582196 6468 582248 6520
rect 63224 6400 63276 6452
rect 130016 6400 130068 6452
rect 155960 6400 156012 6452
rect 394240 6400 394292 6452
rect 48964 6332 49016 6384
rect 128544 6332 128596 6384
rect 156052 6332 156104 6384
rect 400128 6332 400180 6384
rect 44272 6264 44324 6316
rect 129280 6264 129332 6316
rect 160100 6264 160152 6316
rect 446220 6264 446272 6316
rect 33600 6196 33652 6248
rect 127164 6196 127216 6248
rect 162952 6196 163004 6248
rect 493508 6196 493560 6248
rect 24216 6128 24268 6180
rect 122104 6128 122156 6180
rect 168380 6128 168432 6180
rect 562048 6128 562100 6180
rect 101036 5380 101088 5432
rect 133144 5380 133196 5432
rect 97448 5312 97500 5364
rect 133328 5312 133380 5364
rect 136732 5312 136784 5364
rect 150624 5312 150676 5364
rect 85672 5244 85724 5296
rect 131396 5244 131448 5296
rect 138296 5244 138348 5296
rect 171968 5244 172020 5296
rect 15936 5176 15988 5228
rect 46204 5176 46256 5228
rect 59636 5176 59688 5228
rect 129924 5176 129976 5228
rect 151544 5176 151596 5228
rect 329196 5176 329248 5228
rect 30104 5108 30156 5160
rect 127532 5108 127584 5160
rect 136916 5108 136968 5160
rect 148324 5108 148376 5160
rect 153200 5108 153252 5160
rect 358728 5108 358780 5160
rect 28908 5040 28960 5092
rect 127808 5040 127860 5092
rect 137008 5040 137060 5092
rect 151820 5040 151872 5092
rect 157340 5040 157392 5092
rect 414296 5040 414348 5092
rect 19432 4972 19484 5024
rect 124864 4972 124916 5024
rect 138112 4972 138164 5024
rect 167184 4972 167236 5024
rect 170680 4972 170732 5024
rect 480536 4972 480588 5024
rect 13544 4904 13596 4956
rect 126520 4904 126572 4956
rect 137100 4904 137152 4956
rect 154212 4904 154264 4956
rect 162860 4904 162912 4956
rect 491116 4904 491168 4956
rect 11152 4836 11204 4888
rect 125876 4836 125928 4888
rect 8760 4768 8812 4820
rect 125784 4768 125836 4820
rect 136824 4700 136876 4752
rect 157800 4836 157852 4888
rect 168196 4836 168248 4888
rect 545488 4836 545540 4888
rect 138204 4768 138256 4820
rect 162492 4768 162544 4820
rect 169760 4768 169812 4820
rect 576308 4768 576360 4820
rect 135996 4156 136048 4208
rect 141240 4156 141292 4208
rect 119896 4088 119948 4140
rect 124956 4088 125008 4140
rect 125876 4088 125928 4140
rect 134524 4088 134576 4140
rect 137744 4088 137796 4140
rect 144736 4088 144788 4140
rect 138940 4020 138992 4072
rect 143540 4020 143592 4072
rect 12348 3952 12400 4004
rect 126428 3952 126480 4004
rect 138664 3952 138716 4004
rect 145932 3952 145984 4004
rect 144460 3884 144512 3936
rect 153016 3884 153068 3936
rect 86868 3816 86920 3868
rect 131856 3816 131908 3868
rect 135720 3816 135772 3868
rect 140044 3816 140096 3868
rect 140136 3816 140188 3868
rect 149520 3816 149572 3868
rect 211804 3816 211856 3868
rect 83280 3748 83332 3800
rect 79692 3680 79744 3732
rect 131304 3680 131356 3732
rect 131764 3748 131816 3800
rect 135812 3748 135864 3800
rect 142988 3748 143040 3800
rect 155408 3748 155460 3800
rect 172060 3748 172112 3800
rect 212172 3748 212224 3800
rect 242900 3816 242952 3868
rect 244096 3816 244148 3868
rect 251180 3816 251232 3868
rect 252376 3816 252428 3868
rect 284300 3816 284352 3868
rect 285036 3816 285088 3868
rect 344560 3748 344612 3800
rect 132040 3680 132092 3732
rect 135444 3680 135496 3732
rect 137652 3680 137704 3732
rect 144920 3680 144972 3732
rect 72608 3612 72660 3664
rect 126244 3612 126296 3664
rect 69112 3544 69164 3596
rect 130660 3612 130712 3664
rect 132960 3612 133012 3664
rect 135536 3612 135588 3664
rect 135628 3612 135680 3664
rect 138848 3612 138900 3664
rect 139952 3612 140004 3664
rect 149980 3680 150032 3732
rect 163688 3680 163740 3732
rect 171784 3680 171836 3732
rect 445024 3680 445076 3732
rect 126980 3544 127032 3596
rect 130384 3544 130436 3596
rect 135352 3544 135404 3596
rect 136456 3544 136508 3596
rect 142804 3544 142856 3596
rect 169576 3612 169628 3664
rect 171876 3612 171928 3664
rect 465172 3612 465224 3664
rect 23020 3476 23072 3528
rect 88156 3476 88208 3528
rect 93860 3476 93912 3528
rect 94780 3476 94832 3528
rect 110420 3476 110472 3528
rect 111616 3476 111668 3528
rect 124680 3476 124732 3528
rect 134616 3476 134668 3528
rect 135168 3476 135220 3528
rect 147128 3476 147180 3528
rect 166080 3544 166132 3596
rect 172152 3544 172204 3596
rect 468668 3544 468720 3596
rect 35900 3408 35952 3460
rect 36820 3408 36872 3460
rect 60740 3408 60792 3460
rect 61660 3408 61712 3460
rect 139032 3408 139084 3460
rect 163780 3476 163832 3528
rect 164884 3476 164936 3528
rect 172244 3476 172296 3528
rect 475752 3544 475804 3596
rect 471244 3476 471296 3528
rect 472256 3476 472308 3528
rect 506480 3476 506532 3528
rect 507308 3476 507360 3528
rect 539600 3476 539652 3528
rect 540428 3476 540480 3528
rect 173256 3408 173308 3460
rect 512460 3408 512512 3460
rect 170772 3340 170824 3392
rect 307760 3340 307812 3392
rect 309048 3340 309100 3392
rect 316040 3340 316092 3392
rect 317328 3340 317380 3392
rect 324412 3340 324464 3392
rect 325608 3340 325660 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 340972 3340 341024 3392
rect 342168 3340 342220 3392
rect 365720 3340 365772 3392
rect 367008 3340 367060 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 382372 3340 382424 3392
rect 383568 3340 383620 3392
rect 390652 3340 390704 3392
rect 391848 3340 391900 3392
rect 407120 3340 407172 3392
rect 408408 3340 408460 3392
rect 415400 3340 415452 3392
rect 416688 3340 416740 3392
rect 432052 3340 432104 3392
rect 433248 3340 433300 3392
rect 440332 3340 440384 3392
rect 441528 3340 441580 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 456800 3340 456852 3392
rect 458088 3340 458140 3392
rect 168380 3272 168432 3324
rect 152832 3136 152884 3188
rect 156604 3136 156656 3188
rect 478144 3136 478196 3188
rect 479340 3136 479392 3188
rect 173164 3068 173216 3120
rect 179052 3068 179104 3120
rect 349160 1368 349212 1420
rect 350448 1368 350500 1420
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 2778 671256 2834 671265
rect 2778 671191 2834 671200
rect 2792 670750 2820 671191
rect 2780 670744 2832 670750
rect 2780 670686 2832 670692
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3054 566944 3110 566953
rect 3054 566879 3110 566888
rect 3068 565894 3096 566879
rect 3056 565888 3108 565894
rect 3056 565830 3108 565836
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 2778 514856 2834 514865
rect 2778 514791 2780 514800
rect 2832 514791 2834 514800
rect 2780 514762 2832 514768
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3238 462632 3294 462641
rect 3238 462567 3240 462576
rect 3292 462567 3294 462576
rect 3240 462538 3292 462544
rect 3146 423600 3202 423609
rect 3146 423535 3202 423544
rect 3160 422958 3188 423535
rect 3148 422952 3200 422958
rect 3148 422894 3200 422900
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 409902 3188 410479
rect 3148 409896 3200 409902
rect 3148 409838 3200 409844
rect 3238 371376 3294 371385
rect 3238 371311 3294 371320
rect 3252 371278 3280 371311
rect 3240 371272 3292 371278
rect 3240 371214 3292 371220
rect 3238 358456 3294 358465
rect 3238 358391 3294 358400
rect 3252 357610 3280 358391
rect 3240 357604 3292 357610
rect 3240 357546 3292 357552
rect 3238 319288 3294 319297
rect 3238 319223 3294 319232
rect 3252 318850 3280 319223
rect 3240 318844 3292 318850
rect 3240 318786 3292 318792
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 2778 293176 2834 293185
rect 2778 293111 2834 293120
rect 2792 292874 2820 293111
rect 2780 292868 2832 292874
rect 2780 292810 2832 292816
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3160 253978 3188 254079
rect 3148 253972 3200 253978
rect 3148 253914 3200 253920
rect 2778 241088 2834 241097
rect 2778 241023 2834 241032
rect 2792 240242 2820 241023
rect 2780 240236 2832 240242
rect 2780 240178 2832 240184
rect 2962 201920 3018 201929
rect 2962 201855 3018 201864
rect 2976 201550 3004 201855
rect 2964 201544 3016 201550
rect 2964 201486 3016 201492
rect 3252 181490 3280 306167
rect 3344 231130 3372 475623
rect 3332 231124 3384 231130
rect 3332 231066 3384 231072
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3344 213994 3372 214911
rect 3332 213988 3384 213994
rect 3332 213930 3384 213936
rect 3330 188864 3386 188873
rect 3330 188799 3386 188808
rect 3344 187746 3372 188799
rect 3332 187740 3384 187746
rect 3332 187682 3384 187688
rect 3240 181484 3292 181490
rect 3240 181426 3292 181432
rect 3332 162920 3384 162926
rect 3330 162888 3332 162897
rect 3384 162888 3386 162897
rect 3330 162823 3386 162832
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3344 149122 3372 149767
rect 3332 149116 3384 149122
rect 3332 149058 3384 149064
rect 3436 138786 3464 684247
rect 6184 670744 6236 670750
rect 6184 670686 6236 670692
rect 3606 632088 3662 632097
rect 3606 632023 3662 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3424 138780 3476 138786
rect 3424 138722 3476 138728
rect 3422 136776 3478 136785
rect 3422 136711 3424 136720
rect 3476 136711 3478 136720
rect 3424 136682 3476 136688
rect 3424 133952 3476 133958
rect 3424 133894 3476 133900
rect 3332 131164 3384 131170
rect 3332 131106 3384 131112
rect 3240 111784 3292 111790
rect 3240 111726 3292 111732
rect 3252 110673 3280 111726
rect 3238 110664 3294 110673
rect 3238 110599 3294 110608
rect 3344 97617 3372 131106
rect 3330 97608 3386 97617
rect 3330 97543 3386 97552
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3160 84250 3188 84623
rect 3148 84244 3200 84250
rect 3148 84186 3200 84192
rect 1398 73808 1454 73817
rect 1398 73743 1454 73752
rect 572 8968 624 8974
rect 572 8910 624 8916
rect 584 480 612 8910
rect 542 -960 654 480
rect 1412 354 1440 73743
rect 2778 72448 2834 72457
rect 2778 72383 2834 72392
rect 2792 16574 2820 72383
rect 3436 19417 3464 133894
rect 3528 76537 3556 606047
rect 3620 138854 3648 632023
rect 3698 553888 3754 553897
rect 3698 553823 3754 553832
rect 3608 138848 3660 138854
rect 3608 138790 3660 138796
rect 3608 132524 3660 132530
rect 3608 132466 3660 132472
rect 3514 76528 3570 76537
rect 3514 76463 3570 76472
rect 3516 71732 3568 71738
rect 3516 71674 3568 71680
rect 3528 71641 3556 71674
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 3620 58585 3648 132466
rect 3712 78033 3740 553823
rect 4804 514820 4856 514826
rect 4804 514762 4856 514768
rect 3790 501800 3846 501809
rect 3790 501735 3846 501744
rect 3698 78024 3754 78033
rect 3698 77959 3754 77968
rect 3804 76673 3832 501735
rect 3882 449576 3938 449585
rect 3882 449511 3938 449520
rect 3896 78266 3924 449511
rect 3974 397488 4030 397497
rect 3974 397423 4030 397432
rect 3884 78260 3936 78266
rect 3884 78202 3936 78208
rect 3988 76945 4016 397423
rect 4066 345400 4122 345409
rect 4066 345335 4122 345344
rect 4080 84194 4108 345335
rect 4816 120086 4844 514762
rect 4896 292868 4948 292874
rect 4896 292810 4948 292816
rect 4804 120080 4856 120086
rect 4804 120022 4856 120028
rect 4080 84166 4200 84194
rect 4172 84130 4200 84166
rect 4080 84102 4200 84130
rect 4080 78402 4108 84102
rect 4908 78538 4936 292810
rect 4988 240236 5040 240242
rect 4988 240178 5040 240184
rect 4896 78532 4948 78538
rect 4896 78474 4948 78480
rect 4068 78396 4120 78402
rect 4068 78338 4120 78344
rect 3974 76936 4030 76945
rect 3974 76871 4030 76880
rect 3790 76664 3846 76673
rect 5000 76634 5028 240178
rect 6196 115938 6224 670686
rect 6276 422952 6328 422958
rect 6276 422894 6328 422900
rect 6288 142934 6316 422894
rect 6368 357604 6420 357610
rect 6368 357546 6420 357552
rect 6276 142928 6328 142934
rect 6276 142870 6328 142876
rect 6380 124166 6408 357546
rect 6368 124160 6420 124166
rect 6368 124102 6420 124108
rect 6184 115932 6236 115938
rect 6184 115874 6236 115880
rect 6932 78169 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 700330 24348 703520
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 33784 700324 33836 700330
rect 33784 700266 33836 700272
rect 15844 618316 15896 618322
rect 15844 618258 15896 618264
rect 8944 462596 8996 462602
rect 8944 462538 8996 462544
rect 8956 121446 8984 462538
rect 10324 409896 10376 409902
rect 10324 409838 10376 409844
rect 10336 122806 10364 409838
rect 10324 122800 10376 122806
rect 10324 122742 10376 122748
rect 8944 121440 8996 121446
rect 8944 121382 8996 121388
rect 15856 117298 15884 618258
rect 19984 579692 20036 579698
rect 19984 579634 20036 579640
rect 19996 141642 20024 579634
rect 20076 527196 20128 527202
rect 20076 527138 20128 527144
rect 20088 143002 20116 527138
rect 24124 371272 24176 371278
rect 24124 371214 24176 371220
rect 22744 253972 22796 253978
rect 22744 253914 22796 253920
rect 20076 142996 20128 143002
rect 20076 142938 20128 142944
rect 19984 141636 20036 141642
rect 19984 141578 20036 141584
rect 19984 136672 20036 136678
rect 19984 136614 20036 136620
rect 15844 117292 15896 117298
rect 15844 117234 15896 117240
rect 19996 111790 20024 136614
rect 22756 126954 22784 253914
rect 22836 201544 22888 201550
rect 22836 201486 22888 201492
rect 22848 128314 22876 201486
rect 24136 143070 24164 371214
rect 24216 318844 24268 318850
rect 24216 318786 24268 318792
rect 24228 163538 24256 318786
rect 24216 163532 24268 163538
rect 24216 163474 24268 163480
rect 24216 149116 24268 149122
rect 24216 149058 24268 149064
rect 24124 143064 24176 143070
rect 24124 143006 24176 143012
rect 24228 129742 24256 149058
rect 24216 129736 24268 129742
rect 24216 129678 24268 129684
rect 22836 128308 22888 128314
rect 22836 128250 22888 128256
rect 22744 126948 22796 126954
rect 22744 126890 22796 126896
rect 33796 113150 33824 700266
rect 40052 141710 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 43444 565888 43496 565894
rect 43444 565830 43496 565836
rect 40684 266416 40736 266422
rect 40684 266358 40736 266364
rect 40696 163606 40724 266358
rect 40684 163600 40736 163606
rect 40684 163542 40736 163548
rect 40040 141704 40092 141710
rect 40040 141646 40092 141652
rect 43456 118658 43484 565830
rect 64144 457496 64196 457502
rect 64144 457438 64196 457444
rect 64156 445058 64184 457438
rect 48412 445052 48464 445058
rect 48412 444994 48464 445000
rect 64144 445052 64196 445058
rect 64144 444994 64196 445000
rect 48424 442338 48452 444994
rect 46664 442332 46716 442338
rect 46664 442274 46716 442280
rect 48412 442332 48464 442338
rect 48412 442274 48464 442280
rect 46676 436898 46704 442274
rect 45008 436892 45060 436898
rect 45008 436834 45060 436840
rect 46664 436892 46716 436898
rect 46664 436834 46716 436840
rect 44916 240916 44968 240922
rect 44916 240858 44968 240864
rect 44824 239760 44876 239766
rect 44824 239702 44876 239708
rect 44836 231742 44864 239702
rect 44824 231736 44876 231742
rect 44824 231678 44876 231684
rect 44928 226302 44956 240858
rect 45020 229090 45048 436834
rect 69664 396772 69716 396778
rect 69664 396714 69716 396720
rect 69676 385014 69704 396714
rect 68284 385008 68336 385014
rect 68284 384950 68336 384956
rect 69664 385008 69716 385014
rect 69664 384950 69716 384956
rect 64236 380180 64288 380186
rect 64236 380122 64288 380128
rect 64144 358148 64196 358154
rect 64144 358090 64196 358096
rect 60188 356516 60240 356522
rect 60188 356458 60240 356464
rect 60200 354006 60228 356458
rect 49608 354000 49660 354006
rect 49608 353942 49660 353948
rect 60188 354000 60240 354006
rect 60188 353942 60240 353948
rect 49620 350606 49648 353942
rect 46204 350600 46256 350606
rect 46204 350542 46256 350548
rect 49608 350600 49660 350606
rect 49608 350542 49660 350548
rect 46216 342990 46244 350542
rect 45376 342984 45428 342990
rect 45376 342926 45428 342932
rect 46204 342984 46256 342990
rect 46204 342926 46256 342932
rect 45388 248414 45416 342926
rect 62856 331900 62908 331906
rect 62856 331842 62908 331848
rect 62764 319456 62816 319462
rect 62764 319398 62816 319404
rect 61476 318436 61528 318442
rect 61476 318378 61528 318384
rect 61488 311234 61516 318378
rect 60004 311228 60056 311234
rect 60004 311170 60056 311176
rect 61476 311228 61528 311234
rect 61476 311170 61528 311176
rect 60016 291174 60044 311170
rect 62776 299470 62804 319398
rect 62868 318442 62896 331842
rect 64156 319462 64184 358090
rect 64248 356522 64276 380122
rect 68296 358834 68324 384950
rect 65432 358828 65484 358834
rect 65432 358770 65484 358776
rect 68284 358828 68336 358834
rect 68284 358770 68336 358776
rect 65444 358154 65472 358770
rect 65432 358148 65484 358154
rect 65432 358090 65484 358096
rect 64236 356516 64288 356522
rect 64236 356458 64288 356464
rect 64144 319456 64196 319462
rect 64144 319398 64196 319404
rect 62856 318436 62908 318442
rect 62856 318378 62908 318384
rect 60832 299464 60884 299470
rect 60832 299406 60884 299412
rect 62764 299464 62816 299470
rect 62764 299406 62816 299412
rect 60844 294030 60872 299406
rect 60096 294024 60148 294030
rect 60096 293966 60148 293972
rect 60832 294024 60884 294030
rect 60832 293966 60884 293972
rect 58624 291168 58676 291174
rect 58624 291110 58676 291116
rect 60004 291168 60056 291174
rect 60004 291110 60056 291116
rect 57244 287700 57296 287706
rect 57244 287642 57296 287648
rect 56508 284300 56560 284306
rect 56508 284242 56560 284248
rect 56520 281178 56548 284242
rect 54300 281172 54352 281178
rect 54300 281114 54352 281120
rect 56508 281172 56560 281178
rect 56508 281114 56560 281120
rect 54312 278866 54340 281114
rect 53288 278860 53340 278866
rect 53288 278802 53340 278808
rect 54300 278860 54352 278866
rect 54300 278802 54352 278808
rect 54484 278860 54536 278866
rect 54484 278802 54536 278808
rect 53104 274712 53156 274718
rect 53104 274654 53156 274660
rect 51816 272128 51868 272134
rect 51816 272070 51868 272076
rect 51724 264920 51776 264926
rect 51724 264862 51776 264868
rect 49700 263628 49752 263634
rect 49700 263570 49752 263576
rect 49712 259010 49740 263570
rect 46940 259004 46992 259010
rect 46940 258946 46992 258952
rect 49700 259004 49752 259010
rect 49700 258946 49752 258952
rect 46952 255338 46980 258946
rect 50436 256692 50488 256698
rect 50436 256634 50488 256640
rect 45560 255332 45612 255338
rect 45560 255274 45612 255280
rect 46940 255332 46992 255338
rect 46940 255274 46992 255280
rect 45296 248386 45416 248414
rect 45192 245608 45244 245614
rect 45192 245550 45244 245556
rect 45100 240984 45152 240990
rect 45100 240926 45152 240932
rect 45112 231946 45140 240926
rect 45100 231940 45152 231946
rect 45100 231882 45152 231888
rect 45204 231062 45232 245550
rect 45296 231878 45324 248386
rect 45376 240848 45428 240854
rect 45376 240790 45428 240796
rect 45388 232014 45416 240790
rect 45468 238808 45520 238814
rect 45468 238750 45520 238756
rect 45480 232966 45508 238750
rect 45468 232960 45520 232966
rect 45468 232902 45520 232908
rect 45376 232008 45428 232014
rect 45376 231950 45428 231956
rect 45284 231872 45336 231878
rect 45284 231814 45336 231820
rect 45192 231056 45244 231062
rect 45192 230998 45244 231004
rect 45008 229084 45060 229090
rect 45008 229026 45060 229032
rect 44916 226296 44968 226302
rect 44916 226238 44968 226244
rect 45572 201482 45600 255274
rect 50448 253978 50476 256634
rect 47584 253972 47636 253978
rect 47584 253914 47636 253920
rect 50436 253972 50488 253978
rect 50436 253914 50488 253920
rect 46204 253904 46256 253910
rect 46204 253846 46256 253852
rect 45836 245676 45888 245682
rect 45836 245618 45888 245624
rect 45744 242888 45796 242894
rect 45744 242830 45796 242836
rect 45652 240440 45704 240446
rect 45652 240382 45704 240388
rect 45664 233034 45692 240382
rect 45756 233102 45784 242830
rect 45848 238814 45876 245618
rect 46216 245614 46244 253846
rect 47596 245682 47624 253914
rect 50344 250844 50396 250850
rect 50344 250786 50396 250792
rect 47584 245676 47636 245682
rect 47584 245618 47636 245624
rect 49700 245676 49752 245682
rect 49700 245618 49752 245624
rect 46204 245608 46256 245614
rect 46204 245550 46256 245556
rect 49712 242962 49740 245618
rect 49700 242956 49752 242962
rect 49700 242898 49752 242904
rect 46848 240780 46900 240786
rect 46848 240722 46900 240728
rect 46860 239766 46888 240722
rect 50356 240446 50384 250786
rect 51736 245682 51764 264862
rect 51828 263634 51856 272070
rect 51816 263628 51868 263634
rect 51816 263570 51868 263576
rect 53116 252618 53144 274654
rect 53300 272134 53328 278802
rect 53840 277364 53892 277370
rect 53840 277306 53892 277312
rect 53852 274718 53880 277306
rect 53840 274712 53892 274718
rect 53840 274654 53892 274660
rect 53288 272128 53340 272134
rect 53288 272070 53340 272076
rect 54496 266422 54524 278802
rect 57256 277438 57284 287642
rect 58636 284374 58664 291110
rect 58624 284368 58676 284374
rect 58624 284310 58676 284316
rect 60108 282946 60136 293966
rect 71792 287706 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 80704 491972 80756 491978
rect 80704 491914 80756 491920
rect 80716 478922 80744 491914
rect 77944 478916 77996 478922
rect 77944 478858 77996 478864
rect 80704 478916 80756 478922
rect 80704 478858 80756 478864
rect 77956 457502 77984 478858
rect 77944 457496 77996 457502
rect 77944 457438 77996 457444
rect 78588 382968 78640 382974
rect 78588 382910 78640 382916
rect 78600 380186 78628 382910
rect 78588 380180 78640 380186
rect 78588 380122 78640 380128
rect 88352 331906 88380 702406
rect 88984 504416 89036 504422
rect 88984 504358 89036 504364
rect 88996 491978 89024 504358
rect 88984 491972 89036 491978
rect 88984 491914 89036 491920
rect 104164 442944 104216 442950
rect 104164 442886 104216 442892
rect 95884 392624 95936 392630
rect 95884 392566 95936 392572
rect 95896 382974 95924 392566
rect 95884 382968 95936 382974
rect 95884 382910 95936 382916
rect 102784 381540 102836 381546
rect 102784 381482 102836 381488
rect 102140 379228 102192 379234
rect 102140 379170 102192 379176
rect 102152 375018 102180 379170
rect 101404 375012 101456 375018
rect 101404 374954 101456 374960
rect 102140 375012 102192 375018
rect 102140 374954 102192 374960
rect 95884 369912 95936 369918
rect 95884 369854 95936 369860
rect 95896 352442 95924 369854
rect 101416 362982 101444 374954
rect 102796 369918 102824 381482
rect 104176 379234 104204 442886
rect 104164 379228 104216 379234
rect 104164 379170 104216 379176
rect 102784 369912 102836 369918
rect 102784 369854 102836 369860
rect 100024 362976 100076 362982
rect 100024 362918 100076 362924
rect 101404 362976 101456 362982
rect 101404 362918 101456 362924
rect 93124 352436 93176 352442
rect 93124 352378 93176 352384
rect 95884 352436 95936 352442
rect 95884 352378 95936 352384
rect 88340 331900 88392 331906
rect 88340 331842 88392 331848
rect 91744 329452 91796 329458
rect 91744 329394 91796 329400
rect 84844 315308 84896 315314
rect 84844 315250 84896 315256
rect 71780 287700 71832 287706
rect 71780 287642 71832 287648
rect 84856 284374 84884 315250
rect 90364 298104 90416 298110
rect 90364 298046 90416 298052
rect 84844 284368 84896 284374
rect 84844 284310 84896 284316
rect 82084 284300 82136 284306
rect 82084 284242 82136 284248
rect 57980 282940 58032 282946
rect 57980 282882 58032 282888
rect 60096 282940 60148 282946
rect 60096 282882 60148 282888
rect 57992 280242 58020 282882
rect 60004 280832 60056 280838
rect 60004 280774 60056 280780
rect 57900 280214 58020 280242
rect 57900 278866 57928 280214
rect 57888 278860 57940 278866
rect 57888 278802 57940 278808
rect 57244 277432 57296 277438
rect 57244 277374 57296 277380
rect 55864 276684 55916 276690
rect 55864 276626 55916 276632
rect 55876 266422 55904 276626
rect 60016 268122 60044 280774
rect 82096 276690 82124 284242
rect 82084 276684 82136 276690
rect 82084 276626 82136 276632
rect 90376 270706 90404 298046
rect 86960 270700 87012 270706
rect 86960 270642 87012 270648
rect 90364 270700 90416 270706
rect 90364 270642 90416 270648
rect 86972 268394 87000 270642
rect 77944 268388 77996 268394
rect 77944 268330 77996 268336
rect 86960 268388 87012 268394
rect 86960 268330 87012 268336
rect 56600 268116 56652 268122
rect 56600 268058 56652 268064
rect 60004 268116 60056 268122
rect 60004 268058 60056 268064
rect 56612 267734 56640 268058
rect 56520 267706 56640 267734
rect 53196 266416 53248 266422
rect 53196 266358 53248 266364
rect 54484 266416 54536 266422
rect 54484 266358 54536 266364
rect 54576 266416 54628 266422
rect 54576 266358 54628 266364
rect 55864 266416 55916 266422
rect 55864 266358 55916 266364
rect 53208 254046 53236 266358
rect 54588 263634 54616 266358
rect 56520 264994 56548 267706
rect 56508 264988 56560 264994
rect 56508 264930 56560 264936
rect 53288 263628 53340 263634
rect 53288 263570 53340 263576
rect 54576 263628 54628 263634
rect 54576 263570 54628 263576
rect 53300 256766 53328 263570
rect 53288 256760 53340 256766
rect 53288 256702 53340 256708
rect 53196 254040 53248 254046
rect 53196 253982 53248 253988
rect 51816 252612 51868 252618
rect 51816 252554 51868 252560
rect 53104 252612 53156 252618
rect 53104 252554 53156 252560
rect 51828 250850 51856 252554
rect 51816 250844 51868 250850
rect 51816 250786 51868 250792
rect 77956 249762 77984 268330
rect 91756 249762 91784 329394
rect 93136 298110 93164 352378
rect 100036 332178 100064 362918
rect 94412 332172 94464 332178
rect 94412 332114 94464 332120
rect 100024 332172 100076 332178
rect 100024 332114 100076 332120
rect 94424 329458 94452 332114
rect 94412 329452 94464 329458
rect 94412 329394 94464 329400
rect 104912 315314 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 135996 676864 136048 676870
rect 135996 676806 136048 676812
rect 136008 674490 136036 676806
rect 133880 674484 133932 674490
rect 133880 674426 133932 674432
rect 135996 674484 136048 674490
rect 135996 674426 136048 674432
rect 133892 667554 133920 674426
rect 131764 667548 131816 667554
rect 131764 667490 131816 667496
rect 133880 667548 133932 667554
rect 133880 667490 133932 667496
rect 131776 662454 131804 667490
rect 127624 662448 127676 662454
rect 127624 662390 127676 662396
rect 131764 662448 131816 662454
rect 131764 662390 131816 662396
rect 127636 648650 127664 662390
rect 127624 648644 127676 648650
rect 127624 648586 127676 648592
rect 124864 648576 124916 648582
rect 124864 648518 124916 648524
rect 124876 603158 124904 648518
rect 124864 603152 124916 603158
rect 124864 603094 124916 603100
rect 121460 603084 121512 603090
rect 121460 603026 121512 603032
rect 121472 599622 121500 603026
rect 119988 599616 120040 599622
rect 119988 599558 120040 599564
rect 121460 599616 121512 599622
rect 121460 599558 121512 599564
rect 120000 597242 120028 599558
rect 117688 597236 117740 597242
rect 117688 597178 117740 597184
rect 119988 597236 120040 597242
rect 119988 597178 120040 597184
rect 117700 590646 117728 597178
rect 115204 590640 115256 590646
rect 115204 590582 115256 590588
rect 117688 590640 117740 590646
rect 117688 590582 117740 590588
rect 115216 580990 115244 590582
rect 112444 580984 112496 580990
rect 112444 580926 112496 580932
rect 115204 580984 115256 580990
rect 115204 580926 115256 580932
rect 112456 525842 112484 580926
rect 135904 580712 135956 580718
rect 135904 580654 135956 580660
rect 135916 572014 135944 580654
rect 126244 572008 126296 572014
rect 126244 571950 126296 571956
rect 135904 572008 135956 572014
rect 135904 571950 135956 571956
rect 126256 525842 126284 571950
rect 112444 525836 112496 525842
rect 112444 525778 112496 525784
rect 123484 525836 123536 525842
rect 123484 525778 123536 525784
rect 126244 525836 126296 525842
rect 126244 525778 126296 525784
rect 108948 525768 109000 525774
rect 108948 525710 109000 525716
rect 108960 522578 108988 525710
rect 106924 522572 106976 522578
rect 106924 522514 106976 522520
rect 108948 522572 109000 522578
rect 108948 522514 109000 522520
rect 106936 514826 106964 522514
rect 105544 514820 105596 514826
rect 105544 514762 105596 514768
rect 106924 514820 106976 514826
rect 106924 514762 106976 514768
rect 105556 442950 105584 514762
rect 123496 514078 123524 525778
rect 115204 514072 115256 514078
rect 115204 514014 115256 514020
rect 123484 514072 123536 514078
rect 123484 514014 123536 514020
rect 115216 504422 115244 514014
rect 115204 504416 115256 504422
rect 115204 504358 115256 504364
rect 128544 490612 128596 490618
rect 128544 490554 128596 490560
rect 128556 487558 128584 490554
rect 125692 487552 125744 487558
rect 125692 487494 125744 487500
rect 128544 487552 128596 487558
rect 128544 487494 128596 487500
rect 125704 485110 125732 487494
rect 120724 485104 120776 485110
rect 120724 485046 120776 485052
rect 125692 485104 125744 485110
rect 125692 485046 125744 485052
rect 120736 466138 120764 485046
rect 115572 466132 115624 466138
rect 115572 466074 115624 466080
rect 120724 466132 120776 466138
rect 120724 466074 120776 466080
rect 115584 462398 115612 466074
rect 109684 462392 109736 462398
rect 109684 462334 109736 462340
rect 115572 462392 115624 462398
rect 115572 462334 115624 462340
rect 105544 442944 105596 442950
rect 105544 442886 105596 442892
rect 109696 423638 109724 462334
rect 106924 423632 106976 423638
rect 106924 423574 106976 423580
rect 109684 423632 109736 423638
rect 109684 423574 109736 423580
rect 106936 392630 106964 423574
rect 136652 396778 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 696998 154160 703520
rect 170324 702434 170352 703520
rect 169772 702406 170352 702434
rect 152832 696992 152884 696998
rect 152832 696934 152884 696940
rect 154120 696992 154172 696998
rect 154120 696934 154172 696940
rect 152844 692850 152872 696934
rect 150440 692844 150492 692850
rect 150440 692786 150492 692792
rect 152832 692844 152884 692850
rect 152832 692786 152884 692792
rect 150452 688650 150480 692786
rect 150360 688622 150480 688650
rect 150360 687274 150388 688622
rect 150348 687268 150400 687274
rect 150348 687210 150400 687216
rect 146944 687200 146996 687206
rect 146944 687142 146996 687148
rect 146956 678298 146984 687142
rect 144920 678292 144972 678298
rect 144920 678234 144972 678240
rect 146944 678292 146996 678298
rect 146944 678234 146996 678240
rect 144932 676870 144960 678234
rect 144920 676864 144972 676870
rect 144920 676806 144972 676812
rect 163504 649324 163556 649330
rect 163504 649266 163556 649272
rect 163516 638518 163544 649266
rect 156604 638512 156656 638518
rect 156604 638454 156656 638460
rect 163504 638512 163556 638518
rect 163504 638454 163556 638460
rect 156616 622470 156644 638454
rect 152464 622464 152516 622470
rect 152464 622406 152516 622412
rect 156604 622464 156656 622470
rect 156604 622406 156656 622412
rect 152476 603770 152504 622406
rect 138664 603764 138716 603770
rect 138664 603706 138716 603712
rect 152464 603764 152516 603770
rect 152464 603706 152516 603712
rect 138676 580718 138704 603706
rect 138664 580712 138716 580718
rect 138664 580654 138716 580660
rect 157984 580304 158036 580310
rect 157984 580246 158036 580252
rect 157996 545766 158024 580246
rect 149704 545760 149756 545766
rect 149704 545702 149756 545708
rect 157984 545760 158036 545766
rect 157984 545702 158036 545708
rect 149716 496126 149744 545702
rect 138020 496120 138072 496126
rect 138020 496062 138072 496068
rect 149704 496120 149756 496126
rect 149704 496062 149756 496068
rect 138032 490618 138060 496062
rect 138020 490612 138072 490618
rect 138020 490554 138072 490560
rect 169024 429888 169076 429894
rect 169024 429830 169076 429836
rect 169036 407590 169064 429830
rect 166264 407584 166316 407590
rect 166264 407526 166316 407532
rect 169024 407584 169076 407590
rect 169024 407526 169076 407532
rect 136640 396772 136692 396778
rect 136640 396714 136692 396720
rect 106924 392624 106976 392630
rect 106924 392566 106976 392572
rect 166276 392018 166304 407526
rect 163504 392012 163556 392018
rect 163504 391954 163556 391960
rect 166264 392012 166316 392018
rect 166264 391954 166316 391960
rect 163516 381546 163544 391954
rect 163504 381540 163556 381546
rect 163504 381482 163556 381488
rect 104900 315308 104952 315314
rect 104900 315250 104952 315256
rect 169024 300280 169076 300286
rect 169024 300222 169076 300228
rect 93124 298104 93176 298110
rect 93124 298046 93176 298052
rect 169036 295390 169064 300222
rect 167644 295384 167696 295390
rect 167644 295326 167696 295332
rect 169024 295384 169076 295390
rect 169024 295326 169076 295332
rect 167656 278798 167684 295326
rect 169024 289128 169076 289134
rect 169024 289070 169076 289076
rect 167644 278792 167696 278798
rect 167644 278734 167696 278740
rect 162860 278724 162912 278730
rect 162860 278666 162912 278672
rect 162872 274718 162900 278666
rect 159364 274712 159416 274718
rect 159364 274654 159416 274660
rect 162860 274712 162912 274718
rect 162860 274654 162912 274660
rect 159376 262002 159404 274654
rect 169036 273290 169064 289070
rect 169772 280838 169800 702406
rect 202800 699718 202828 703520
rect 196624 699712 196676 699718
rect 196624 699654 196676 699660
rect 202788 699712 202840 699718
rect 202788 699654 202840 699660
rect 196636 692102 196664 699654
rect 185584 692096 185636 692102
rect 185584 692038 185636 692044
rect 196624 692096 196676 692102
rect 196624 692038 196676 692044
rect 185596 689314 185624 692038
rect 210424 690668 210476 690674
rect 210424 690610 210476 690616
rect 180064 689308 180116 689314
rect 180064 689250 180116 689256
rect 185584 689308 185636 689314
rect 185584 689250 185636 689256
rect 180076 666466 180104 689250
rect 210436 667214 210464 690610
rect 218072 680406 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 235184 699718 235212 703520
rect 229744 699712 229796 699718
rect 229744 699654 229796 699660
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 229756 690674 229784 699654
rect 267660 697338 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 260104 697332 260156 697338
rect 260104 697274 260156 697280
rect 267648 697332 267700 697338
rect 267648 697274 267700 697280
rect 229744 690668 229796 690674
rect 229744 690610 229796 690616
rect 217324 680400 217376 680406
rect 217324 680342 217376 680348
rect 218060 680400 218112 680406
rect 218060 680342 218112 680348
rect 202144 667208 202196 667214
rect 202144 667150 202196 667156
rect 210424 667208 210476 667214
rect 210424 667150 210476 667156
rect 177304 666460 177356 666466
rect 177304 666402 177356 666408
rect 180064 666460 180116 666466
rect 180064 666402 180116 666408
rect 177316 662454 177344 666402
rect 174544 662448 174596 662454
rect 174544 662390 174596 662396
rect 177304 662448 177356 662454
rect 177304 662390 177356 662396
rect 174556 651438 174584 662390
rect 171692 651432 171744 651438
rect 171692 651374 171744 651380
rect 174544 651432 174596 651438
rect 174544 651374 174596 651380
rect 171704 649330 171732 651374
rect 202156 650758 202184 667150
rect 217336 658850 217364 680342
rect 260116 678502 260144 697274
rect 253572 678496 253624 678502
rect 253572 678438 253624 678444
rect 260104 678496 260156 678502
rect 260104 678438 260156 678444
rect 253584 674082 253612 678438
rect 282932 677634 282960 702406
rect 300136 697746 300164 703520
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 300124 697740 300176 697746
rect 300124 697682 300176 697688
rect 307024 697740 307076 697746
rect 307024 697682 307076 697688
rect 307036 684486 307064 697682
rect 307024 684480 307076 684486
rect 307024 684422 307076 684428
rect 310244 684480 310296 684486
rect 310244 684422 310296 684428
rect 310256 678774 310284 684422
rect 310244 678768 310296 678774
rect 310244 678710 310296 678716
rect 315304 678768 315356 678774
rect 315304 678710 315356 678716
rect 282840 677606 282960 677634
rect 282840 674830 282868 677606
rect 278412 674824 278464 674830
rect 278412 674766 278464 674772
rect 282828 674824 282880 674830
rect 282828 674766 282880 674772
rect 250444 674076 250496 674082
rect 250444 674018 250496 674024
rect 253572 674076 253624 674082
rect 253572 674018 253624 674024
rect 250456 663814 250484 674018
rect 278424 669118 278452 674766
rect 276664 669112 276716 669118
rect 276664 669054 276716 669060
rect 278412 669112 278464 669118
rect 278412 669054 278464 669060
rect 247684 663808 247736 663814
rect 247684 663750 247736 663756
rect 250444 663808 250496 663814
rect 250444 663750 250496 663756
rect 214564 658844 214616 658850
rect 214564 658786 214616 658792
rect 217324 658844 217376 658850
rect 217324 658786 217376 658792
rect 195244 650752 195296 650758
rect 195244 650694 195296 650700
rect 202144 650752 202196 650758
rect 202144 650694 202196 650700
rect 171692 649324 171744 649330
rect 171692 649266 171744 649272
rect 195256 623082 195284 650694
rect 186964 623076 187016 623082
rect 186964 623018 187016 623024
rect 195244 623076 195296 623082
rect 195244 623018 195296 623024
rect 186976 612814 187004 623018
rect 184204 612808 184256 612814
rect 184204 612750 184256 612756
rect 186964 612808 187016 612814
rect 186964 612750 187016 612756
rect 184216 603770 184244 612750
rect 214576 609754 214604 658786
rect 247696 645862 247724 663750
rect 276676 661094 276704 669054
rect 273904 661088 273956 661094
rect 273904 661030 273956 661036
rect 276664 661088 276716 661094
rect 276664 661030 276716 661036
rect 273916 650078 273944 661030
rect 315316 653410 315344 678710
rect 331232 674830 331260 702986
rect 348804 702434 348832 703520
rect 347792 702406 348832 702434
rect 347792 688498 347820 702406
rect 364996 699718 365024 703520
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 369124 699712 369176 699718
rect 369124 699654 369176 699660
rect 369136 688634 369164 699654
rect 369124 688628 369176 688634
rect 369124 688570 369176 688576
rect 374644 688628 374696 688634
rect 374644 688570 374696 688576
rect 347780 688492 347832 688498
rect 347780 688434 347832 688440
rect 351920 688492 351972 688498
rect 351920 688434 351972 688440
rect 351932 683806 351960 688434
rect 351920 683800 351972 683806
rect 351920 683742 351972 683748
rect 362224 683800 362276 683806
rect 362224 683742 362276 683748
rect 362236 681018 362264 683742
rect 374656 682310 374684 688570
rect 374644 682304 374696 682310
rect 374644 682246 374696 682252
rect 380256 682304 380308 682310
rect 380256 682246 380308 682252
rect 362224 681012 362276 681018
rect 362224 680954 362276 680960
rect 371240 681012 371292 681018
rect 371240 680954 371292 680960
rect 371252 675510 371280 680954
rect 380268 675510 380296 682246
rect 371240 675504 371292 675510
rect 371240 675446 371292 675452
rect 380164 675504 380216 675510
rect 380164 675446 380216 675452
rect 380256 675504 380308 675510
rect 380256 675446 380308 675452
rect 396448 675504 396500 675510
rect 396448 675446 396500 675452
rect 331220 674824 331272 674830
rect 331220 674766 331272 674772
rect 334624 674824 334676 674830
rect 334624 674766 334676 674772
rect 334636 663066 334664 674766
rect 334624 663060 334676 663066
rect 334624 663002 334676 663008
rect 358084 663060 358136 663066
rect 358084 663002 358136 663008
rect 315304 653404 315356 653410
rect 315304 653346 315356 653352
rect 319812 653404 319864 653410
rect 319812 653346 319864 653352
rect 273904 650072 273956 650078
rect 273904 650014 273956 650020
rect 269764 650004 269816 650010
rect 269764 649946 269816 649952
rect 269776 647970 269804 649946
rect 319824 648922 319852 653346
rect 358096 650010 358124 663002
rect 358084 650004 358136 650010
rect 358084 649946 358136 649952
rect 366364 650004 366416 650010
rect 366364 649946 366416 649952
rect 319812 648916 319864 648922
rect 319812 648858 319864 648864
rect 324964 648916 325016 648922
rect 324964 648858 325016 648864
rect 265624 647964 265676 647970
rect 265624 647906 265676 647912
rect 269764 647964 269816 647970
rect 269764 647906 269816 647912
rect 244924 645856 244976 645862
rect 244924 645798 244976 645804
rect 247684 645856 247736 645862
rect 247684 645798 247736 645804
rect 211804 609748 211856 609754
rect 211804 609690 211856 609696
rect 214564 609748 214616 609754
rect 214564 609690 214616 609696
rect 178040 603764 178092 603770
rect 178040 603706 178092 603712
rect 184204 603764 184256 603770
rect 184204 603706 184256 603712
rect 178052 600370 178080 603706
rect 171784 600364 171836 600370
rect 171784 600306 171836 600312
rect 178040 600364 178092 600370
rect 178040 600306 178092 600312
rect 171796 580310 171824 600306
rect 211816 592074 211844 609690
rect 210424 592068 210476 592074
rect 210424 592010 210476 592016
rect 211804 592068 211856 592074
rect 211804 592010 211856 592016
rect 171784 580304 171836 580310
rect 171784 580246 171836 580252
rect 209044 558204 209096 558210
rect 209044 558146 209096 558152
rect 207664 554464 207716 554470
rect 207664 554406 207716 554412
rect 207676 543794 207704 554406
rect 206284 543788 206336 543794
rect 206284 543730 206336 543736
rect 207664 543788 207716 543794
rect 207664 543730 207716 543736
rect 204904 536852 204956 536858
rect 204904 536794 204956 536800
rect 203524 511964 203576 511970
rect 203524 511906 203576 511912
rect 201868 507884 201920 507890
rect 201868 507826 201920 507832
rect 201880 500274 201908 507826
rect 189724 500268 189776 500274
rect 189724 500210 189776 500216
rect 201868 500268 201920 500274
rect 201868 500210 201920 500216
rect 189736 438938 189764 500210
rect 203536 445874 203564 511906
rect 204916 507890 204944 536794
rect 206296 511970 206324 543730
rect 209056 536858 209084 558146
rect 210436 554470 210464 592010
rect 244936 581194 244964 645798
rect 265636 598806 265664 647906
rect 324976 640286 325004 648858
rect 366376 647222 366404 649946
rect 380176 649330 380204 675446
rect 380164 649324 380216 649330
rect 380164 649266 380216 649272
rect 387064 649324 387116 649330
rect 387064 649266 387116 649272
rect 366364 647216 366416 647222
rect 366364 647158 366416 647164
rect 371884 647216 371936 647222
rect 371884 647158 371936 647164
rect 324964 640280 325016 640286
rect 324964 640222 325016 640228
rect 327724 640280 327776 640286
rect 327724 640222 327776 640228
rect 327736 632534 327764 640222
rect 371896 635526 371924 647158
rect 387076 643793 387104 649266
rect 387062 643784 387118 643793
rect 387062 643719 387118 643728
rect 371884 635520 371936 635526
rect 371884 635462 371936 635468
rect 388904 635520 388956 635526
rect 388904 635462 388956 635468
rect 327724 632528 327776 632534
rect 327724 632470 327776 632476
rect 329932 632528 329984 632534
rect 329932 632470 329984 632476
rect 329944 629950 329972 632470
rect 388916 631718 388944 635462
rect 388904 631712 388956 631718
rect 388904 631654 388956 631660
rect 395344 631712 395396 631718
rect 395344 631654 395396 631660
rect 329932 629944 329984 629950
rect 329932 629886 329984 629892
rect 339500 629944 339552 629950
rect 339500 629886 339552 629892
rect 339512 626550 339540 629886
rect 339500 626544 339552 626550
rect 339500 626486 339552 626492
rect 344008 626544 344060 626550
rect 344008 626486 344060 626492
rect 344020 620294 344048 626486
rect 344008 620288 344060 620294
rect 344008 620230 344060 620236
rect 353300 620288 353352 620294
rect 353300 620230 353352 620236
rect 353312 617574 353340 620230
rect 353300 617568 353352 617574
rect 353300 617510 353352 617516
rect 263600 598800 263652 598806
rect 263600 598742 263652 598748
rect 265624 598800 265676 598806
rect 265624 598742 265676 598748
rect 263612 595474 263640 598742
rect 249064 595468 249116 595474
rect 249064 595410 249116 595416
rect 263600 595468 263652 595474
rect 263600 595410 263652 595416
rect 241612 581188 241664 581194
rect 241612 581130 241664 581136
rect 244924 581188 244976 581194
rect 244924 581130 244976 581136
rect 241624 577658 241652 581130
rect 238760 577652 238812 577658
rect 238760 577594 238812 577600
rect 241612 577652 241664 577658
rect 241612 577594 241664 577600
rect 238772 574122 238800 577594
rect 236644 574116 236696 574122
rect 236644 574058 236696 574064
rect 238760 574116 238812 574122
rect 238760 574058 238812 574064
rect 236656 562154 236684 574058
rect 233240 562148 233292 562154
rect 233240 562090 233292 562096
rect 236644 562148 236696 562154
rect 236644 562090 236696 562096
rect 233252 558210 233280 562090
rect 233240 558204 233292 558210
rect 233240 558146 233292 558152
rect 210424 554464 210476 554470
rect 210424 554406 210476 554412
rect 209044 536852 209096 536858
rect 209044 536794 209096 536800
rect 206284 511964 206336 511970
rect 206284 511906 206336 511912
rect 204904 507884 204956 507890
rect 204904 507826 204956 507832
rect 249076 497486 249104 595410
rect 236644 497480 236696 497486
rect 236644 497422 236696 497428
rect 249064 497480 249116 497486
rect 249064 497422 249116 497428
rect 236656 474706 236684 497422
rect 235264 474700 235316 474706
rect 235264 474642 235316 474648
rect 236644 474700 236696 474706
rect 236644 474642 236696 474648
rect 235276 466478 235304 474642
rect 232504 466472 232556 466478
rect 232504 466414 232556 466420
rect 235264 466472 235316 466478
rect 235264 466414 235316 466420
rect 232516 446418 232544 466414
rect 226432 446412 226484 446418
rect 226432 446354 226484 446360
rect 232504 446412 232556 446418
rect 232504 446354 232556 446360
rect 201592 445868 201644 445874
rect 201592 445810 201644 445816
rect 203524 445868 203576 445874
rect 203524 445810 203576 445816
rect 201604 445398 201632 445810
rect 199384 445392 199436 445398
rect 199384 445334 199436 445340
rect 201592 445392 201644 445398
rect 201592 445334 201644 445340
rect 184204 438932 184256 438938
rect 184204 438874 184256 438880
rect 189724 438932 189776 438938
rect 189724 438874 189776 438880
rect 184216 435402 184244 438874
rect 199396 437510 199424 445334
rect 226444 442474 226472 446354
rect 225604 442468 225656 442474
rect 225604 442410 225656 442416
rect 226432 442468 226484 442474
rect 226432 442410 226484 442416
rect 199384 437504 199436 437510
rect 199384 437446 199436 437452
rect 196624 437436 196676 437442
rect 196624 437378 196676 437384
rect 174544 435396 174596 435402
rect 174544 435338 174596 435344
rect 184204 435396 184256 435402
rect 184204 435338 184256 435344
rect 174556 429894 174584 435338
rect 174544 429888 174596 429894
rect 174544 429830 174596 429836
rect 196636 426902 196664 437378
rect 193864 426896 193916 426902
rect 193864 426838 193916 426844
rect 196624 426896 196676 426902
rect 196624 426838 196676 426844
rect 193876 404394 193904 426838
rect 225616 407386 225644 442410
rect 224224 407380 224276 407386
rect 224224 407322 224276 407328
rect 225604 407380 225656 407386
rect 225604 407322 225656 407328
rect 193864 404388 193916 404394
rect 193864 404330 193916 404336
rect 191104 404320 191156 404326
rect 191104 404262 191156 404268
rect 191116 385082 191144 404262
rect 224236 396030 224264 407322
rect 223028 396024 223080 396030
rect 223028 395966 223080 395972
rect 224224 396024 224276 396030
rect 224224 395966 224276 395972
rect 223040 387122 223068 395966
rect 209044 387116 209096 387122
rect 209044 387058 209096 387064
rect 223028 387116 223080 387122
rect 223028 387058 223080 387064
rect 191104 385076 191156 385082
rect 191104 385018 191156 385024
rect 186964 385008 187016 385014
rect 186964 384950 187016 384956
rect 186976 350606 187004 384950
rect 209056 382294 209084 387058
rect 205640 382288 205692 382294
rect 205640 382230 205692 382236
rect 209044 382288 209096 382294
rect 209044 382230 209096 382236
rect 205652 378146 205680 382230
rect 202144 378140 202196 378146
rect 202144 378082 202196 378088
rect 205640 378140 205692 378146
rect 205640 378082 205692 378088
rect 202156 372638 202184 378082
rect 202144 372632 202196 372638
rect 202144 372574 202196 372580
rect 198004 372564 198056 372570
rect 198004 372506 198056 372512
rect 185584 350600 185636 350606
rect 185584 350542 185636 350548
rect 186964 350600 187016 350606
rect 186964 350542 187016 350548
rect 185596 338774 185624 350542
rect 198016 346390 198044 372506
rect 195244 346384 195296 346390
rect 195244 346326 195296 346332
rect 198004 346384 198056 346390
rect 198004 346326 198056 346332
rect 184204 338768 184256 338774
rect 184204 338710 184256 338716
rect 185584 338768 185636 338774
rect 185584 338710 185636 338716
rect 184216 329186 184244 338710
rect 182824 329180 182876 329186
rect 182824 329122 182876 329128
rect 184204 329180 184256 329186
rect 184204 329122 184256 329128
rect 181444 320204 181496 320210
rect 181444 320146 181496 320152
rect 181456 314702 181484 320146
rect 179512 314696 179564 314702
rect 179512 314638 179564 314644
rect 181444 314696 181496 314702
rect 181444 314638 181496 314644
rect 179524 309602 179552 314638
rect 178684 309596 178736 309602
rect 178684 309538 178736 309544
rect 179512 309596 179564 309602
rect 179512 309538 179564 309544
rect 178696 305250 178724 309538
rect 176660 305244 176712 305250
rect 176660 305186 176712 305192
rect 178684 305244 178736 305250
rect 178684 305186 178736 305192
rect 176672 304298 176700 305186
rect 170128 304292 170180 304298
rect 170128 304234 170180 304240
rect 176660 304292 176712 304298
rect 176660 304234 176712 304240
rect 170140 300286 170168 304234
rect 182836 302122 182864 329122
rect 195256 328098 195284 346326
rect 194048 328092 194100 328098
rect 194048 328034 194100 328040
rect 195244 328092 195296 328098
rect 195244 328034 195296 328040
rect 194060 322250 194088 328034
rect 183376 322244 183428 322250
rect 183376 322186 183428 322192
rect 194048 322244 194100 322250
rect 194048 322186 194100 322192
rect 183388 320210 183416 322186
rect 183376 320204 183428 320210
rect 183376 320146 183428 320152
rect 180064 302116 180116 302122
rect 180064 302058 180116 302064
rect 182824 302116 182876 302122
rect 182824 302058 182876 302064
rect 170128 300280 170180 300286
rect 170128 300222 170180 300228
rect 180076 291038 180104 302058
rect 175648 291032 175700 291038
rect 175648 290974 175700 290980
rect 180064 291032 180116 291038
rect 180064 290974 180116 290980
rect 175660 289134 175688 290974
rect 175648 289128 175700 289134
rect 175648 289070 175700 289076
rect 169760 280832 169812 280838
rect 169760 280774 169812 280780
rect 169024 273284 169076 273290
rect 169024 273226 169076 273232
rect 166264 273216 166316 273222
rect 166264 273158 166316 273164
rect 166276 264994 166304 273158
rect 164240 264988 164292 264994
rect 164240 264930 164292 264936
rect 166264 264988 166316 264994
rect 166264 264930 166316 264936
rect 156604 261996 156656 262002
rect 156604 261938 156656 261944
rect 159364 261996 159416 262002
rect 159364 261938 159416 261944
rect 156616 256766 156644 261938
rect 164252 260098 164280 264930
rect 162124 260092 162176 260098
rect 162124 260034 162176 260040
rect 164240 260092 164292 260098
rect 164240 260034 164292 260040
rect 154028 256760 154080 256766
rect 154028 256702 154080 256708
rect 156604 256760 156656 256766
rect 156604 256702 156656 256708
rect 154040 255338 154068 256702
rect 151084 255332 151136 255338
rect 151084 255274 151136 255280
rect 154028 255332 154080 255338
rect 154028 255274 154080 255280
rect 75184 249756 75236 249762
rect 75184 249698 75236 249704
rect 77944 249756 77996 249762
rect 77944 249698 77996 249704
rect 89168 249756 89220 249762
rect 89168 249698 89220 249704
rect 91744 249756 91796 249762
rect 91744 249698 91796 249704
rect 51724 245676 51776 245682
rect 51724 245618 51776 245624
rect 75092 243024 75144 243030
rect 75092 242966 75144 242972
rect 75104 240990 75132 242966
rect 75092 240984 75144 240990
rect 75092 240926 75144 240932
rect 75196 240922 75224 249698
rect 89180 244934 89208 249698
rect 151096 245682 151124 255274
rect 162136 245954 162164 260034
rect 160100 245948 160152 245954
rect 160100 245890 160152 245896
rect 162124 245948 162176 245954
rect 162124 245890 162176 245896
rect 145196 245676 145248 245682
rect 145196 245618 145248 245624
rect 151084 245676 151136 245682
rect 151084 245618 151136 245624
rect 81440 244928 81492 244934
rect 81440 244870 81492 244876
rect 89168 244928 89220 244934
rect 89168 244870 89220 244876
rect 81452 243030 81480 244870
rect 81440 243024 81492 243030
rect 81440 242966 81492 242972
rect 145208 241874 145236 245618
rect 142988 241868 143040 241874
rect 142988 241810 143040 241816
rect 145196 241868 145248 241874
rect 145196 241810 145248 241816
rect 75184 240916 75236 240922
rect 75184 240858 75236 240864
rect 143000 240854 143028 241810
rect 142988 240848 143040 240854
rect 142988 240790 143040 240796
rect 160112 240786 160140 245890
rect 160100 240780 160152 240786
rect 160100 240722 160152 240728
rect 50344 240440 50396 240446
rect 50344 240382 50396 240388
rect 395356 240038 395384 631654
rect 395436 617568 395488 617574
rect 395436 617510 395488 617516
rect 395344 240032 395396 240038
rect 395344 239974 395396 239980
rect 395448 239834 395476 617510
rect 395436 239828 395488 239834
rect 395436 239770 395488 239776
rect 46848 239760 46900 239766
rect 46848 239702 46900 239708
rect 45836 238808 45888 238814
rect 45836 238750 45888 238756
rect 45744 233096 45796 233102
rect 45744 233038 45796 233044
rect 45652 233028 45704 233034
rect 45652 232970 45704 232976
rect 45836 232960 45888 232966
rect 45836 232902 45888 232908
rect 45848 231198 45876 232902
rect 62764 232416 62816 232422
rect 62764 232358 62816 232364
rect 80704 232416 80756 232422
rect 80704 232358 80756 232364
rect 395436 232416 395488 232422
rect 395436 232358 395488 232364
rect 46572 232008 46624 232014
rect 46572 231950 46624 231956
rect 45836 231192 45888 231198
rect 45836 231134 45888 231140
rect 46584 230518 46612 231950
rect 46848 231872 46900 231878
rect 46848 231814 46900 231820
rect 46572 230512 46624 230518
rect 46572 230454 46624 230460
rect 46860 227610 46888 231814
rect 49148 231804 49200 231810
rect 49148 231746 49200 231752
rect 47032 229084 47084 229090
rect 47032 229026 47084 229032
rect 46860 227582 46980 227610
rect 46952 225010 46980 227582
rect 47044 225758 47072 229026
rect 47032 225752 47084 225758
rect 47032 225694 47084 225700
rect 46940 225004 46992 225010
rect 46940 224946 46992 224952
rect 49160 222222 49188 231746
rect 49792 231736 49844 231742
rect 49792 231678 49844 231684
rect 49700 230444 49752 230450
rect 49700 230386 49752 230392
rect 49712 226370 49740 230386
rect 49804 230178 49832 231678
rect 49792 230172 49844 230178
rect 49792 230114 49844 230120
rect 55128 230172 55180 230178
rect 55128 230114 55180 230120
rect 49700 226364 49752 226370
rect 49700 226306 49752 226312
rect 50436 226296 50488 226302
rect 50436 226238 50488 226244
rect 55140 226250 55168 230114
rect 56232 226296 56284 226302
rect 50344 224936 50396 224942
rect 50344 224878 50396 224884
rect 49148 222216 49200 222222
rect 49148 222158 49200 222164
rect 50356 213926 50384 224878
rect 50448 215150 50476 226238
rect 55140 226222 55260 226250
rect 56232 226238 56284 226244
rect 53840 225752 53892 225758
rect 53840 225694 53892 225700
rect 53852 222902 53880 225694
rect 55232 222970 55260 226222
rect 55220 222964 55272 222970
rect 55220 222906 55272 222912
rect 53840 222896 53892 222902
rect 53840 222838 53892 222844
rect 56244 222154 56272 226238
rect 55128 222148 55180 222154
rect 55128 222090 55180 222096
rect 56232 222148 56284 222154
rect 56232 222090 56284 222096
rect 55140 217682 55168 222090
rect 55140 217654 55260 217682
rect 50436 215144 50488 215150
rect 50436 215086 50488 215092
rect 54484 215144 54536 215150
rect 54484 215086 54536 215092
rect 50344 213920 50396 213926
rect 50344 213862 50396 213868
rect 53104 213920 53156 213926
rect 53104 213862 53156 213868
rect 53116 209506 53144 213862
rect 53104 209500 53156 209506
rect 53104 209442 53156 209448
rect 45560 201476 45612 201482
rect 45560 201418 45612 201424
rect 47584 201476 47636 201482
rect 47584 201418 47636 201424
rect 46204 181484 46256 181490
rect 46204 181426 46256 181432
rect 46216 137290 46244 181426
rect 47596 171834 47624 201418
rect 54496 186998 54524 215086
rect 55232 214130 55260 217654
rect 55220 214124 55272 214130
rect 55220 214066 55272 214072
rect 54576 209500 54628 209506
rect 54576 209442 54628 209448
rect 54588 197334 54616 209442
rect 54576 197328 54628 197334
rect 54576 197270 54628 197276
rect 56508 197328 56560 197334
rect 56508 197270 56560 197276
rect 56520 190454 56548 197270
rect 56612 195974 56640 230588
rect 57336 222964 57388 222970
rect 57336 222906 57388 222912
rect 57244 222148 57296 222154
rect 57244 222090 57296 222096
rect 57256 211138 57284 222090
rect 57348 217326 57376 222906
rect 57336 217320 57388 217326
rect 57336 217262 57388 217268
rect 62776 215966 62804 232358
rect 64880 231056 64932 231062
rect 64880 230998 64932 231004
rect 64892 226370 64920 230998
rect 64880 226364 64932 226370
rect 64880 226306 64932 226312
rect 69572 226364 69624 226370
rect 69572 226306 69624 226312
rect 69584 219434 69612 226306
rect 69664 222896 69716 222902
rect 69664 222838 69716 222844
rect 69676 220114 69704 222838
rect 69664 220108 69716 220114
rect 69664 220050 69716 220056
rect 79324 220108 79376 220114
rect 79324 220050 79376 220056
rect 69584 219406 69704 219434
rect 69676 218686 69704 219406
rect 69664 218680 69716 218686
rect 69664 218622 69716 218628
rect 71872 218680 71924 218686
rect 71872 218622 71924 218628
rect 67548 217320 67600 217326
rect 67548 217262 67600 217268
rect 62764 215960 62816 215966
rect 62764 215902 62816 215908
rect 67560 215626 67588 217262
rect 70400 215960 70452 215966
rect 70400 215902 70452 215908
rect 67548 215620 67600 215626
rect 67548 215562 67600 215568
rect 69020 215620 69072 215626
rect 69020 215562 69072 215568
rect 57336 214124 57388 214130
rect 57336 214066 57388 214072
rect 57244 211132 57296 211138
rect 57244 211074 57296 211080
rect 57348 208418 57376 214066
rect 69032 213586 69060 215562
rect 69020 213580 69072 213586
rect 69020 213522 69072 213528
rect 70412 213042 70440 215902
rect 71884 214606 71912 218622
rect 71872 214600 71924 214606
rect 71872 214542 71924 214548
rect 73988 214600 74040 214606
rect 73988 214542 74040 214548
rect 71044 213580 71096 213586
rect 71044 213522 71096 213528
rect 70400 213036 70452 213042
rect 70400 212978 70452 212984
rect 58624 211132 58676 211138
rect 58624 211074 58676 211080
rect 57336 208412 57388 208418
rect 57336 208354 57388 208360
rect 58636 202842 58664 211074
rect 71056 208962 71084 213522
rect 73804 213036 73856 213042
rect 73804 212978 73856 212984
rect 71044 208956 71096 208962
rect 71044 208898 71096 208904
rect 63500 208344 63552 208350
rect 63500 208286 63552 208292
rect 63512 204270 63540 208286
rect 63500 204264 63552 204270
rect 63500 204206 63552 204212
rect 65524 204264 65576 204270
rect 65524 204206 65576 204212
rect 58624 202836 58676 202842
rect 58624 202778 58676 202784
rect 63500 202836 63552 202842
rect 63500 202778 63552 202784
rect 63512 198014 63540 202778
rect 63500 198008 63552 198014
rect 63500 197950 63552 197956
rect 56600 195968 56652 195974
rect 56600 195910 56652 195916
rect 56520 190426 56640 190454
rect 54484 186992 54536 186998
rect 54484 186934 54536 186940
rect 56612 186454 56640 190426
rect 56600 186448 56652 186454
rect 56600 186390 56652 186396
rect 58624 186448 58676 186454
rect 58624 186390 58676 186396
rect 58636 175234 58664 186390
rect 58624 175228 58676 175234
rect 58624 175170 58676 175176
rect 60648 175228 60700 175234
rect 60648 175170 60700 175176
rect 60660 172582 60688 175170
rect 60648 172576 60700 172582
rect 60648 172518 60700 172524
rect 65536 172514 65564 204206
rect 73816 199442 73844 212978
rect 74000 209778 74028 214542
rect 73988 209772 74040 209778
rect 73988 209714 74040 209720
rect 75460 209772 75512 209778
rect 75460 209714 75512 209720
rect 73896 208956 73948 208962
rect 73896 208898 73948 208904
rect 73804 199436 73856 199442
rect 73804 199378 73856 199384
rect 69572 198008 69624 198014
rect 69572 197950 69624 197956
rect 69584 196178 69612 197950
rect 73908 197334 73936 208898
rect 75472 208350 75500 209714
rect 79336 209098 79364 220050
rect 80716 214606 80744 232358
rect 393964 231872 394016 231878
rect 393964 231814 394016 231820
rect 142160 231192 142212 231198
rect 142160 231134 142212 231140
rect 80704 214600 80756 214606
rect 80704 214542 80756 214548
rect 79324 209092 79376 209098
rect 79324 209034 79376 209040
rect 75460 208344 75512 208350
rect 75460 208286 75512 208292
rect 77576 208344 77628 208350
rect 77576 208286 77628 208292
rect 77588 204882 77616 208286
rect 77576 204876 77628 204882
rect 77576 204818 77628 204824
rect 80060 204876 80112 204882
rect 80060 204818 80112 204824
rect 80072 202842 80100 204818
rect 80060 202836 80112 202842
rect 80060 202778 80112 202784
rect 81808 202836 81860 202842
rect 81808 202778 81860 202784
rect 81820 199442 81848 202778
rect 81440 199436 81492 199442
rect 81440 199378 81492 199384
rect 81808 199436 81860 199442
rect 81808 199378 81860 199384
rect 73896 197328 73948 197334
rect 73896 197270 73948 197276
rect 76288 197328 76340 197334
rect 76288 197270 76340 197276
rect 69572 196172 69624 196178
rect 69572 196114 69624 196120
rect 71780 196172 71832 196178
rect 71780 196114 71832 196120
rect 71792 193186 71820 196114
rect 76300 195906 76328 197270
rect 81452 196654 81480 199378
rect 81440 196648 81492 196654
rect 81440 196590 81492 196596
rect 86972 195906 87000 230588
rect 115952 230574 116518 230602
rect 91744 214600 91796 214606
rect 91744 214542 91796 214548
rect 91100 209092 91152 209098
rect 91100 209034 91152 209040
rect 91112 206310 91140 209034
rect 91756 208350 91784 214542
rect 91744 208344 91796 208350
rect 91744 208286 91796 208292
rect 95148 208344 95200 208350
rect 95148 208286 95200 208292
rect 91100 206304 91152 206310
rect 91100 206246 91152 206252
rect 95160 204950 95188 208286
rect 104716 206304 104768 206310
rect 104716 206246 104768 206252
rect 95148 204944 95200 204950
rect 95148 204886 95200 204892
rect 104728 202842 104756 206246
rect 106648 204944 106700 204950
rect 106648 204886 106700 204892
rect 104716 202836 104768 202842
rect 104716 202778 104768 202784
rect 106660 202774 106688 204886
rect 108672 202836 108724 202842
rect 108672 202778 108724 202784
rect 106648 202768 106700 202774
rect 106648 202710 106700 202716
rect 88984 199436 89036 199442
rect 88984 199378 89036 199384
rect 88340 196648 88392 196654
rect 88340 196590 88392 196596
rect 76288 195900 76340 195906
rect 76288 195842 76340 195848
rect 77944 195900 77996 195906
rect 77944 195842 77996 195848
rect 86960 195900 87012 195906
rect 86960 195842 87012 195848
rect 71780 193180 71832 193186
rect 71780 193122 71832 193128
rect 74264 193180 74316 193186
rect 74264 193122 74316 193128
rect 68284 186992 68336 186998
rect 68284 186934 68336 186940
rect 68296 176662 68324 186934
rect 74276 186318 74304 193122
rect 74264 186312 74316 186318
rect 74264 186254 74316 186260
rect 76564 186312 76616 186318
rect 76564 186254 76616 186260
rect 68284 176656 68336 176662
rect 68284 176598 68336 176604
rect 76576 172514 76604 186254
rect 76656 176656 76708 176662
rect 76656 176598 76708 176604
rect 63500 172508 63552 172514
rect 63500 172450 63552 172456
rect 65524 172508 65576 172514
rect 65524 172450 65576 172456
rect 66260 172508 66312 172514
rect 66260 172450 66312 172456
rect 76564 172508 76616 172514
rect 76564 172450 76616 172456
rect 47584 171828 47636 171834
rect 47584 171770 47636 171776
rect 61660 171828 61712 171834
rect 61660 171770 61712 171776
rect 61672 168774 61700 171770
rect 63512 169590 63540 172450
rect 66272 169590 66300 172450
rect 63500 169584 63552 169590
rect 63500 169526 63552 169532
rect 65616 169584 65668 169590
rect 65616 169526 65668 169532
rect 66260 169584 66312 169590
rect 66260 169526 66312 169532
rect 69664 169584 69716 169590
rect 69664 169526 69716 169532
rect 61660 168768 61712 168774
rect 61660 168710 61712 168716
rect 63500 168768 63552 168774
rect 63500 168710 63552 168716
rect 63512 166326 63540 168710
rect 63500 166320 63552 166326
rect 63500 166262 63552 166268
rect 65628 162858 65656 169526
rect 65616 162852 65668 162858
rect 65616 162794 65668 162800
rect 69676 144906 69704 169526
rect 75184 166320 75236 166326
rect 75184 166262 75236 166268
rect 71044 162852 71096 162858
rect 71044 162794 71096 162800
rect 71056 153882 71084 162794
rect 75196 158030 75224 166262
rect 76668 164218 76696 176598
rect 77956 175234 77984 195842
rect 88352 193594 88380 196590
rect 88340 193588 88392 193594
rect 88340 193530 88392 193536
rect 88996 190670 89024 199378
rect 108684 197538 108712 202778
rect 110236 202768 110288 202774
rect 110236 202710 110288 202716
rect 110248 198014 110276 202710
rect 110236 198008 110288 198014
rect 110236 197950 110288 197956
rect 108672 197532 108724 197538
rect 108672 197474 108724 197480
rect 111064 197532 111116 197538
rect 111064 197474 111116 197480
rect 91744 193588 91796 193594
rect 91744 193530 91796 193536
rect 88984 190664 89036 190670
rect 88984 190606 89036 190612
rect 77944 175228 77996 175234
rect 77944 175170 77996 175176
rect 79416 175228 79468 175234
rect 79416 175170 79468 175176
rect 79324 172508 79376 172514
rect 79324 172450 79376 172456
rect 76656 164212 76708 164218
rect 76656 164154 76708 164160
rect 75184 158024 75236 158030
rect 75184 157966 75236 157972
rect 71044 153876 71096 153882
rect 71044 153818 71096 153824
rect 69664 144900 69716 144906
rect 69664 144842 69716 144848
rect 71044 144900 71096 144906
rect 71044 144842 71096 144848
rect 46204 137284 46256 137290
rect 46204 137226 46256 137232
rect 71056 132054 71084 144842
rect 71044 132048 71096 132054
rect 71044 131990 71096 131996
rect 72516 132048 72568 132054
rect 72516 131990 72568 131996
rect 72528 125594 72556 131990
rect 72516 125588 72568 125594
rect 72516 125530 72568 125536
rect 73896 125588 73948 125594
rect 73896 125530 73948 125536
rect 73908 122738 73936 125530
rect 73896 122732 73948 122738
rect 73896 122674 73948 122680
rect 75460 122732 75512 122738
rect 75460 122674 75512 122680
rect 43444 118652 43496 118658
rect 43444 118594 43496 118600
rect 75472 114578 75500 122674
rect 79336 118318 79364 172450
rect 79428 143546 79456 175170
rect 91756 171222 91784 193530
rect 93860 190664 93912 190670
rect 93860 190606 93912 190612
rect 93872 187950 93900 190606
rect 93860 187944 93912 187950
rect 93860 187886 93912 187892
rect 95884 187944 95936 187950
rect 95884 187886 95936 187892
rect 95896 175302 95924 187886
rect 111076 186318 111104 197474
rect 115952 194614 115980 230574
rect 142172 228342 142200 231134
rect 180800 231124 180852 231130
rect 180800 231066 180852 231072
rect 385684 231124 385736 231130
rect 385684 231066 385736 231072
rect 146312 230574 146510 230602
rect 142160 228336 142212 228342
rect 142160 228278 142212 228284
rect 143540 228336 143592 228342
rect 143540 228278 143592 228284
rect 143552 220114 143580 228278
rect 143540 220108 143592 220114
rect 143540 220050 143592 220056
rect 119436 218068 119488 218074
rect 119436 218010 119488 218016
rect 117320 198008 117372 198014
rect 117320 197950 117372 197956
rect 115940 194608 115992 194614
rect 115940 194550 115992 194556
rect 117332 194410 117360 197950
rect 117320 194404 117372 194410
rect 117320 194346 117372 194352
rect 116584 187740 116636 187746
rect 116584 187682 116636 187688
rect 111064 186312 111116 186318
rect 111064 186254 111116 186260
rect 113824 186312 113876 186318
rect 113824 186254 113876 186260
rect 113836 178974 113864 186254
rect 113824 178968 113876 178974
rect 113824 178910 113876 178916
rect 95884 175296 95936 175302
rect 95884 175238 95936 175244
rect 100024 175228 100076 175234
rect 100024 175170 100076 175176
rect 91744 171216 91796 171222
rect 91744 171158 91796 171164
rect 94504 171216 94556 171222
rect 94504 171158 94556 171164
rect 94516 164218 94544 171158
rect 100036 165646 100064 175170
rect 100024 165640 100076 165646
rect 100024 165582 100076 165588
rect 102784 165572 102836 165578
rect 102784 165514 102836 165520
rect 81808 164212 81860 164218
rect 81808 164154 81860 164160
rect 94504 164212 94556 164218
rect 94504 164154 94556 164160
rect 97264 164212 97316 164218
rect 97264 164154 97316 164160
rect 81820 161294 81848 164154
rect 81808 161288 81860 161294
rect 81808 161230 81860 161236
rect 85488 161288 85540 161294
rect 85488 161230 85540 161236
rect 85500 155922 85528 161230
rect 86132 158024 86184 158030
rect 86132 157966 86184 157972
rect 85488 155916 85540 155922
rect 85488 155858 85540 155864
rect 86144 154562 86172 157966
rect 90364 155916 90416 155922
rect 90364 155858 90416 155864
rect 86132 154556 86184 154562
rect 86132 154498 86184 154504
rect 79416 143540 79468 143546
rect 79416 143482 79468 143488
rect 80704 143540 80756 143546
rect 80704 143482 80756 143488
rect 80716 120698 80744 143482
rect 90376 140622 90404 155858
rect 91744 154556 91796 154562
rect 91744 154498 91796 154504
rect 90364 140616 90416 140622
rect 90364 140558 90416 140564
rect 91756 134638 91784 154498
rect 97276 152318 97304 164154
rect 100024 153876 100076 153882
rect 100024 153818 100076 153824
rect 97264 152312 97316 152318
rect 97264 152254 97316 152260
rect 94504 140616 94556 140622
rect 94504 140558 94556 140564
rect 94516 136542 94544 140558
rect 100036 138922 100064 153818
rect 102796 151434 102824 165514
rect 103612 152312 103664 152318
rect 103612 152254 103664 152260
rect 102784 151428 102836 151434
rect 102784 151370 102836 151376
rect 103624 149598 103652 152254
rect 104532 151428 104584 151434
rect 104532 151370 104584 151376
rect 103612 149592 103664 149598
rect 103612 149534 103664 149540
rect 104544 148918 104572 151370
rect 109684 149592 109736 149598
rect 109684 149534 109736 149540
rect 104532 148912 104584 148918
rect 104532 148854 104584 148860
rect 106280 148912 106332 148918
rect 106280 148854 106332 148860
rect 106292 142186 106320 148854
rect 106280 142180 106332 142186
rect 106280 142122 106332 142128
rect 100024 138916 100076 138922
rect 100024 138858 100076 138864
rect 94504 136536 94556 136542
rect 94504 136478 94556 136484
rect 100116 136536 100168 136542
rect 100116 136478 100168 136484
rect 91744 134632 91796 134638
rect 91744 134574 91796 134580
rect 94228 134632 94280 134638
rect 94228 134574 94280 134580
rect 94240 131238 94268 134574
rect 100128 131986 100156 136478
rect 100116 131980 100168 131986
rect 100116 131922 100168 131928
rect 105544 131980 105596 131986
rect 105544 131922 105596 131928
rect 94228 131232 94280 131238
rect 94228 131174 94280 131180
rect 99380 131232 99432 131238
rect 99380 131174 99432 131180
rect 99392 126886 99420 131174
rect 99380 126880 99432 126886
rect 99380 126822 99432 126828
rect 80704 120692 80756 120698
rect 80704 120634 80756 120640
rect 82820 120692 82872 120698
rect 82820 120634 82872 120640
rect 82832 118590 82860 120634
rect 105556 119134 105584 131922
rect 106188 126880 106240 126886
rect 106188 126822 106240 126828
rect 106200 123486 106228 126822
rect 106188 123480 106240 123486
rect 106188 123422 106240 123428
rect 105544 119128 105596 119134
rect 105544 119070 105596 119076
rect 82820 118584 82872 118590
rect 82820 118526 82872 118532
rect 86224 118584 86276 118590
rect 86224 118526 86276 118532
rect 79324 118312 79376 118318
rect 79324 118254 79376 118260
rect 81072 118312 81124 118318
rect 81072 118254 81124 118260
rect 81084 115870 81112 118254
rect 81072 115864 81124 115870
rect 81072 115806 81124 115812
rect 82728 115864 82780 115870
rect 82728 115806 82780 115812
rect 75460 114572 75512 114578
rect 75460 114514 75512 114520
rect 81348 114504 81400 114510
rect 81348 114446 81400 114452
rect 33784 113144 33836 113150
rect 33784 113086 33836 113092
rect 19984 111784 20036 111790
rect 19984 111726 20036 111732
rect 81360 110498 81388 114446
rect 81348 110492 81400 110498
rect 81348 110434 81400 110440
rect 82740 110378 82768 115806
rect 86236 112470 86264 118526
rect 86224 112464 86276 112470
rect 86224 112406 86276 112412
rect 87420 112464 87472 112470
rect 87420 112406 87472 112412
rect 82740 110350 82860 110378
rect 82832 107642 82860 110350
rect 87432 109750 87460 112406
rect 87420 109744 87472 109750
rect 87420 109686 87472 109692
rect 97908 109744 97960 109750
rect 97908 109686 97960 109692
rect 97920 109002 97948 109686
rect 97908 108996 97960 109002
rect 97908 108938 97960 108944
rect 82820 107636 82872 107642
rect 82820 107578 82872 107584
rect 109696 107574 109724 149534
rect 109776 142112 109828 142118
rect 109776 142054 109828 142060
rect 109788 121990 109816 142054
rect 115296 123480 115348 123486
rect 115296 123422 115348 123428
rect 109776 121984 109828 121990
rect 109776 121926 109828 121932
rect 111800 121984 111852 121990
rect 111800 121926 111852 121932
rect 109776 119128 109828 119134
rect 109776 119070 109828 119076
rect 109684 107568 109736 107574
rect 109684 107510 109736 107516
rect 109788 102066 109816 119070
rect 111812 117230 111840 121926
rect 111800 117224 111852 117230
rect 111800 117166 111852 117172
rect 115204 117224 115256 117230
rect 115204 117166 115256 117172
rect 112444 107568 112496 107574
rect 112444 107510 112496 107516
rect 109776 102060 109828 102066
rect 109776 102002 109828 102008
rect 6918 78160 6974 78169
rect 6918 78095 6974 78104
rect 112456 77994 112484 107510
rect 115216 97986 115244 117166
rect 115308 111790 115336 123422
rect 115296 111784 115348 111790
rect 115296 111726 115348 111732
rect 115848 102060 115900 102066
rect 115848 102002 115900 102008
rect 115204 97980 115256 97986
rect 115204 97922 115256 97928
rect 115860 95198 115888 102002
rect 115848 95192 115900 95198
rect 115848 95134 115900 95140
rect 112444 77988 112496 77994
rect 112444 77930 112496 77936
rect 116596 77178 116624 187682
rect 117964 178968 118016 178974
rect 117964 178910 118016 178916
rect 117872 138032 117924 138038
rect 117872 137974 117924 137980
rect 117320 137284 117372 137290
rect 117320 137226 117372 137232
rect 117332 137193 117360 137226
rect 117318 137184 117374 137193
rect 117318 137119 117374 137128
rect 116676 136740 116728 136746
rect 116676 136682 116728 136688
rect 116584 77172 116636 77178
rect 116584 77114 116636 77120
rect 116688 77110 116716 136682
rect 117318 134056 117374 134065
rect 117318 133991 117374 134000
rect 117332 133958 117360 133991
rect 117320 133952 117372 133958
rect 117320 133894 117372 133900
rect 117318 132560 117374 132569
rect 117318 132495 117320 132504
rect 117372 132495 117374 132504
rect 117320 132466 117372 132472
rect 117318 131200 117374 131209
rect 117318 131135 117320 131144
rect 117372 131135 117374 131144
rect 117320 131106 117372 131112
rect 117320 129736 117372 129742
rect 117318 129704 117320 129713
rect 117372 129704 117374 129713
rect 117318 129639 117374 129648
rect 117320 128308 117372 128314
rect 117320 128250 117372 128256
rect 117332 128217 117360 128250
rect 117318 128208 117374 128217
rect 117318 128143 117374 128152
rect 117320 126948 117372 126954
rect 117320 126890 117372 126896
rect 117332 126857 117360 126890
rect 117318 126848 117374 126857
rect 117318 126783 117374 126792
rect 117320 124160 117372 124166
rect 117320 124102 117372 124108
rect 117332 123865 117360 124102
rect 117318 123856 117374 123865
rect 117318 123791 117374 123800
rect 117320 122800 117372 122806
rect 117318 122768 117320 122777
rect 117372 122768 117374 122777
rect 117318 122703 117374 122712
rect 117320 121440 117372 121446
rect 117320 121382 117372 121388
rect 117332 121281 117360 121382
rect 117318 121272 117374 121281
rect 117318 121207 117374 121216
rect 117320 120080 117372 120086
rect 117320 120022 117372 120028
rect 117332 119785 117360 120022
rect 117318 119776 117374 119785
rect 117318 119711 117374 119720
rect 117320 118652 117372 118658
rect 117320 118594 117372 118600
rect 117332 118289 117360 118594
rect 117318 118280 117374 118289
rect 117318 118215 117374 118224
rect 117320 117292 117372 117298
rect 117320 117234 117372 117240
rect 117332 116793 117360 117234
rect 117318 116784 117374 116793
rect 117318 116719 117374 116728
rect 117320 115932 117372 115938
rect 117320 115874 117372 115880
rect 117332 115297 117360 115874
rect 117318 115288 117374 115297
rect 117318 115223 117374 115232
rect 117320 113144 117372 113150
rect 117318 113112 117320 113121
rect 117372 113112 117374 113121
rect 117318 113047 117374 113056
rect 117320 111784 117372 111790
rect 117318 111752 117320 111761
rect 117372 111752 117374 111761
rect 117318 111687 117374 111696
rect 117320 110424 117372 110430
rect 117320 110366 117372 110372
rect 117332 110265 117360 110366
rect 117318 110256 117374 110265
rect 117318 110191 117374 110200
rect 117320 108996 117372 109002
rect 117320 108938 117372 108944
rect 117332 108905 117360 108938
rect 117318 108896 117374 108905
rect 117318 108831 117374 108840
rect 117320 107636 117372 107642
rect 117320 107578 117372 107584
rect 117332 107545 117360 107578
rect 117318 107536 117374 107545
rect 117318 107471 117374 107480
rect 116768 97980 116820 97986
rect 116768 97922 116820 97928
rect 116780 89010 116808 97922
rect 116768 89004 116820 89010
rect 116768 88946 116820 88952
rect 117884 83745 117912 137974
rect 117976 98734 118004 178910
rect 118700 171828 118752 171834
rect 118700 171770 118752 171776
rect 118332 142860 118384 142866
rect 118332 142802 118384 142808
rect 118146 137184 118202 137193
rect 118146 137119 118202 137128
rect 118160 125497 118188 137119
rect 118238 135552 118294 135561
rect 118238 135487 118294 135496
rect 118146 125488 118202 125497
rect 118146 125423 118202 125432
rect 118148 114844 118200 114850
rect 118148 114786 118200 114792
rect 117964 98728 118016 98734
rect 117964 98670 118016 98676
rect 117964 89004 118016 89010
rect 117964 88946 118016 88952
rect 117870 83736 117926 83745
rect 117870 83671 117926 83680
rect 117976 81462 118004 88946
rect 118160 86873 118188 114786
rect 118252 95169 118280 135487
rect 118238 95160 118294 95169
rect 118238 95095 118294 95104
rect 118344 91089 118372 142802
rect 118516 141568 118568 141574
rect 118516 141510 118568 141516
rect 118424 141500 118476 141506
rect 118424 141442 118476 141448
rect 118330 91080 118386 91089
rect 118330 91015 118386 91024
rect 118436 89729 118464 141442
rect 118422 89720 118478 89729
rect 118422 89655 118478 89664
rect 118528 88233 118556 141510
rect 118608 124160 118660 124166
rect 118608 124102 118660 124108
rect 118620 106185 118648 124102
rect 118606 106176 118662 106185
rect 118606 106111 118662 106120
rect 118712 92449 118740 171770
rect 118792 146940 118844 146946
rect 118792 146882 118844 146888
rect 118698 92440 118754 92449
rect 118698 92375 118754 92384
rect 118514 88224 118570 88233
rect 118514 88159 118570 88168
rect 118146 86864 118202 86873
rect 118146 86799 118202 86808
rect 118804 85377 118832 146882
rect 119068 145580 119120 145586
rect 119068 145522 119120 145528
rect 118976 144220 119028 144226
rect 118976 144162 119028 144168
rect 118884 140072 118936 140078
rect 118884 140014 118936 140020
rect 118896 93809 118924 140014
rect 118988 100337 119016 144162
rect 119080 103193 119108 145522
rect 119160 141432 119212 141438
rect 119160 141374 119212 141380
rect 119066 103184 119122 103193
rect 119066 103119 119122 103128
rect 118974 100328 119030 100337
rect 118974 100263 119030 100272
rect 119172 98841 119200 141374
rect 119344 140208 119396 140214
rect 119344 140150 119396 140156
rect 119252 138712 119304 138718
rect 119252 138654 119304 138660
rect 119158 98832 119214 98841
rect 119158 98767 119214 98776
rect 119264 97345 119292 138654
rect 119356 104825 119384 140150
rect 119448 114850 119476 218010
rect 146312 197418 146340 230574
rect 176672 229770 176700 230588
rect 166264 229764 166316 229770
rect 166264 229706 166316 229712
rect 176660 229764 176712 229770
rect 176660 229706 176712 229712
rect 157984 228472 158036 228478
rect 157984 228414 158036 228420
rect 155960 199436 156012 199442
rect 155960 199378 156012 199384
rect 148968 198008 149020 198014
rect 148968 197950 149020 197956
rect 146142 197390 146340 197418
rect 148980 197404 149008 197950
rect 155972 197470 156000 199378
rect 154488 197464 154540 197470
rect 154146 197412 154488 197418
rect 154146 197406 154540 197412
rect 155960 197464 156012 197470
rect 155960 197406 156012 197412
rect 154146 197390 154528 197406
rect 157996 197334 158024 228414
rect 158628 220108 158680 220114
rect 158628 220050 158680 220056
rect 158640 219434 158668 220050
rect 158640 219406 158760 219434
rect 158732 213926 158760 219406
rect 158720 213920 158772 213926
rect 158720 213862 158772 213868
rect 160100 213920 160152 213926
rect 160100 213862 160152 213868
rect 160112 211206 160140 213862
rect 160100 211200 160152 211206
rect 160100 211142 160152 211148
rect 162860 211132 162912 211138
rect 162860 211074 162912 211080
rect 162872 209166 162900 211074
rect 162860 209160 162912 209166
rect 162860 209102 162912 209108
rect 164240 209160 164292 209166
rect 164240 209102 164292 209108
rect 164252 206718 164280 209102
rect 164240 206712 164292 206718
rect 164240 206654 164292 206660
rect 152740 197328 152792 197334
rect 152582 197276 152740 197282
rect 152582 197270 152792 197276
rect 157984 197328 158036 197334
rect 157984 197270 158036 197276
rect 152582 197254 152780 197270
rect 166276 196790 166304 229706
rect 166356 206712 166408 206718
rect 166356 206654 166408 206660
rect 147956 196784 148008 196790
rect 147798 196732 147956 196738
rect 147798 196726 148008 196732
rect 166264 196784 166316 196790
rect 166264 196726 166316 196732
rect 147798 196710 147996 196726
rect 160836 196716 160888 196722
rect 160836 196658 160888 196664
rect 151176 196648 151228 196654
rect 150926 196596 151176 196602
rect 150926 196590 151228 196596
rect 150926 196574 151216 196590
rect 140424 196030 140530 196058
rect 157366 196030 157564 196058
rect 138112 195968 138164 195974
rect 138110 195936 138112 195945
rect 140424 195945 140452 196030
rect 157536 195974 157564 196030
rect 157524 195968 157576 195974
rect 138164 195936 138166 195945
rect 140410 195936 140466 195945
rect 138110 195871 138166 195880
rect 139400 195900 139452 195906
rect 158916 195937 158944 196044
rect 160848 195945 160876 196658
rect 157524 195910 157576 195916
rect 158902 195928 158958 195937
rect 140410 195871 140466 195880
rect 157432 195900 157484 195906
rect 139400 195842 139452 195848
rect 158902 195863 158958 195872
rect 160834 195936 160890 195945
rect 160834 195871 160890 195880
rect 157432 195842 157484 195848
rect 139412 195537 139440 195842
rect 140778 195664 140834 195673
rect 140778 195599 140834 195608
rect 157154 195664 157210 195673
rect 157444 195650 157472 195842
rect 157210 195622 157472 195650
rect 157154 195599 157210 195608
rect 139398 195528 139454 195537
rect 139398 195463 139454 195472
rect 140792 194614 140820 195599
rect 140780 194608 140832 194614
rect 140780 194550 140832 194556
rect 120724 194404 120776 194410
rect 120724 194346 120776 194352
rect 120736 189310 120764 194346
rect 166368 193186 166396 206654
rect 166356 193180 166408 193186
rect 166356 193122 166408 193128
rect 168472 193180 168524 193186
rect 168472 193122 168524 193128
rect 140962 191856 141018 191865
rect 140962 191791 141018 191800
rect 140870 191720 140926 191729
rect 140870 191655 140926 191664
rect 140778 191584 140834 191593
rect 140778 191519 140834 191528
rect 140792 190618 140820 191519
rect 140700 190590 140820 190618
rect 140700 190454 140728 190590
rect 140780 190528 140832 190534
rect 140780 190470 140832 190476
rect 140608 190426 140728 190454
rect 140608 190074 140636 190426
rect 140792 190398 140820 190470
rect 140780 190392 140832 190398
rect 140884 190369 140912 191655
rect 140976 191010 141004 191791
rect 144550 191040 144606 191049
rect 140964 191004 141016 191010
rect 144302 190998 144550 191026
rect 144550 190975 144606 190984
rect 140964 190946 141016 190952
rect 140962 190904 141018 190913
rect 140962 190839 141018 190848
rect 140780 190334 140832 190340
rect 140870 190360 140926 190369
rect 140870 190295 140926 190304
rect 140872 190256 140924 190262
rect 140872 190198 140924 190204
rect 140608 190046 140820 190074
rect 120724 189304 120776 189310
rect 120724 189246 120776 189252
rect 123668 189304 123720 189310
rect 123668 189246 123720 189252
rect 123680 182170 123708 189246
rect 140792 184249 140820 190046
rect 140778 184240 140834 184249
rect 140778 184175 140834 184184
rect 140884 184113 140912 190198
rect 140976 184385 141004 190839
rect 144460 190528 144512 190534
rect 144380 190476 144460 190482
rect 144380 190470 144512 190476
rect 144380 190454 144500 190470
rect 140962 184376 141018 184385
rect 140962 184311 141018 184320
rect 140870 184104 140926 184113
rect 140870 184039 140926 184048
rect 123668 182164 123720 182170
rect 123668 182106 123720 182112
rect 126520 182164 126572 182170
rect 126520 182106 126572 182112
rect 136376 182158 136758 182186
rect 121460 180124 121512 180130
rect 121460 180066 121512 180072
rect 120724 140140 120776 140146
rect 120724 140082 120776 140088
rect 120632 138984 120684 138990
rect 120632 138926 120684 138932
rect 119528 137284 119580 137290
rect 119528 137226 119580 137232
rect 119540 124166 119568 137226
rect 120644 136241 120672 138926
rect 120630 136232 120686 136241
rect 120630 136167 120686 136176
rect 119528 124160 119580 124166
rect 119528 124102 119580 124108
rect 119436 114844 119488 114850
rect 119436 114786 119488 114792
rect 119342 104816 119398 104825
rect 119342 104751 119398 104760
rect 120736 103514 120764 140082
rect 121472 137986 121500 180066
rect 124864 178764 124916 178770
rect 124864 178706 124916 178712
rect 124220 177336 124272 177342
rect 124220 177278 124272 177284
rect 124232 151814 124260 177278
rect 124232 151786 124536 151814
rect 123668 139800 123720 139806
rect 123668 139742 123720 139748
rect 123680 137986 123708 139742
rect 121472 137958 121808 137986
rect 123372 137958 123708 137986
rect 124508 137986 124536 151786
rect 124876 139806 124904 178706
rect 126532 178702 126560 182106
rect 136376 180130 136404 182158
rect 144380 182036 144408 190454
rect 145012 190324 145064 190330
rect 145012 190266 145064 190272
rect 145024 188970 145052 190266
rect 145852 189774 145958 189802
rect 145852 189009 145880 189774
rect 166106 189366 166212 189394
rect 145838 189000 145894 189009
rect 144644 188964 144696 188970
rect 144644 188906 144696 188912
rect 145012 188964 145064 188970
rect 145838 188935 145894 188944
rect 145012 188906 145064 188912
rect 144656 181558 144684 188906
rect 144918 182200 144974 182209
rect 144918 182135 144974 182144
rect 144644 181552 144696 181558
rect 144644 181494 144696 181500
rect 144932 181257 144960 182135
rect 145196 181552 145248 181558
rect 145196 181494 145248 181500
rect 145208 181257 145236 181494
rect 144918 181248 144974 181257
rect 144918 181183 144974 181192
rect 145194 181248 145250 181257
rect 145194 181183 145250 181192
rect 144642 180976 144698 180985
rect 136468 180934 136758 180962
rect 144578 180934 144642 180962
rect 136364 180124 136416 180130
rect 136364 180066 136416 180072
rect 136364 178832 136416 178838
rect 136364 178774 136416 178780
rect 126520 178696 126572 178702
rect 126520 178638 126572 178644
rect 135996 177812 136048 177818
rect 135996 177754 136048 177760
rect 136008 176118 136036 177754
rect 126980 176112 127032 176118
rect 126980 176054 127032 176060
rect 135996 176112 136048 176118
rect 135996 176054 136048 176060
rect 125600 175976 125652 175982
rect 125600 175918 125652 175924
rect 125612 151814 125640 175918
rect 126992 151814 127020 176054
rect 136376 176050 136404 178774
rect 136468 178770 136496 180934
rect 144642 180911 144698 180920
rect 136560 179982 136758 180010
rect 136456 178764 136508 178770
rect 136456 178706 136508 178712
rect 136560 177970 136588 179982
rect 165172 179382 165200 188020
rect 166184 187678 166212 189366
rect 166172 187672 166224 187678
rect 166172 187614 166224 187620
rect 168484 184890 168512 193122
rect 180064 191888 180116 191894
rect 180064 191830 180116 191836
rect 168472 184884 168524 184890
rect 168472 184826 168524 184832
rect 170404 184884 170456 184890
rect 170404 184826 170456 184832
rect 158812 179376 158864 179382
rect 158812 179318 158864 179324
rect 165160 179376 165212 179382
rect 165160 179318 165212 179324
rect 136744 178838 136772 179044
rect 144090 178936 144146 178945
rect 144090 178871 144146 178880
rect 136732 178832 136784 178838
rect 136732 178774 136784 178780
rect 141606 178800 141662 178809
rect 141606 178735 141662 178744
rect 141790 178800 141846 178809
rect 141790 178735 141846 178744
rect 136468 177942 136588 177970
rect 136468 177342 136496 177942
rect 136744 177834 136772 177956
rect 136652 177818 136772 177834
rect 136640 177812 136772 177818
rect 136692 177806 136772 177812
rect 136640 177754 136692 177760
rect 136456 177336 136508 177342
rect 136456 177278 136508 177284
rect 136468 176990 136758 177018
rect 136364 176044 136416 176050
rect 136364 175986 136416 175992
rect 136468 175234 136496 176990
rect 136560 175902 136758 175930
rect 128360 175228 128412 175234
rect 128360 175170 128412 175176
rect 136456 175228 136508 175234
rect 136456 175170 136508 175176
rect 128372 151814 128400 175170
rect 133880 173936 133932 173942
rect 133880 173878 133932 173884
rect 136560 173894 136588 175902
rect 141620 175710 141648 178735
rect 141804 176118 141832 178735
rect 142066 178664 142122 178673
rect 142066 178599 142122 178608
rect 141792 176112 141844 176118
rect 141792 176054 141844 176060
rect 141608 175704 141660 175710
rect 141608 175646 141660 175652
rect 131120 172576 131172 172582
rect 131120 172518 131172 172524
rect 125612 151786 126100 151814
rect 126992 151786 127664 151814
rect 128372 151786 129228 151814
rect 124864 139800 124916 139806
rect 124864 139742 124916 139748
rect 126072 137986 126100 151786
rect 127636 137986 127664 151786
rect 129200 137986 129228 151786
rect 131132 137986 131160 172518
rect 132500 171148 132552 171154
rect 132500 171090 132552 171096
rect 132512 137986 132540 171090
rect 133892 137986 133920 173878
rect 136560 173866 136680 173894
rect 136652 172582 136680 173866
rect 136640 172576 136692 172582
rect 136640 172518 136692 172524
rect 135260 171964 135312 171970
rect 135260 171906 135312 171912
rect 135272 151814 135300 171906
rect 136744 171154 136772 174964
rect 142080 174894 142108 178599
rect 144104 174962 144132 178871
rect 153936 178696 153988 178702
rect 153988 178644 154436 178650
rect 153936 178638 154436 178644
rect 153948 178622 154436 178638
rect 145470 177440 145526 177449
rect 145470 177375 145526 177384
rect 144460 175568 144512 175574
rect 144460 175510 144512 175516
rect 144092 174956 144144 174962
rect 144092 174898 144144 174904
rect 142068 174888 142120 174894
rect 142068 174830 142120 174836
rect 137284 173936 137336 173942
rect 137336 173884 137586 173890
rect 137284 173878 137586 173884
rect 137296 173862 137586 173878
rect 138676 171970 138704 173196
rect 139596 173182 139702 173210
rect 138664 171964 138716 171970
rect 138664 171906 138716 171912
rect 136732 171148 136784 171154
rect 136732 171090 136784 171096
rect 138020 171148 138072 171154
rect 138020 171090 138072 171096
rect 138032 151814 138060 171090
rect 135272 151786 135484 151814
rect 138032 151786 138612 151814
rect 135456 137986 135484 151786
rect 137744 139732 137796 139738
rect 137744 139674 137796 139680
rect 137756 137986 137784 139674
rect 124508 137958 124936 137986
rect 126072 137958 126500 137986
rect 127636 137958 128064 137986
rect 129200 137958 129628 137986
rect 131132 137958 131192 137986
rect 132512 137958 132756 137986
rect 133892 137958 134320 137986
rect 135456 137958 135884 137986
rect 137448 137958 137784 137986
rect 138584 137986 138612 151786
rect 139596 139738 139624 173182
rect 140792 171154 140820 173196
rect 140780 171148 140832 171154
rect 140780 171090 140832 171096
rect 142264 140758 142292 173196
rect 142526 172952 142582 172961
rect 142526 172887 142582 172896
rect 142436 166320 142488 166326
rect 142436 166262 142488 166268
rect 142448 142154 142476 166262
rect 142356 142126 142476 142154
rect 140688 140752 140740 140758
rect 140688 140694 140740 140700
rect 142252 140752 142304 140758
rect 142252 140694 142304 140700
rect 139584 139732 139636 139738
rect 139584 139674 139636 139680
rect 140700 137986 140728 140694
rect 142356 139482 142384 142126
rect 142540 140282 142568 172887
rect 142632 166326 142660 173196
rect 142620 166320 142672 166326
rect 142620 166262 142672 166268
rect 143644 161474 143672 173196
rect 143552 161446 143672 161474
rect 142528 140276 142580 140282
rect 142528 140218 142580 140224
rect 138584 137958 139012 137986
rect 140576 137958 140728 137986
rect 142080 139454 142384 139482
rect 142080 137986 142108 139454
rect 143552 137986 143580 161446
rect 144472 140350 144500 175510
rect 144460 140344 144512 140350
rect 144460 140286 144512 140292
rect 144932 137986 144960 173196
rect 145484 171902 145512 177375
rect 149244 176656 149296 176662
rect 149244 176598 149296 176604
rect 149256 175817 149284 176598
rect 154408 176458 154436 178622
rect 158824 176497 158852 179318
rect 158810 176488 158866 176497
rect 154396 176452 154448 176458
rect 158810 176423 158866 176432
rect 154396 176394 154448 176400
rect 160468 175976 160520 175982
rect 160468 175918 160520 175924
rect 159180 175908 159232 175914
rect 159180 175850 159232 175856
rect 159088 175840 159140 175846
rect 149242 175808 149298 175817
rect 159192 175817 159220 175850
rect 159088 175782 159140 175788
rect 159178 175808 159234 175817
rect 149242 175743 149298 175752
rect 149336 175704 149388 175710
rect 149336 175646 149388 175652
rect 148692 175568 148744 175574
rect 148692 175510 148744 175516
rect 148704 175273 148732 175510
rect 149348 175409 149376 175646
rect 159100 175409 159128 175782
rect 159178 175743 159234 175752
rect 149334 175400 149390 175409
rect 149334 175335 149390 175344
rect 159086 175400 159142 175409
rect 159086 175335 159142 175344
rect 148690 175264 148746 175273
rect 148690 175199 148746 175208
rect 154578 175264 154634 175273
rect 154634 175222 154974 175250
rect 154578 175199 154634 175208
rect 145472 171896 145524 171902
rect 145472 171838 145524 171844
rect 146312 151814 146340 173196
rect 146680 161474 146708 173196
rect 147600 161474 147628 173196
rect 149348 170066 149376 173196
rect 149336 170060 149388 170066
rect 149336 170002 149388 170008
rect 149624 161474 149652 173196
rect 150440 170060 150492 170066
rect 150440 170002 150492 170008
rect 146496 161446 146708 161474
rect 147508 161446 147628 161474
rect 149532 161446 149652 161474
rect 146312 151786 146432 151814
rect 146404 137986 146432 151786
rect 146496 139806 146524 161446
rect 146484 139800 146536 139806
rect 146484 139742 146536 139748
rect 147508 139738 147536 161446
rect 148048 139800 148100 139806
rect 148048 139742 148100 139748
rect 147496 139732 147548 139738
rect 147496 139674 147548 139680
rect 148060 137986 148088 139742
rect 149532 139670 149560 161446
rect 150452 139754 150480 170002
rect 150636 161474 150664 173196
rect 152384 170338 152412 173196
rect 152372 170332 152424 170338
rect 152372 170274 152424 170280
rect 152660 161474 152688 173196
rect 150544 161446 150664 161474
rect 152476 161446 152688 161474
rect 153488 173182 153686 173210
rect 150544 140554 150572 161446
rect 150532 140548 150584 140554
rect 150532 140490 150584 140496
rect 149612 139732 149664 139738
rect 150452 139726 151124 139754
rect 152476 139738 152504 161446
rect 153488 139806 153516 173182
rect 158442 172952 158498 172961
rect 158442 172887 158498 172896
rect 157984 171896 158036 171902
rect 157984 171838 158036 171844
rect 156512 170332 156564 170338
rect 156512 170274 156564 170280
rect 154486 169552 154542 169561
rect 154486 169487 154542 169496
rect 154500 152522 154528 169487
rect 154488 152516 154540 152522
rect 154488 152458 154540 152464
rect 154580 140548 154632 140554
rect 154580 140490 154632 140496
rect 153476 139800 153528 139806
rect 153476 139742 153528 139748
rect 149612 139674 149664 139680
rect 149520 139664 149572 139670
rect 149520 139606 149572 139612
rect 149624 137986 149652 139674
rect 151096 137986 151124 139726
rect 152464 139732 152516 139738
rect 152464 139674 152516 139680
rect 152740 139664 152792 139670
rect 152740 139606 152792 139612
rect 152752 137986 152780 139606
rect 154592 137986 154620 140490
rect 156524 137986 156552 170274
rect 157996 145654 158024 171838
rect 157984 145648 158036 145654
rect 157984 145590 158036 145596
rect 157432 139732 157484 139738
rect 157432 139674 157484 139680
rect 142080 137958 142140 137986
rect 143552 137958 143704 137986
rect 144932 137958 145268 137986
rect 146404 137958 146832 137986
rect 148060 137958 148396 137986
rect 149624 137958 149960 137986
rect 151096 137958 151524 137986
rect 152752 137958 153088 137986
rect 154592 137958 154652 137986
rect 156216 137958 156552 137986
rect 157444 137986 157472 139674
rect 158456 138990 158484 172887
rect 160480 172514 160508 175918
rect 163596 175908 163648 175914
rect 163596 175850 163648 175856
rect 162492 175840 162544 175846
rect 162492 175782 162544 175788
rect 163608 175794 163636 175850
rect 164238 175808 164294 175817
rect 161480 174548 161532 174554
rect 161480 174490 161532 174496
rect 160468 172508 160520 172514
rect 160468 172450 160520 172456
rect 161492 151814 161520 174490
rect 162504 172938 162532 175782
rect 163608 175766 164238 175794
rect 164238 175743 164294 175752
rect 166998 175808 167054 175817
rect 166998 175743 167054 175752
rect 162504 172910 162900 172938
rect 162124 172508 162176 172514
rect 162124 172450 162176 172456
rect 162136 160750 162164 172450
rect 162872 166994 162900 172910
rect 162872 166966 163176 166994
rect 162124 160744 162176 160750
rect 162124 160686 162176 160692
rect 163148 151814 163176 166966
rect 161492 151786 162072 151814
rect 163148 151786 163452 151814
rect 160560 140344 160612 140350
rect 160560 140286 160612 140292
rect 158996 139800 159048 139806
rect 158996 139742 159048 139748
rect 158444 138984 158496 138990
rect 158444 138926 158496 138932
rect 159008 137986 159036 139742
rect 160572 137986 160600 140286
rect 162044 137986 162072 151786
rect 163424 138122 163452 151786
rect 163516 140350 163544 175100
rect 163608 151814 163636 173196
rect 164528 173182 164634 173210
rect 163608 151786 163728 151814
rect 163700 140486 163728 151786
rect 163688 140480 163740 140486
rect 163688 140422 163740 140428
rect 164528 140418 164556 173182
rect 165436 172984 165488 172990
rect 165436 172926 165488 172932
rect 164976 145648 165028 145654
rect 164976 145590 165028 145596
rect 164988 143546 165016 145590
rect 164976 143540 165028 143546
rect 164976 143482 165028 143488
rect 164516 140412 164568 140418
rect 164516 140354 164568 140360
rect 163504 140344 163556 140350
rect 163504 140286 163556 140292
rect 163424 138094 163636 138122
rect 163608 137986 163636 138094
rect 165448 137986 165476 172926
rect 167012 137986 167040 175743
rect 170416 153950 170444 184826
rect 179512 162920 179564 162926
rect 179512 162862 179564 162868
rect 179420 160744 179472 160750
rect 179420 160686 179472 160692
rect 171138 157992 171194 158001
rect 171138 157927 171194 157936
rect 170404 153944 170456 153950
rect 170404 153886 170456 153892
rect 169760 152516 169812 152522
rect 169760 152458 169812 152464
rect 169772 151814 169800 152458
rect 171152 151814 171180 157927
rect 172520 153944 172572 153950
rect 172520 153886 172572 153892
rect 169772 151786 169892 151814
rect 171152 151786 171456 151814
rect 168380 143540 168432 143546
rect 168380 143482 168432 143488
rect 168392 137986 168420 143482
rect 169864 137986 169892 151786
rect 171428 137986 171456 151786
rect 172532 150550 172560 153886
rect 172520 150544 172572 150550
rect 172520 150486 172572 150492
rect 176568 150544 176620 150550
rect 176568 150486 176620 150492
rect 176580 149002 176608 150486
rect 176580 148974 176700 149002
rect 176672 146266 176700 148974
rect 176660 146260 176712 146266
rect 176660 146202 176712 146208
rect 178684 146260 178736 146266
rect 178684 146202 178736 146208
rect 174636 140480 174688 140486
rect 174636 140422 174688 140428
rect 173072 140276 173124 140282
rect 173072 140218 173124 140224
rect 173084 137986 173112 140218
rect 174648 137986 174676 140422
rect 176200 140412 176252 140418
rect 176200 140354 176252 140360
rect 176212 137986 176240 140354
rect 178040 140344 178092 140350
rect 178040 140286 178092 140292
rect 178052 137986 178080 140286
rect 178696 140010 178724 146202
rect 178684 140004 178736 140010
rect 178684 139946 178736 139952
rect 157444 137958 157780 137986
rect 159008 137958 159344 137986
rect 160572 137958 160908 137986
rect 162044 137958 162472 137986
rect 163608 137958 164036 137986
rect 165448 137958 165600 137986
rect 167012 137958 167164 137986
rect 168392 137958 168728 137986
rect 169864 137958 170292 137986
rect 171428 137958 171856 137986
rect 173084 137958 173420 137986
rect 174648 137958 174984 137986
rect 176212 137958 176548 137986
rect 178052 137958 178112 137986
rect 179432 111897 179460 160686
rect 179524 131753 179552 162862
rect 179696 140004 179748 140010
rect 179696 139946 179748 139952
rect 179604 138848 179656 138854
rect 179604 138790 179656 138796
rect 179510 131744 179566 131753
rect 179510 131679 179566 131688
rect 179616 118289 179644 138790
rect 179708 137970 179736 139946
rect 179696 137964 179748 137970
rect 179696 137906 179748 137912
rect 179602 118280 179658 118289
rect 179602 118215 179658 118224
rect 179418 111888 179474 111897
rect 179418 111823 179474 111832
rect 120644 103486 120764 103514
rect 120644 101833 120672 103486
rect 120630 101824 120686 101833
rect 120630 101759 120686 101768
rect 120908 98728 120960 98734
rect 120908 98670 120960 98676
rect 119250 97336 119306 97345
rect 119250 97271 119306 97280
rect 120816 95192 120868 95198
rect 120816 95134 120868 95140
rect 118882 93800 118938 93809
rect 118882 93735 118938 93744
rect 118790 85368 118846 85377
rect 118790 85303 118846 85312
rect 120828 84946 120856 95134
rect 120920 85066 120948 98670
rect 120908 85060 120960 85066
rect 120908 85002 120960 85008
rect 120828 84918 121040 84946
rect 120908 84856 120960 84862
rect 120908 84798 120960 84804
rect 120724 84244 120776 84250
rect 120724 84186 120776 84192
rect 120630 81560 120686 81569
rect 120630 81495 120686 81504
rect 117964 81456 118016 81462
rect 117964 81398 118016 81404
rect 118514 80200 118570 80209
rect 118514 80135 118570 80144
rect 118422 78704 118478 78713
rect 118422 78639 118478 78648
rect 116676 77104 116728 77110
rect 116676 77046 116728 77052
rect 3790 76599 3846 76608
rect 4988 76628 5040 76634
rect 4988 76570 5040 76576
rect 110420 75404 110472 75410
rect 110420 75346 110472 75352
rect 57244 75336 57296 75342
rect 57244 75278 57296 75284
rect 46204 75268 46256 75274
rect 46204 75210 46256 75216
rect 22744 75200 22796 75206
rect 22744 75142 22796 75148
rect 20718 73944 20774 73953
rect 20718 73879 20774 73888
rect 16580 72548 16632 72554
rect 16580 72490 16632 72496
rect 6920 72480 6972 72486
rect 6920 72422 6972 72428
rect 3606 58576 3662 58585
rect 3606 58511 3662 58520
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 3516 33040 3568 33046
rect 3516 32982 3568 32988
rect 3528 32473 3556 32982
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3516 23248 3568 23254
rect 3516 23190 3568 23196
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 2792 16546 2912 16574
rect 2884 480 2912 16546
rect 3528 6497 3556 23190
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 4172 16574 4200 18566
rect 6932 16574 6960 72422
rect 16592 16574 16620 72490
rect 20732 16574 20760 73879
rect 4172 16546 5304 16574
rect 6932 16546 7696 16574
rect 16592 16546 17080 16574
rect 20732 16546 21864 16574
rect 3514 6488 3570 6497
rect 3514 6423 3570 6432
rect 4066 3360 4122 3369
rect 4066 3295 4122 3304
rect 4080 480 4108 3295
rect 5276 480 5304 16546
rect 6460 7676 6512 7682
rect 6460 7618 6512 7624
rect 6472 480 6500 7618
rect 7668 480 7696 16546
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8772 480 8800 4762
rect 9968 480 9996 8978
rect 13544 4956 13596 4962
rect 13544 4898 13596 4904
rect 11152 4888 11204 4894
rect 11152 4830 11204 4836
rect 11164 480 11192 4830
rect 12348 4004 12400 4010
rect 12348 3946 12400 3952
rect 12360 480 12388 3946
rect 13556 480 13584 4898
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 15846
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 15948 480 15976 5170
rect 17052 480 17080 16546
rect 18236 7608 18288 7614
rect 18236 7550 18288 7556
rect 18248 480 18276 7550
rect 20626 6216 20682 6225
rect 20626 6151 20682 6160
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19444 480 19472 4966
rect 20640 480 20668 6151
rect 21836 480 21864 16546
rect 22756 7682 22784 75142
rect 44180 73908 44232 73914
rect 44180 73850 44232 73856
rect 30380 73840 30432 73846
rect 30380 73782 30432 73788
rect 26240 71052 26292 71058
rect 26240 70994 26292 71000
rect 25320 10328 25372 10334
rect 25320 10270 25372 10276
rect 22744 7676 22796 7682
rect 22744 7618 22796 7624
rect 24216 6180 24268 6186
rect 24216 6122 24268 6128
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 23032 480 23060 3470
rect 24228 480 24256 6122
rect 25332 480 25360 10270
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 70994
rect 30392 16574 30420 73782
rect 42800 72616 42852 72622
rect 42800 72558 42852 72564
rect 35898 71088 35954 71097
rect 35898 71023 35954 71032
rect 30392 16546 30880 16574
rect 27712 7676 27764 7682
rect 27712 7618 27764 7624
rect 27724 480 27752 7618
rect 30104 5160 30156 5166
rect 30104 5102 30156 5108
rect 28908 5092 28960 5098
rect 28908 5034 28960 5040
rect 28920 480 28948 5034
rect 30116 480 30144 5102
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31944 14476 31996 14482
rect 31944 14418 31996 14424
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 14418
rect 34796 9104 34848 9110
rect 34796 9046 34848 9052
rect 33600 6248 33652 6254
rect 33600 6190 33652 6196
rect 33612 480 33640 6190
rect 34808 480 34836 9046
rect 35912 3466 35940 71023
rect 35992 44872 36044 44878
rect 35992 44814 36044 44820
rect 35900 3460 35952 3466
rect 35900 3402 35952 3408
rect 36004 480 36032 44814
rect 38660 17264 38712 17270
rect 38660 17206 38712 17212
rect 38672 16574 38700 17206
rect 38672 16546 39160 16574
rect 38382 8936 38438 8945
rect 38382 8871 38438 8880
rect 36820 3460 36872 3466
rect 36820 3402 36872 3408
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 36832 354 36860 3402
rect 38396 480 38424 8871
rect 37158 354 37270 480
rect 36832 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 41878 9072 41934 9081
rect 41878 9007 41934 9016
rect 40682 6352 40738 6361
rect 40682 6287 40738 6296
rect 40696 480 40724 6287
rect 41892 480 41920 9007
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 39550 -960 39662 326
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 42812 354 42840 72558
rect 44192 16574 44220 73850
rect 45560 21412 45612 21418
rect 45560 21354 45612 21360
rect 45572 16574 45600 21354
rect 44192 16546 45048 16574
rect 45572 16546 46152 16574
rect 44272 6316 44324 6322
rect 44272 6258 44324 6264
rect 44284 480 44312 6258
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46124 3482 46152 16546
rect 46216 5234 46244 75210
rect 51080 72752 51132 72758
rect 51080 72694 51132 72700
rect 46940 71120 46992 71126
rect 46940 71062 46992 71068
rect 46952 16574 46980 71062
rect 46952 16546 47440 16574
rect 46204 5228 46256 5234
rect 46204 5170 46256 5176
rect 46124 3454 46704 3482
rect 46676 480 46704 3454
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 50160 9172 50212 9178
rect 50160 9114 50212 9120
rect 48964 6384 49016 6390
rect 48964 6326 49016 6332
rect 48976 480 49004 6326
rect 50172 480 50200 9114
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 47830 -960 47942 326
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 72694
rect 53838 72584 53894 72593
rect 53838 72519 53894 72528
rect 52460 22840 52512 22846
rect 52460 22782 52512 22788
rect 52472 16574 52500 22782
rect 53852 16574 53880 72519
rect 52472 16546 52592 16574
rect 53852 16546 54984 16574
rect 52564 480 52592 16546
rect 53748 9240 53800 9246
rect 53748 9182 53800 9188
rect 53760 480 53788 9182
rect 54956 480 54984 16546
rect 57256 10334 57284 75278
rect 102140 74180 102192 74186
rect 102140 74122 102192 74128
rect 93860 74112 93912 74118
rect 93860 74054 93912 74060
rect 86960 74044 87012 74050
rect 86960 73986 87012 73992
rect 69020 73976 69072 73982
rect 69020 73918 69072 73924
rect 57978 72720 58034 72729
rect 57978 72655 58034 72664
rect 60740 72684 60792 72690
rect 57992 16574 58020 72655
rect 60740 72626 60792 72632
rect 57992 16546 58480 16574
rect 57244 10328 57296 10334
rect 57244 10270 57296 10276
rect 57242 9208 57298 9217
rect 57242 9143 57298 9152
rect 56046 7576 56102 7585
rect 56046 7511 56102 7520
rect 56060 480 56088 7511
rect 57256 480 57284 9143
rect 58452 480 58480 16546
rect 59636 5228 59688 5234
rect 59636 5170 59688 5176
rect 59648 480 59676 5170
rect 60752 3466 60780 72626
rect 64880 71188 64932 71194
rect 64880 71130 64932 71136
rect 64892 16574 64920 71130
rect 69032 16574 69060 73918
rect 75920 71256 75972 71262
rect 75920 71198 75972 71204
rect 70400 19984 70452 19990
rect 70400 19926 70452 19932
rect 70412 16574 70440 19926
rect 64892 16546 65104 16574
rect 69032 16546 69888 16574
rect 70412 16546 71544 16574
rect 64328 10396 64380 10402
rect 64328 10338 64380 10344
rect 60832 10328 60884 10334
rect 60832 10270 60884 10276
rect 60740 3460 60792 3466
rect 60740 3402 60792 3408
rect 60844 480 60872 10270
rect 63224 6452 63276 6458
rect 63224 6394 63276 6400
rect 61660 3460 61712 3466
rect 61660 3402 61712 3408
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61672 354 61700 3402
rect 63236 480 63264 6394
rect 64340 480 64368 10338
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 67640 10464 67692 10470
rect 67640 10406 67692 10412
rect 66720 6520 66772 6526
rect 66720 6462 66772 6468
rect 66732 480 66760 6462
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 10406
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 69124 480 69152 3538
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71516 480 71544 16546
rect 74998 11656 75054 11665
rect 74998 11591 75054 11600
rect 73802 6488 73858 6497
rect 73802 6423 73858 6432
rect 72608 3664 72660 3670
rect 72608 3606 72660 3612
rect 72620 480 72648 3606
rect 73816 480 73844 6423
rect 75012 480 75040 11591
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 71198
rect 86972 16574 87000 73986
rect 89718 71224 89774 71233
rect 89718 71159 89774 71168
rect 88340 36576 88392 36582
rect 88340 36518 88392 36524
rect 88352 16574 88380 36518
rect 89732 16574 89760 71159
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 81624 10600 81676 10606
rect 81624 10542 81676 10548
rect 78128 10532 78180 10538
rect 78128 10474 78180 10480
rect 77392 7744 77444 7750
rect 77392 7686 77444 7692
rect 77404 480 77432 7686
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 10474
rect 80888 7812 80940 7818
rect 80888 7754 80940 7760
rect 79692 3732 79744 3738
rect 79692 3674 79744 3680
rect 79704 480 79732 3674
rect 80900 480 80928 7754
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 78558 -960 78670 326
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 81636 354 81664 10542
rect 84476 7880 84528 7886
rect 84476 7822 84528 7828
rect 83280 3800 83332 3806
rect 83280 3742 83332 3748
rect 83292 480 83320 3742
rect 84488 480 84516 7822
rect 85672 5296 85724 5302
rect 85672 5238 85724 5244
rect 85684 480 85712 5238
rect 86868 3868 86920 3874
rect 86868 3810 86920 3816
rect 86880 480 86908 3810
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87524 354 87552 16546
rect 88154 6624 88210 6633
rect 88154 6559 88210 6568
rect 88168 3534 88196 6559
rect 88156 3528 88208 3534
rect 88156 3470 88208 3476
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 92478 10296 92534 10305
rect 92478 10231 92534 10240
rect 91558 7712 91614 7721
rect 91558 7647 91614 7656
rect 91572 480 91600 7647
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 10231
rect 93872 3534 93900 74054
rect 93952 71324 94004 71330
rect 93952 71266 94004 71272
rect 93860 3528 93912 3534
rect 93860 3470 93912 3476
rect 93964 480 93992 71266
rect 95240 55888 95292 55894
rect 95240 55830 95292 55836
rect 95252 16574 95280 55830
rect 95252 16546 95832 16574
rect 94780 3528 94832 3534
rect 94780 3470 94832 3476
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 3470
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 99840 10668 99892 10674
rect 99840 10610 99892 10616
rect 98644 7948 98696 7954
rect 98644 7890 98696 7896
rect 97448 5364 97500 5370
rect 97448 5306 97500 5312
rect 97460 480 97488 5306
rect 98656 480 98684 7890
rect 99852 480 99880 10610
rect 102152 6914 102180 74122
rect 107660 72820 107712 72826
rect 107660 72762 107712 72768
rect 102232 54528 102284 54534
rect 102232 54470 102284 54476
rect 102244 16574 102272 54470
rect 106280 20052 106332 20058
rect 106280 19994 106332 20000
rect 106292 16574 106320 19994
rect 107672 16574 107700 72762
rect 102244 16546 103376 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102152 6886 102272 6914
rect 101036 5432 101088 5438
rect 101036 5374 101088 5380
rect 101048 480 101076 5374
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 105728 8084 105780 8090
rect 105728 8026 105780 8032
rect 104532 8016 104584 8022
rect 104532 7958 104584 7964
rect 104544 480 104572 7958
rect 105740 480 105768 8026
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 109314 9344 109370 9353
rect 109314 9279 109370 9288
rect 109328 480 109356 9279
rect 110432 3534 110460 75346
rect 111798 74080 111854 74089
rect 111798 74015 111854 74024
rect 111812 16574 111840 74015
rect 114560 69692 114612 69698
rect 114560 69634 114612 69640
rect 114572 16574 114600 69634
rect 118436 22778 118464 78639
rect 118528 60722 118556 80135
rect 120644 78674 120672 81495
rect 120632 78668 120684 78674
rect 120632 78610 120684 78616
rect 118792 78260 118844 78266
rect 118792 78202 118844 78208
rect 118804 77246 118832 78202
rect 119804 77648 119856 77654
rect 119804 77590 119856 77596
rect 118792 77240 118844 77246
rect 118792 77182 118844 77188
rect 119816 75274 119844 77590
rect 120736 77042 120764 84186
rect 120816 81388 120868 81394
rect 120816 81330 120868 81336
rect 120724 77036 120776 77042
rect 120724 76978 120776 76984
rect 119804 75268 119856 75274
rect 119804 75210 119856 75216
rect 120724 74724 120776 74730
rect 120724 74666 120776 74672
rect 118700 71392 118752 71398
rect 118700 71334 118752 71340
rect 118516 60716 118568 60722
rect 118516 60658 118568 60664
rect 118424 22772 118476 22778
rect 118424 22714 118476 22720
rect 118712 16574 118740 71334
rect 120080 40316 120132 40322
rect 120080 40258 120132 40264
rect 120092 16574 120120 40258
rect 120736 17270 120764 74666
rect 120828 73642 120856 81330
rect 120920 73710 120948 84798
rect 121012 74254 121040 84918
rect 178960 79348 179012 79354
rect 178960 79290 179012 79296
rect 124772 78668 124996 78674
rect 124824 78646 124996 78668
rect 124772 78610 124824 78616
rect 124968 78606 124996 78646
rect 174544 78668 174596 78674
rect 174544 78610 174596 78616
rect 124956 78600 125008 78606
rect 124956 78542 125008 78548
rect 174340 78254 174492 78282
rect 122104 78124 122156 78130
rect 122104 78066 122156 78072
rect 125428 78118 125580 78146
rect 121644 77852 121696 77858
rect 121644 77794 121696 77800
rect 121368 76492 121420 76498
rect 121368 76434 121420 76440
rect 121092 75880 121144 75886
rect 121092 75822 121144 75828
rect 121000 74248 121052 74254
rect 121000 74190 121052 74196
rect 120908 73704 120960 73710
rect 120908 73646 120960 73652
rect 120816 73636 120868 73642
rect 120816 73578 120868 73584
rect 121104 70394 121132 75822
rect 121380 73953 121408 76434
rect 121366 73944 121422 73953
rect 121366 73879 121422 73888
rect 121460 72888 121512 72894
rect 121460 72830 121512 72836
rect 120828 70366 121132 70394
rect 120828 21418 120856 70366
rect 120816 21412 120868 21418
rect 120816 21354 120868 21360
rect 120724 17264 120776 17270
rect 120724 17206 120776 17212
rect 121472 16574 121500 72830
rect 121656 72486 121684 77794
rect 121644 72480 121696 72486
rect 121644 72422 121696 72428
rect 111812 16546 112392 16574
rect 114572 16546 114784 16574
rect 118712 16546 118832 16574
rect 120092 16546 120672 16574
rect 121472 16546 122052 16574
rect 110510 10432 110566 10441
rect 110510 10367 110566 10376
rect 110420 3528 110472 3534
rect 110420 3470 110472 3476
rect 110524 480 110552 10367
rect 111616 3528 111668 3534
rect 111616 3470 111668 3476
rect 111628 480 111656 3470
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114006 10568 114062 10577
rect 114006 10503 114062 10512
rect 114020 480 114048 10503
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 117320 11756 117372 11762
rect 117320 11698 117372 11704
rect 116400 9308 116452 9314
rect 116400 9250 116452 9256
rect 116412 480 116440 9250
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 11698
rect 118804 480 118832 16546
rect 119896 4140 119948 4146
rect 119896 4082 119948 4088
rect 119908 480 119936 4082
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122024 3482 122052 16546
rect 122116 6186 122144 78066
rect 124864 78056 124916 78062
rect 124864 77998 124916 78004
rect 124772 77988 124824 77994
rect 124772 77930 124824 77936
rect 123758 77888 123814 77897
rect 123758 77823 123814 77832
rect 123772 75206 123800 77823
rect 124784 77217 124812 77930
rect 124770 77208 124826 77217
rect 124770 77143 124826 77152
rect 124772 76764 124824 76770
rect 124772 76706 124824 76712
rect 123760 75200 123812 75206
rect 123760 75142 123812 75148
rect 123484 74996 123536 75002
rect 123484 74938 123536 74944
rect 122840 74452 122892 74458
rect 122840 74394 122892 74400
rect 122196 73908 122248 73914
rect 122196 73850 122248 73856
rect 122208 14482 122236 73850
rect 122852 16574 122880 74394
rect 123496 40322 123524 74938
rect 124784 73982 124812 76706
rect 124772 73976 124824 73982
rect 124772 73918 124824 73924
rect 124220 72412 124272 72418
rect 124220 72354 124272 72360
rect 123484 40316 123536 40322
rect 123484 40258 123536 40264
rect 122852 16546 123064 16574
rect 122196 14476 122248 14482
rect 122196 14418 122248 14424
rect 122104 6180 122156 6186
rect 122104 6122 122156 6128
rect 122024 3454 122328 3482
rect 122300 480 122328 3454
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124232 8974 124260 72354
rect 124220 8968 124272 8974
rect 124220 8910 124272 8916
rect 124876 5030 124904 77998
rect 125324 77920 125376 77926
rect 125324 77862 125376 77868
rect 125048 77512 125100 77518
rect 125048 77454 125100 77460
rect 124956 74520 125008 74526
rect 124956 74462 125008 74468
rect 124864 5024 124916 5030
rect 124864 4966 124916 4972
rect 124968 4146 124996 74462
rect 125060 15910 125088 77454
rect 125232 75812 125284 75818
rect 125232 75754 125284 75760
rect 125140 74860 125192 74866
rect 125140 74802 125192 74808
rect 125152 36582 125180 74802
rect 125244 54534 125272 75754
rect 125336 75177 125364 77862
rect 125322 75168 125378 75177
rect 125322 75103 125378 75112
rect 125324 75064 125376 75070
rect 125324 75006 125376 75012
rect 125336 55894 125364 75006
rect 125428 72418 125456 78118
rect 125658 77908 125686 78132
rect 125520 77880 125686 77908
rect 125520 73817 125548 77880
rect 125750 77840 125778 78132
rect 125842 77926 125870 78132
rect 125830 77920 125882 77926
rect 125830 77862 125882 77868
rect 125704 77812 125778 77840
rect 125506 73808 125562 73817
rect 125506 73743 125562 73752
rect 125704 72457 125732 77812
rect 125934 77772 125962 78132
rect 126026 77897 126054 78132
rect 126012 77888 126068 77897
rect 126118 77858 126146 78132
rect 126210 77858 126238 78132
rect 126302 77897 126330 78132
rect 126288 77888 126344 77897
rect 126012 77823 126068 77832
rect 126106 77852 126158 77858
rect 126106 77794 126158 77800
rect 126198 77852 126250 77858
rect 126394 77858 126422 78132
rect 126288 77823 126344 77832
rect 126382 77852 126434 77858
rect 126198 77794 126250 77800
rect 126382 77794 126434 77800
rect 125842 77744 125962 77772
rect 126242 77752 126298 77761
rect 125842 77636 125870 77744
rect 126152 77716 126204 77722
rect 126242 77687 126298 77696
rect 126336 77716 126388 77722
rect 126152 77658 126204 77664
rect 125842 77608 126008 77636
rect 125876 77444 125928 77450
rect 125876 77386 125928 77392
rect 125784 76356 125836 76362
rect 125784 76298 125836 76304
rect 125690 72448 125746 72457
rect 125416 72412 125468 72418
rect 125690 72383 125746 72392
rect 125416 72354 125468 72360
rect 125324 55888 125376 55894
rect 125324 55830 125376 55836
rect 125232 54528 125284 54534
rect 125232 54470 125284 54476
rect 125140 36576 125192 36582
rect 125140 36518 125192 36524
rect 125048 15904 125100 15910
rect 125048 15846 125100 15852
rect 125796 4826 125824 76298
rect 125888 74534 125916 77386
rect 125980 76242 126008 77608
rect 126164 76362 126192 77658
rect 126152 76356 126204 76362
rect 126152 76298 126204 76304
rect 125980 76214 126192 76242
rect 126060 76152 126112 76158
rect 126060 76094 126112 76100
rect 125888 74506 126008 74534
rect 125876 73568 125928 73574
rect 125876 73510 125928 73516
rect 125888 4894 125916 73510
rect 125980 7614 126008 74506
rect 126072 9042 126100 76094
rect 126164 18630 126192 76214
rect 126256 76158 126284 77687
rect 126336 77658 126388 77664
rect 126244 76152 126296 76158
rect 126244 76094 126296 76100
rect 126348 73574 126376 77658
rect 126486 77636 126514 78132
rect 126440 77608 126514 77636
rect 126336 73568 126388 73574
rect 126336 73510 126388 73516
rect 126336 72548 126388 72554
rect 126336 72490 126388 72496
rect 126242 71904 126298 71913
rect 126242 71839 126298 71848
rect 126152 18624 126204 18630
rect 126152 18566 126204 18572
rect 126060 9036 126112 9042
rect 126060 8978 126112 8984
rect 125968 7608 126020 7614
rect 125968 7550 126020 7556
rect 125876 4888 125928 4894
rect 125876 4830 125928 4836
rect 125784 4820 125836 4826
rect 125784 4762 125836 4768
rect 124956 4140 125008 4146
rect 124956 4082 125008 4088
rect 125876 4140 125928 4146
rect 125876 4082 125928 4088
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 124692 480 124720 3470
rect 125888 480 125916 4082
rect 126256 3670 126284 71839
rect 126348 10402 126376 72490
rect 126336 10396 126388 10402
rect 126336 10338 126388 10344
rect 126440 4010 126468 77608
rect 126578 77568 126606 78132
rect 126670 77722 126698 78132
rect 126658 77716 126710 77722
rect 126658 77658 126710 77664
rect 126762 77602 126790 78132
rect 126854 77636 126882 78132
rect 126946 77926 126974 78132
rect 127038 77926 127066 78132
rect 127130 77926 127158 78132
rect 127222 77926 127250 78132
rect 126934 77920 126986 77926
rect 126934 77862 126986 77868
rect 127026 77920 127078 77926
rect 127026 77862 127078 77868
rect 127118 77920 127170 77926
rect 127118 77862 127170 77868
rect 127210 77920 127262 77926
rect 127210 77862 127262 77868
rect 127314 77858 127342 78132
rect 127406 77858 127434 78132
rect 127498 77926 127526 78132
rect 127486 77920 127538 77926
rect 127590 77897 127618 78132
rect 127682 77926 127710 78132
rect 127774 77926 127802 78132
rect 127866 77926 127894 78132
rect 127958 77926 127986 78132
rect 127670 77920 127722 77926
rect 127486 77862 127538 77868
rect 127576 77888 127632 77897
rect 127302 77852 127354 77858
rect 127302 77794 127354 77800
rect 127394 77852 127446 77858
rect 127670 77862 127722 77868
rect 127762 77920 127814 77926
rect 127762 77862 127814 77868
rect 127854 77920 127906 77926
rect 127854 77862 127906 77868
rect 127946 77920 127998 77926
rect 128050 77897 128078 78132
rect 128142 77926 128170 78132
rect 128234 77926 128262 78132
rect 128326 77926 128354 78132
rect 128130 77920 128182 77926
rect 127946 77862 127998 77868
rect 128036 77888 128092 77897
rect 127576 77823 127632 77832
rect 128130 77862 128182 77868
rect 128222 77920 128274 77926
rect 128222 77862 128274 77868
rect 128314 77920 128366 77926
rect 128314 77862 128366 77868
rect 128036 77823 128092 77832
rect 127394 77794 127446 77800
rect 127072 77784 127124 77790
rect 127808 77784 127860 77790
rect 127072 77726 127124 77732
rect 127530 77752 127586 77761
rect 126980 77716 127032 77722
rect 126980 77658 127032 77664
rect 126854 77608 126928 77636
rect 126716 77574 126790 77602
rect 126578 77540 126652 77568
rect 126624 76106 126652 77540
rect 126716 77382 126744 77574
rect 126704 77376 126756 77382
rect 126704 77318 126756 77324
rect 126624 76078 126744 76106
rect 126610 75440 126666 75449
rect 126610 75375 126666 75384
rect 126624 72554 126652 75375
rect 126612 72548 126664 72554
rect 126612 72490 126664 72496
rect 126610 71360 126666 71369
rect 126610 71295 126666 71304
rect 126624 71058 126652 71295
rect 126612 71052 126664 71058
rect 126612 70994 126664 71000
rect 126716 69014 126744 76078
rect 126796 75132 126848 75138
rect 126796 75074 126848 75080
rect 126808 74458 126836 75074
rect 126796 74452 126848 74458
rect 126796 74394 126848 74400
rect 126900 72486 126928 77608
rect 126992 76498 127020 77658
rect 126980 76492 127032 76498
rect 126980 76434 127032 76440
rect 127084 76401 127112 77726
rect 127808 77726 127860 77732
rect 127900 77784 127952 77790
rect 127900 77726 127952 77732
rect 127530 77687 127586 77696
rect 127624 77716 127676 77722
rect 127256 77648 127308 77654
rect 127256 77590 127308 77596
rect 127440 77648 127492 77654
rect 127440 77590 127492 77596
rect 127268 76809 127296 77590
rect 127348 77444 127400 77450
rect 127348 77386 127400 77392
rect 127254 76800 127310 76809
rect 127254 76735 127310 76744
rect 127070 76392 127126 76401
rect 127070 76327 127126 76336
rect 127256 76356 127308 76362
rect 127256 76298 127308 76304
rect 127164 74928 127216 74934
rect 127164 74870 127216 74876
rect 127072 73704 127124 73710
rect 127072 73646 127124 73652
rect 127084 73574 127112 73646
rect 127072 73568 127124 73574
rect 127072 73510 127124 73516
rect 126888 72480 126940 72486
rect 126888 72422 126940 72428
rect 126532 68986 126744 69014
rect 126532 4962 126560 68986
rect 127176 6254 127204 74870
rect 127268 7682 127296 76298
rect 127360 9110 127388 77386
rect 127452 75342 127480 77590
rect 127440 75336 127492 75342
rect 127440 75278 127492 75284
rect 127440 75132 127492 75138
rect 127440 75074 127492 75080
rect 127452 44878 127480 75074
rect 127544 73914 127572 77687
rect 127624 77658 127676 77664
rect 127636 76362 127664 77658
rect 127716 77512 127768 77518
rect 127716 77454 127768 77460
rect 127624 76356 127676 76362
rect 127624 76298 127676 76304
rect 127624 76220 127676 76226
rect 127624 76162 127676 76168
rect 127532 73908 127584 73914
rect 127532 73850 127584 73856
rect 127532 73364 127584 73370
rect 127532 73306 127584 73312
rect 127440 44872 127492 44878
rect 127440 44814 127492 44820
rect 127348 9104 127400 9110
rect 127348 9046 127400 9052
rect 127256 7676 127308 7682
rect 127256 7618 127308 7624
rect 127164 6248 127216 6254
rect 127164 6190 127216 6196
rect 127544 5166 127572 73306
rect 127636 71126 127664 76162
rect 127624 71120 127676 71126
rect 127624 71062 127676 71068
rect 127728 64874 127756 77454
rect 127636 64846 127756 64874
rect 127636 9178 127664 64846
rect 127624 9172 127676 9178
rect 127624 9114 127676 9120
rect 127532 5160 127584 5166
rect 127532 5102 127584 5108
rect 127820 5098 127848 77726
rect 127912 73370 127940 77726
rect 127992 77716 128044 77722
rect 127992 77658 128044 77664
rect 128084 77716 128136 77722
rect 128314 77716 128366 77722
rect 128084 77658 128136 77664
rect 128188 77676 128314 77704
rect 128004 73778 128032 77658
rect 128096 74934 128124 77658
rect 128188 75138 128216 77676
rect 128418 77704 128446 78132
rect 128510 77926 128538 78132
rect 128602 77926 128630 78132
rect 128694 77926 128722 78132
rect 128498 77920 128550 77926
rect 128498 77862 128550 77868
rect 128590 77920 128642 77926
rect 128590 77862 128642 77868
rect 128682 77920 128734 77926
rect 128682 77862 128734 77868
rect 128786 77704 128814 78132
rect 128418 77676 128492 77704
rect 128314 77658 128366 77664
rect 128464 76809 128492 77676
rect 128740 77676 128814 77704
rect 128544 77580 128596 77586
rect 128544 77522 128596 77528
rect 128636 77580 128688 77586
rect 128636 77522 128688 77528
rect 128450 76800 128506 76809
rect 128450 76735 128506 76744
rect 128450 76392 128506 76401
rect 128450 76327 128506 76336
rect 128464 75596 128492 76327
rect 128556 75857 128584 77522
rect 128542 75848 128598 75857
rect 128542 75783 128598 75792
rect 128544 75744 128596 75750
rect 128544 75686 128596 75692
rect 128372 75568 128492 75596
rect 128176 75132 128228 75138
rect 128176 75074 128228 75080
rect 128084 74928 128136 74934
rect 128084 74870 128136 74876
rect 128084 74384 128136 74390
rect 128084 74326 128136 74332
rect 127992 73772 128044 73778
rect 127992 73714 128044 73720
rect 128096 73642 128124 74326
rect 128372 73846 128400 75568
rect 128452 74928 128504 74934
rect 128452 74870 128504 74876
rect 128360 73840 128412 73846
rect 128360 73782 128412 73788
rect 128084 73636 128136 73642
rect 128084 73578 128136 73584
rect 127900 73364 127952 73370
rect 127900 73306 127952 73312
rect 128360 73160 128412 73166
rect 128360 73102 128412 73108
rect 128372 6914 128400 73102
rect 128464 10538 128492 74870
rect 128452 10532 128504 10538
rect 128452 10474 128504 10480
rect 128372 6886 128492 6914
rect 127808 5092 127860 5098
rect 127808 5034 127860 5040
rect 126520 4956 126572 4962
rect 126520 4898 126572 4904
rect 126428 4004 126480 4010
rect 126428 3946 126480 3952
rect 126244 3664 126296 3670
rect 126244 3606 126296 3612
rect 126980 3596 127032 3602
rect 126980 3538 127032 3544
rect 126992 480 127020 3538
rect 128174 3360 128230 3369
rect 128174 3295 128230 3304
rect 128188 480 128216 3295
rect 128464 490 128492 6886
rect 128556 6390 128584 75686
rect 128648 74730 128676 77522
rect 128740 75585 128768 77676
rect 128878 77636 128906 78132
rect 128970 77772 128998 78132
rect 129062 77897 129090 78132
rect 129154 77926 129182 78132
rect 129142 77920 129194 77926
rect 129048 77888 129104 77897
rect 129142 77862 129194 77868
rect 129246 77858 129274 78132
rect 129338 77926 129366 78132
rect 129430 77926 129458 78132
rect 129522 77926 129550 78132
rect 129614 77926 129642 78132
rect 129326 77920 129378 77926
rect 129326 77862 129378 77868
rect 129418 77920 129470 77926
rect 129418 77862 129470 77868
rect 129510 77920 129562 77926
rect 129510 77862 129562 77868
rect 129602 77920 129654 77926
rect 129602 77862 129654 77868
rect 129048 77823 129104 77832
rect 129234 77852 129286 77858
rect 129234 77794 129286 77800
rect 129464 77784 129516 77790
rect 128970 77744 129044 77772
rect 128878 77608 128952 77636
rect 128820 77512 128872 77518
rect 128820 77454 128872 77460
rect 128832 76129 128860 77454
rect 128818 76120 128874 76129
rect 128818 76055 128874 76064
rect 128726 75576 128782 75585
rect 128726 75511 128782 75520
rect 128728 75336 128780 75342
rect 128728 75278 128780 75284
rect 128636 74724 128688 74730
rect 128636 74666 128688 74672
rect 128634 74216 128690 74225
rect 128634 74151 128690 74160
rect 128648 74118 128676 74151
rect 128636 74112 128688 74118
rect 128636 74054 128688 74060
rect 128636 72480 128688 72486
rect 128636 72422 128688 72428
rect 128648 9246 128676 72422
rect 128740 22846 128768 75278
rect 128924 74534 128952 77608
rect 129016 75834 129044 77744
rect 129706 77772 129734 78132
rect 129464 77726 129516 77732
rect 129660 77744 129734 77772
rect 129096 77716 129148 77722
rect 129096 77658 129148 77664
rect 129372 77716 129424 77722
rect 129372 77658 129424 77664
rect 129108 76226 129136 77658
rect 129188 77648 129240 77654
rect 129188 77590 129240 77596
rect 129096 76220 129148 76226
rect 129096 76162 129148 76168
rect 129200 75954 129228 77590
rect 129280 77444 129332 77450
rect 129280 77386 129332 77392
rect 129292 77217 129320 77386
rect 129278 77208 129334 77217
rect 129278 77143 129334 77152
rect 129188 75948 129240 75954
rect 129188 75890 129240 75896
rect 129016 75806 129320 75834
rect 129188 75268 129240 75274
rect 129188 75210 129240 75216
rect 128924 74506 129136 74534
rect 129108 73154 129136 74506
rect 128924 73126 129136 73154
rect 128924 72622 128952 73126
rect 128912 72616 128964 72622
rect 128912 72558 128964 72564
rect 129200 70394 129228 75210
rect 129108 70366 129228 70394
rect 128728 22840 128780 22846
rect 128728 22782 128780 22788
rect 129108 10334 129136 70366
rect 129096 10328 129148 10334
rect 129096 10270 129148 10276
rect 128636 9240 128688 9246
rect 128636 9182 128688 9188
rect 128544 6384 128596 6390
rect 128544 6326 128596 6332
rect 129292 6322 129320 75806
rect 129384 75750 129412 77658
rect 129372 75744 129424 75750
rect 129372 75686 129424 75692
rect 129372 75132 129424 75138
rect 129372 75074 129424 75080
rect 129384 72826 129412 75074
rect 129372 72820 129424 72826
rect 129372 72762 129424 72768
rect 129476 72758 129504 77726
rect 129556 77716 129608 77722
rect 129556 77658 129608 77664
rect 129568 75342 129596 77658
rect 129556 75336 129608 75342
rect 129556 75278 129608 75284
rect 129464 72752 129516 72758
rect 129464 72694 129516 72700
rect 129660 72486 129688 77744
rect 129798 77704 129826 78132
rect 129890 77897 129918 78132
rect 129982 77926 130010 78132
rect 129970 77920 130022 77926
rect 129876 77888 129932 77897
rect 129970 77862 130022 77868
rect 129876 77823 129932 77832
rect 129924 77784 129976 77790
rect 130074 77772 130102 78132
rect 130166 77926 130194 78132
rect 130258 77926 130286 78132
rect 130154 77920 130206 77926
rect 130154 77862 130206 77868
rect 130246 77920 130298 77926
rect 130246 77862 130298 77868
rect 130350 77772 130378 78132
rect 129924 77726 129976 77732
rect 130028 77744 130102 77772
rect 130304 77744 130378 77772
rect 129752 77676 129826 77704
rect 129752 76401 129780 77676
rect 129738 76392 129794 76401
rect 129738 76327 129794 76336
rect 129832 76356 129884 76362
rect 129832 76298 129884 76304
rect 129740 74792 129792 74798
rect 129740 74734 129792 74740
rect 129648 72480 129700 72486
rect 129648 72422 129700 72428
rect 129752 70394 129780 74734
rect 129844 72729 129872 76298
rect 129830 72720 129886 72729
rect 129830 72655 129886 72664
rect 129752 70366 129872 70394
rect 129844 64874 129872 70366
rect 129752 64846 129872 64874
rect 129752 16574 129780 64846
rect 129752 16546 129872 16574
rect 129280 6316 129332 6322
rect 129280 6258 129332 6264
rect 129844 3482 129872 16546
rect 129936 5234 129964 77726
rect 130028 77704 130056 77744
rect 130200 77716 130252 77722
rect 130028 77676 130148 77704
rect 130016 77580 130068 77586
rect 130016 77522 130068 77528
rect 130028 76401 130056 77522
rect 130014 76392 130070 76401
rect 130120 76362 130148 77676
rect 130200 77658 130252 77664
rect 130014 76327 130070 76336
rect 130108 76356 130160 76362
rect 130108 76298 130160 76304
rect 130016 76288 130068 76294
rect 130016 76230 130068 76236
rect 130028 6458 130056 76230
rect 130108 75336 130160 75342
rect 130108 75278 130160 75284
rect 130120 6526 130148 75278
rect 130212 75274 130240 77658
rect 130304 76362 130332 77744
rect 130442 77738 130470 78132
rect 130534 77897 130562 78132
rect 130626 77926 130654 78132
rect 130718 77926 130746 78132
rect 130810 77926 130838 78132
rect 130614 77920 130666 77926
rect 130520 77888 130576 77897
rect 130614 77862 130666 77868
rect 130706 77920 130758 77926
rect 130706 77862 130758 77868
rect 130798 77920 130850 77926
rect 130798 77862 130850 77868
rect 130520 77823 130576 77832
rect 130660 77784 130712 77790
rect 130442 77710 130516 77738
rect 130660 77726 130712 77732
rect 130752 77784 130804 77790
rect 130902 77772 130930 78132
rect 130994 77926 131022 78132
rect 130982 77920 131034 77926
rect 130982 77862 131034 77868
rect 131086 77772 131114 78132
rect 131178 77926 131206 78132
rect 131270 77926 131298 78132
rect 131166 77920 131218 77926
rect 131166 77862 131218 77868
rect 131258 77920 131310 77926
rect 131258 77862 131310 77868
rect 130856 77761 130930 77772
rect 130752 77726 130804 77732
rect 130842 77752 130930 77761
rect 130292 76356 130344 76362
rect 130292 76298 130344 76304
rect 130488 76294 130516 77710
rect 130568 77376 130620 77382
rect 130568 77318 130620 77324
rect 130476 76288 130528 76294
rect 130476 76230 130528 76236
rect 130580 75800 130608 77318
rect 130488 75772 130608 75800
rect 130200 75268 130252 75274
rect 130200 75210 130252 75216
rect 130488 74984 130516 75772
rect 130566 75712 130622 75721
rect 130566 75647 130622 75656
rect 130212 74956 130516 74984
rect 130212 10470 130240 74956
rect 130292 74452 130344 74458
rect 130292 74394 130344 74400
rect 130304 19990 130332 74394
rect 130382 71768 130438 71777
rect 130382 71703 130438 71712
rect 130292 19984 130344 19990
rect 130292 19926 130344 19932
rect 130200 10464 130252 10470
rect 130200 10406 130252 10412
rect 130108 6520 130160 6526
rect 130108 6462 130160 6468
rect 130016 6452 130068 6458
rect 130016 6394 130068 6400
rect 129924 5228 129976 5234
rect 129924 5170 129976 5176
rect 130396 3602 130424 71703
rect 130580 16574 130608 75647
rect 130672 75342 130700 77726
rect 130764 77382 130792 77726
rect 130898 77744 130930 77752
rect 131040 77744 131114 77772
rect 131212 77784 131264 77790
rect 130842 77687 130898 77696
rect 130844 77648 130896 77654
rect 130844 77590 130896 77596
rect 130936 77648 130988 77654
rect 130936 77590 130988 77596
rect 130752 77376 130804 77382
rect 130752 77318 130804 77324
rect 130752 76356 130804 76362
rect 130752 76298 130804 76304
rect 130660 75336 130712 75342
rect 130660 75278 130712 75284
rect 130764 72690 130792 76298
rect 130752 72684 130804 72690
rect 130752 72626 130804 72632
rect 130856 71194 130884 77590
rect 130948 76770 130976 77590
rect 130936 76764 130988 76770
rect 130936 76706 130988 76712
rect 131040 74458 131068 77744
rect 131362 77772 131390 78132
rect 131454 77926 131482 78132
rect 131546 77926 131574 78132
rect 131442 77920 131494 77926
rect 131442 77862 131494 77868
rect 131534 77920 131586 77926
rect 131534 77862 131586 77868
rect 131638 77772 131666 78132
rect 131730 77897 131758 78132
rect 131822 77926 131850 78132
rect 131914 77926 131942 78132
rect 131810 77920 131862 77926
rect 131716 77888 131772 77897
rect 131810 77862 131862 77868
rect 131902 77920 131954 77926
rect 132006 77897 132034 78132
rect 131902 77862 131954 77868
rect 131992 77888 132048 77897
rect 131716 77823 131772 77832
rect 131992 77823 132048 77832
rect 131212 77726 131264 77732
rect 131316 77744 131390 77772
rect 131500 77744 131666 77772
rect 131946 77752 132002 77761
rect 131120 77648 131172 77654
rect 131120 77590 131172 77596
rect 131132 74905 131160 77590
rect 131118 74896 131174 74905
rect 131118 74831 131174 74840
rect 131224 74769 131252 77726
rect 131210 74760 131266 74769
rect 131210 74695 131266 74704
rect 131316 74633 131344 77744
rect 131394 77480 131450 77489
rect 131394 77415 131450 77424
rect 131302 74624 131358 74633
rect 131212 74588 131264 74594
rect 131302 74559 131358 74568
rect 131212 74530 131264 74536
rect 131028 74452 131080 74458
rect 131028 74394 131080 74400
rect 131120 74452 131172 74458
rect 131120 74394 131172 74400
rect 131132 73574 131160 74394
rect 131120 73568 131172 73574
rect 131120 73510 131172 73516
rect 131224 71262 131252 74530
rect 131408 74202 131436 77415
rect 131500 74934 131528 77744
rect 131946 77687 132002 77696
rect 131580 77648 131632 77654
rect 131580 77590 131632 77596
rect 131488 74928 131540 74934
rect 131488 74870 131540 74876
rect 131316 74174 131436 74202
rect 131212 71256 131264 71262
rect 131212 71198 131264 71204
rect 130844 71188 130896 71194
rect 130844 71130 130896 71136
rect 130580 16546 130700 16574
rect 130672 3670 130700 16546
rect 131316 3738 131344 74174
rect 131396 74112 131448 74118
rect 131396 74054 131448 74060
rect 131408 5302 131436 74054
rect 131488 74044 131540 74050
rect 131488 73986 131540 73992
rect 131500 7886 131528 73986
rect 131488 7880 131540 7886
rect 131488 7822 131540 7828
rect 131592 7750 131620 77590
rect 131672 77580 131724 77586
rect 131672 77522 131724 77528
rect 131684 7818 131712 77522
rect 131764 77512 131816 77518
rect 131764 77454 131816 77460
rect 131776 10606 131804 77454
rect 131856 77444 131908 77450
rect 131856 77386 131908 77392
rect 131868 74594 131896 77386
rect 131856 74588 131908 74594
rect 131856 74530 131908 74536
rect 131856 74248 131908 74254
rect 131856 74190 131908 74196
rect 131764 10600 131816 10606
rect 131764 10542 131816 10548
rect 131672 7812 131724 7818
rect 131672 7754 131724 7760
rect 131580 7744 131632 7750
rect 131580 7686 131632 7692
rect 131396 5296 131448 5302
rect 131396 5238 131448 5244
rect 131868 3874 131896 74190
rect 131960 74186 131988 77687
rect 132098 77636 132126 78132
rect 132190 77926 132218 78132
rect 132282 77926 132310 78132
rect 132178 77920 132230 77926
rect 132178 77862 132230 77868
rect 132270 77920 132322 77926
rect 132374 77897 132402 78132
rect 132466 77926 132494 78132
rect 132454 77920 132506 77926
rect 132270 77862 132322 77868
rect 132360 77888 132416 77897
rect 132558 77897 132586 78132
rect 132650 77926 132678 78132
rect 132742 77926 132770 78132
rect 132638 77920 132690 77926
rect 132454 77862 132506 77868
rect 132544 77888 132600 77897
rect 132360 77823 132416 77832
rect 132638 77862 132690 77868
rect 132730 77920 132782 77926
rect 132730 77862 132782 77868
rect 132544 77823 132600 77832
rect 132834 77790 132862 78132
rect 132926 77897 132954 78132
rect 132912 77888 132968 77897
rect 132912 77823 132968 77832
rect 132592 77784 132644 77790
rect 132592 77726 132644 77732
rect 132822 77784 132874 77790
rect 133018 77738 133046 78132
rect 133110 77926 133138 78132
rect 133098 77920 133150 77926
rect 133202 77897 133230 78132
rect 133098 77862 133150 77868
rect 133188 77888 133244 77897
rect 133188 77823 133244 77832
rect 133294 77772 133322 78132
rect 133386 77926 133414 78132
rect 133478 77926 133506 78132
rect 133570 77926 133598 78132
rect 133374 77920 133426 77926
rect 133374 77862 133426 77868
rect 133466 77920 133518 77926
rect 133466 77862 133518 77868
rect 133558 77920 133610 77926
rect 133662 77897 133690 78132
rect 133754 77926 133782 78132
rect 133742 77920 133794 77926
rect 133558 77862 133610 77868
rect 133648 77888 133704 77897
rect 133846 77897 133874 78132
rect 133938 77926 133966 78132
rect 134030 77926 134058 78132
rect 134122 77926 134150 78132
rect 134214 77926 134242 78132
rect 133926 77920 133978 77926
rect 133742 77862 133794 77868
rect 133832 77888 133888 77897
rect 133648 77823 133704 77832
rect 133926 77862 133978 77868
rect 134018 77920 134070 77926
rect 134018 77862 134070 77868
rect 134110 77920 134162 77926
rect 134110 77862 134162 77868
rect 134202 77920 134254 77926
rect 134202 77862 134254 77868
rect 133832 77823 133888 77832
rect 133880 77784 133932 77790
rect 133294 77744 133368 77772
rect 132822 77726 132874 77732
rect 132316 77716 132368 77722
rect 132316 77658 132368 77664
rect 132224 77648 132276 77654
rect 132098 77608 132172 77636
rect 132038 77480 132094 77489
rect 132038 77415 132094 77424
rect 131948 74180 132000 74186
rect 131948 74122 132000 74128
rect 131856 3868 131908 3874
rect 131856 3810 131908 3816
rect 131764 3800 131816 3806
rect 131764 3742 131816 3748
rect 131304 3732 131356 3738
rect 131304 3674 131356 3680
rect 130660 3664 130712 3670
rect 130660 3606 130712 3612
rect 130384 3596 130436 3602
rect 130384 3538 130436 3544
rect 129844 3454 130608 3482
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128464 462 128952 490
rect 130580 480 130608 3454
rect 131776 480 131804 3742
rect 132052 3738 132080 77415
rect 132144 74050 132172 77608
rect 132224 77590 132276 77596
rect 132236 74254 132264 77590
rect 132328 74866 132356 77658
rect 132408 77580 132460 77586
rect 132408 77522 132460 77528
rect 132316 74860 132368 74866
rect 132316 74802 132368 74808
rect 132224 74248 132276 74254
rect 132224 74190 132276 74196
rect 132420 74118 132448 77522
rect 132498 77208 132554 77217
rect 132604 77194 132632 77726
rect 132972 77710 133046 77738
rect 132684 77648 132736 77654
rect 132684 77590 132736 77596
rect 132696 77294 132724 77590
rect 132696 77266 132816 77294
rect 132604 77166 132724 77194
rect 132498 77143 132554 77152
rect 132408 74112 132460 74118
rect 132408 74054 132460 74060
rect 132132 74044 132184 74050
rect 132132 73986 132184 73992
rect 132512 71233 132540 77143
rect 132590 76392 132646 76401
rect 132590 76327 132646 76336
rect 132604 74225 132632 76327
rect 132696 75041 132724 77166
rect 132682 75032 132738 75041
rect 132682 74967 132738 74976
rect 132788 74497 132816 77266
rect 132866 76256 132922 76265
rect 132866 76191 132922 76200
rect 132774 74488 132830 74497
rect 132774 74423 132830 74432
rect 132776 74248 132828 74254
rect 132590 74216 132646 74225
rect 132776 74190 132828 74196
rect 132590 74151 132646 74160
rect 132684 74112 132736 74118
rect 132684 74054 132736 74060
rect 132592 73228 132644 73234
rect 132592 73170 132644 73176
rect 132604 71330 132632 73170
rect 132592 71324 132644 71330
rect 132592 71266 132644 71272
rect 132498 71224 132554 71233
rect 132498 71159 132554 71168
rect 132696 8022 132724 74054
rect 132788 8090 132816 74190
rect 132776 8084 132828 8090
rect 132776 8026 132828 8032
rect 132684 8016 132736 8022
rect 132684 7958 132736 7964
rect 132880 7954 132908 76191
rect 132972 75070 133000 77710
rect 133236 77648 133288 77654
rect 133236 77590 133288 77596
rect 133052 77580 133104 77586
rect 133052 77522 133104 77528
rect 133144 77580 133196 77586
rect 133144 77522 133196 77528
rect 132960 75064 133012 75070
rect 132960 75006 133012 75012
rect 133064 74474 133092 77522
rect 132972 74446 133092 74474
rect 132972 73234 133000 74446
rect 133052 74316 133104 74322
rect 133052 74258 133104 74264
rect 132960 73228 133012 73234
rect 132960 73170 133012 73176
rect 132960 73024 133012 73030
rect 132960 72966 133012 72972
rect 132972 10674 133000 72966
rect 133064 20058 133092 74258
rect 133052 20052 133104 20058
rect 133052 19994 133104 20000
rect 132960 10668 133012 10674
rect 132960 10610 133012 10616
rect 132868 7948 132920 7954
rect 132868 7890 132920 7896
rect 133156 5438 133184 77522
rect 133248 70394 133276 77590
rect 133340 73030 133368 77744
rect 133510 77752 133566 77761
rect 133510 77687 133566 77696
rect 133786 77752 133842 77761
rect 134306 77772 134334 78132
rect 134398 77897 134426 78132
rect 134490 77926 134518 78132
rect 134582 77926 134610 78132
rect 134478 77920 134530 77926
rect 134384 77888 134440 77897
rect 134478 77862 134530 77868
rect 134570 77920 134622 77926
rect 134570 77862 134622 77868
rect 134384 77823 134440 77832
rect 133880 77726 133932 77732
rect 134260 77744 134334 77772
rect 134432 77784 134484 77790
rect 133786 77687 133842 77696
rect 133524 77568 133552 77687
rect 133696 77580 133748 77586
rect 133524 77540 133644 77568
rect 133420 77512 133472 77518
rect 133420 77454 133472 77460
rect 133432 74186 133460 77454
rect 133512 77444 133564 77450
rect 133512 77386 133564 77392
rect 133524 75818 133552 77386
rect 133512 75812 133564 75818
rect 133512 75754 133564 75760
rect 133512 75064 133564 75070
rect 133512 75006 133564 75012
rect 133420 74180 133472 74186
rect 133420 74122 133472 74128
rect 133524 73166 133552 75006
rect 133616 74118 133644 77540
rect 133696 77522 133748 77528
rect 133708 74254 133736 77522
rect 133800 74322 133828 77687
rect 133892 75138 133920 77726
rect 134064 77648 134116 77654
rect 134064 77590 134116 77596
rect 133972 77512 134024 77518
rect 133972 77454 134024 77460
rect 133984 75410 134012 77454
rect 133972 75404 134024 75410
rect 133972 75346 134024 75352
rect 133880 75132 133932 75138
rect 133880 75074 133932 75080
rect 133972 75132 134024 75138
rect 133972 75074 134024 75080
rect 133984 74984 134012 75074
rect 134076 75041 134104 77590
rect 134154 77344 134210 77353
rect 134154 77279 134156 77288
rect 134208 77279 134210 77288
rect 134156 77250 134208 77256
rect 134260 76208 134288 77744
rect 134674 77772 134702 78132
rect 134766 77897 134794 78132
rect 134858 77926 134886 78132
rect 134950 77926 134978 78132
rect 135042 77926 135070 78132
rect 134846 77920 134898 77926
rect 134752 77888 134808 77897
rect 134846 77862 134898 77868
rect 134938 77920 134990 77926
rect 134938 77862 134990 77868
rect 135030 77920 135082 77926
rect 135030 77862 135082 77868
rect 134752 77823 134808 77832
rect 134432 77726 134484 77732
rect 134522 77752 134578 77761
rect 134340 77580 134392 77586
rect 134340 77522 134392 77528
rect 134352 76401 134380 77522
rect 134338 76392 134394 76401
rect 134338 76327 134394 76336
rect 134168 76180 134288 76208
rect 133892 74956 134012 74984
rect 134062 75032 134118 75041
rect 134062 74967 134118 74976
rect 133788 74316 133840 74322
rect 133788 74258 133840 74264
rect 133696 74248 133748 74254
rect 133696 74190 133748 74196
rect 133604 74112 133656 74118
rect 133604 74054 133656 74060
rect 133512 73160 133564 73166
rect 133512 73102 133564 73108
rect 133328 73024 133380 73030
rect 133328 72966 133380 72972
rect 133248 70366 133368 70394
rect 133144 5432 133196 5438
rect 133144 5374 133196 5380
rect 133340 5370 133368 70366
rect 133328 5364 133380 5370
rect 133328 5306 133380 5312
rect 132040 3732 132092 3738
rect 132040 3674 132092 3680
rect 132960 3664 133012 3670
rect 132960 3606 133012 3612
rect 132972 480 133000 3606
rect 128924 354 128952 462
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133892 354 133920 74956
rect 134064 74860 134116 74866
rect 134064 74802 134116 74808
rect 133972 74248 134024 74254
rect 133972 74190 134024 74196
rect 133984 69698 134012 74190
rect 134076 71398 134104 74802
rect 134168 74361 134196 76180
rect 134154 74352 134210 74361
rect 134154 74287 134210 74296
rect 134444 74254 134472 77726
rect 134522 77687 134578 77696
rect 134628 77744 134702 77772
rect 135134 77772 135162 78132
rect 135226 77926 135254 78132
rect 135318 77926 135346 78132
rect 135214 77920 135266 77926
rect 135214 77862 135266 77868
rect 135306 77920 135358 77926
rect 135306 77862 135358 77868
rect 135410 77795 135438 78132
rect 135502 77926 135530 78132
rect 135594 77926 135622 78132
rect 135686 77926 135714 78132
rect 135490 77920 135542 77926
rect 135490 77862 135542 77868
rect 135582 77920 135634 77926
rect 135582 77862 135634 77868
rect 135674 77920 135726 77926
rect 135674 77862 135726 77868
rect 135396 77786 135452 77795
rect 135134 77744 135208 77772
rect 134536 74866 134564 77687
rect 134524 74860 134576 74866
rect 134524 74802 134576 74808
rect 134628 74338 134656 77744
rect 134800 77716 134852 77722
rect 134800 77658 134852 77664
rect 134892 77716 134944 77722
rect 134892 77658 134944 77664
rect 134984 77716 135036 77722
rect 134984 77658 135036 77664
rect 134708 77580 134760 77586
rect 134708 77522 134760 77528
rect 134536 74310 134656 74338
rect 134432 74248 134484 74254
rect 134432 74190 134484 74196
rect 134536 74100 134564 74310
rect 134616 74248 134668 74254
rect 134616 74190 134668 74196
rect 134168 74072 134564 74100
rect 134064 71392 134116 71398
rect 134064 71334 134116 71340
rect 133972 69692 134024 69698
rect 133972 69634 134024 69640
rect 134168 11762 134196 74072
rect 134524 73976 134576 73982
rect 134524 73918 134576 73924
rect 134156 11756 134208 11762
rect 134156 11698 134208 11704
rect 134536 4146 134564 73918
rect 134524 4140 134576 4146
rect 134524 4082 134576 4088
rect 134628 3534 134656 74190
rect 134720 9314 134748 77522
rect 134812 74662 134840 77658
rect 134904 75002 134932 77658
rect 134892 74996 134944 75002
rect 134892 74938 134944 74944
rect 134800 74656 134852 74662
rect 134800 74598 134852 74604
rect 134996 72894 135024 77658
rect 135180 76616 135208 77744
rect 135778 77772 135806 78132
rect 135870 77926 135898 78132
rect 135962 77926 135990 78132
rect 135858 77920 135910 77926
rect 135858 77862 135910 77868
rect 135950 77920 136002 77926
rect 136054 77897 136082 78132
rect 135950 77862 136002 77868
rect 136040 77888 136096 77897
rect 136146 77858 136174 78132
rect 136238 77897 136266 78132
rect 136224 77888 136280 77897
rect 136040 77823 136096 77832
rect 136134 77852 136186 77858
rect 136224 77823 136280 77832
rect 136134 77794 136186 77800
rect 136330 77772 136358 78132
rect 136422 77897 136450 78132
rect 136514 77926 136542 78132
rect 136502 77920 136554 77926
rect 136408 77888 136464 77897
rect 136502 77862 136554 77868
rect 136606 77858 136634 78132
rect 136698 77897 136726 78132
rect 136790 77926 136818 78132
rect 136778 77920 136830 77926
rect 136684 77888 136740 77897
rect 136408 77823 136464 77832
rect 136594 77852 136646 77858
rect 136882 77897 136910 78132
rect 136778 77862 136830 77868
rect 136868 77888 136924 77897
rect 136684 77823 136740 77832
rect 136868 77823 136924 77832
rect 136594 77794 136646 77800
rect 135778 77744 135852 77772
rect 135260 77716 135312 77722
rect 135396 77721 135452 77730
rect 135260 77658 135312 77664
rect 135628 77716 135680 77722
rect 135628 77658 135680 77664
rect 135088 76588 135208 76616
rect 135088 75206 135116 76588
rect 135076 75200 135128 75206
rect 135076 75142 135128 75148
rect 135076 74996 135128 75002
rect 135076 74938 135128 74944
rect 134984 72888 135036 72894
rect 134984 72830 135036 72836
rect 135088 70394 135116 74938
rect 135272 74848 135300 77658
rect 135352 77648 135404 77654
rect 135352 77590 135404 77596
rect 135444 77648 135496 77654
rect 135444 77590 135496 77596
rect 135180 74820 135300 74848
rect 135180 74254 135208 74820
rect 135260 74724 135312 74730
rect 135260 74666 135312 74672
rect 135168 74248 135220 74254
rect 135168 74190 135220 74196
rect 135272 70394 135300 74666
rect 135364 73982 135392 77590
rect 135456 75041 135484 77590
rect 135536 77512 135588 77518
rect 135536 77454 135588 77460
rect 135548 75070 135576 77454
rect 135536 75064 135588 75070
rect 135442 75032 135498 75041
rect 135536 75006 135588 75012
rect 135442 74967 135498 74976
rect 135536 74928 135588 74934
rect 135536 74870 135588 74876
rect 135444 74860 135496 74866
rect 135444 74802 135496 74808
rect 135352 73976 135404 73982
rect 135352 73918 135404 73924
rect 135088 70366 135208 70394
rect 135272 70366 135392 70394
rect 134708 9308 134760 9314
rect 134708 9250 134760 9256
rect 135180 3534 135208 70366
rect 135364 3602 135392 70366
rect 135456 3738 135484 74802
rect 135444 3732 135496 3738
rect 135444 3674 135496 3680
rect 135548 3670 135576 74870
rect 135640 74798 135668 77658
rect 135720 75064 135772 75070
rect 135720 75006 135772 75012
rect 135628 74792 135680 74798
rect 135628 74734 135680 74740
rect 135628 74656 135680 74662
rect 135628 74598 135680 74604
rect 135640 3670 135668 74598
rect 135732 3874 135760 75006
rect 135720 3868 135772 3874
rect 135720 3810 135772 3816
rect 135824 3806 135852 77744
rect 136178 77752 136234 77761
rect 136088 77716 136140 77722
rect 136330 77744 136404 77772
rect 136178 77687 136234 77696
rect 136088 77658 136140 77664
rect 135904 77648 135956 77654
rect 135904 77590 135956 77596
rect 135916 74934 135944 77590
rect 135996 77580 136048 77586
rect 135996 77522 136048 77528
rect 135904 74928 135956 74934
rect 135904 74870 135956 74876
rect 135904 74792 135956 74798
rect 135904 74734 135956 74740
rect 135916 16574 135944 74734
rect 136008 20670 136036 77522
rect 136100 75138 136128 77658
rect 136088 75132 136140 75138
rect 136088 75074 136140 75080
rect 136086 75032 136142 75041
rect 136086 74967 136142 74976
rect 135996 20664 136048 20670
rect 135996 20606 136048 20612
rect 135916 16546 136036 16574
rect 136008 4214 136036 16546
rect 135996 4208 136048 4214
rect 135996 4150 136048 4156
rect 135812 3800 135864 3806
rect 135812 3742 135864 3748
rect 135536 3664 135588 3670
rect 135536 3606 135588 3612
rect 135628 3664 135680 3670
rect 135628 3606 135680 3612
rect 135352 3596 135404 3602
rect 135352 3538 135404 3544
rect 134616 3528 134668 3534
rect 134616 3470 134668 3476
rect 135168 3528 135220 3534
rect 136100 3482 136128 74967
rect 136192 74866 136220 77687
rect 136272 77648 136324 77654
rect 136272 77590 136324 77596
rect 136180 74860 136232 74866
rect 136180 74802 136232 74808
rect 136284 74730 136312 77590
rect 136272 74724 136324 74730
rect 136272 74666 136324 74672
rect 136376 74662 136404 77744
rect 136822 77752 136878 77761
rect 136732 77716 136784 77722
rect 136822 77687 136878 77696
rect 136974 77704 137002 78132
rect 137066 77858 137094 78132
rect 137054 77852 137106 77858
rect 137054 77794 137106 77800
rect 136732 77658 136784 77664
rect 136640 77648 136692 77654
rect 136640 77590 136692 77596
rect 136548 77580 136600 77586
rect 136468 77540 136548 77568
rect 136468 74798 136496 77540
rect 136548 77522 136600 77528
rect 136546 77480 136602 77489
rect 136546 77415 136602 77424
rect 136560 75070 136588 77415
rect 136548 75064 136600 75070
rect 136548 75006 136600 75012
rect 136652 74866 136680 77590
rect 136744 75002 136772 77658
rect 136732 74996 136784 75002
rect 136732 74938 136784 74944
rect 136640 74860 136692 74866
rect 136640 74802 136692 74808
rect 136456 74792 136508 74798
rect 136456 74734 136508 74740
rect 136364 74656 136416 74662
rect 136364 74598 136416 74604
rect 136836 74066 136864 77687
rect 136974 77676 137048 77704
rect 136916 77580 136968 77586
rect 136916 77522 136968 77528
rect 136744 74038 136864 74066
rect 136744 73710 136772 74038
rect 136824 73976 136876 73982
rect 136824 73918 136876 73924
rect 136732 73704 136784 73710
rect 136732 73646 136784 73652
rect 136732 73500 136784 73506
rect 136732 73442 136784 73448
rect 136744 5370 136772 73442
rect 136732 5364 136784 5370
rect 136732 5306 136784 5312
rect 136836 4758 136864 73918
rect 136928 5166 136956 77522
rect 137020 75070 137048 77676
rect 137158 77636 137186 78132
rect 137250 77738 137278 78132
rect 137342 77926 137370 78132
rect 137330 77920 137382 77926
rect 137434 77897 137462 78132
rect 137526 77926 137554 78132
rect 137618 77926 137646 78132
rect 137514 77920 137566 77926
rect 137330 77862 137382 77868
rect 137420 77888 137476 77897
rect 137514 77862 137566 77868
rect 137606 77920 137658 77926
rect 137606 77862 137658 77868
rect 137420 77823 137476 77832
rect 137374 77752 137430 77761
rect 137250 77710 137324 77738
rect 137158 77608 137232 77636
rect 137008 75064 137060 75070
rect 137008 75006 137060 75012
rect 137008 74860 137060 74866
rect 137008 74802 137060 74808
rect 136916 5160 136968 5166
rect 136916 5102 136968 5108
rect 137020 5098 137048 74802
rect 137100 74316 137152 74322
rect 137100 74258 137152 74264
rect 137008 5092 137060 5098
rect 137008 5034 137060 5040
rect 137112 4962 137140 74258
rect 137204 57934 137232 77608
rect 137296 73506 137324 77710
rect 137374 77687 137430 77696
rect 137468 77716 137520 77722
rect 137284 73500 137336 73506
rect 137284 73442 137336 73448
rect 137282 73400 137338 73409
rect 137282 73335 137338 73344
rect 137296 62150 137324 73335
rect 137388 73302 137416 77687
rect 137710 77704 137738 78132
rect 137802 77926 137830 78132
rect 137894 77926 137922 78132
rect 137986 77926 138014 78132
rect 137790 77920 137842 77926
rect 137790 77862 137842 77868
rect 137882 77920 137934 77926
rect 137882 77862 137934 77868
rect 137974 77920 138026 77926
rect 137974 77862 138026 77868
rect 137836 77784 137888 77790
rect 138078 77772 138106 78132
rect 138170 77926 138198 78132
rect 138262 77926 138290 78132
rect 138354 77926 138382 78132
rect 138158 77920 138210 77926
rect 138158 77862 138210 77868
rect 138250 77920 138302 77926
rect 138250 77862 138302 77868
rect 138342 77920 138394 77926
rect 138342 77862 138394 77868
rect 137836 77726 137888 77732
rect 138032 77744 138106 77772
rect 138296 77784 138348 77790
rect 137710 77676 137784 77704
rect 137468 77658 137520 77664
rect 137480 74322 137508 77658
rect 137652 77580 137704 77586
rect 137652 77522 137704 77528
rect 137468 74316 137520 74322
rect 137468 74258 137520 74264
rect 137376 73296 137428 73302
rect 137376 73238 137428 73244
rect 137664 71670 137692 77522
rect 137756 75206 137784 77676
rect 137744 75200 137796 75206
rect 137744 75142 137796 75148
rect 137744 74996 137796 75002
rect 137744 74938 137796 74944
rect 137652 71664 137704 71670
rect 137652 71606 137704 71612
rect 137284 62144 137336 62150
rect 137284 62086 137336 62092
rect 137192 57928 137244 57934
rect 137192 57870 137244 57876
rect 137100 4956 137152 4962
rect 137100 4898 137152 4904
rect 136824 4752 136876 4758
rect 136824 4694 136876 4700
rect 137756 4146 137784 74938
rect 137848 73982 137876 77726
rect 137928 77716 137980 77722
rect 137928 77658 137980 77664
rect 137940 75041 137968 77658
rect 137926 75032 137982 75041
rect 137926 74967 137982 74976
rect 137836 73976 137888 73982
rect 137836 73918 137888 73924
rect 138032 73817 138060 77744
rect 138296 77726 138348 77732
rect 138204 77716 138256 77722
rect 138204 77658 138256 77664
rect 138112 77580 138164 77586
rect 138112 77522 138164 77528
rect 138124 77489 138152 77522
rect 138110 77480 138166 77489
rect 138110 77415 138166 77424
rect 138112 74928 138164 74934
rect 138112 74870 138164 74876
rect 138018 73808 138074 73817
rect 138018 73743 138074 73752
rect 138124 5030 138152 74870
rect 138112 5024 138164 5030
rect 138112 4966 138164 4972
rect 138216 4826 138244 77658
rect 138308 74118 138336 77726
rect 138446 77636 138474 78132
rect 138538 77926 138566 78132
rect 138630 77926 138658 78132
rect 138526 77920 138578 77926
rect 138526 77862 138578 77868
rect 138618 77920 138670 77926
rect 138618 77862 138670 77868
rect 138722 77738 138750 78132
rect 138814 77926 138842 78132
rect 138802 77920 138854 77926
rect 138802 77862 138854 77868
rect 138906 77772 138934 78132
rect 138998 77926 139026 78132
rect 138986 77920 139038 77926
rect 138986 77862 139038 77868
rect 138860 77761 138934 77772
rect 138676 77710 138750 77738
rect 138846 77752 138934 77761
rect 138446 77608 138520 77636
rect 138386 77480 138442 77489
rect 138386 77415 138442 77424
rect 138296 74112 138348 74118
rect 138296 74054 138348 74060
rect 138294 73944 138350 73953
rect 138294 73879 138350 73888
rect 138308 5302 138336 73879
rect 138400 9246 138428 77415
rect 138492 62218 138520 77608
rect 138676 77568 138704 77710
rect 138902 77744 138934 77752
rect 139090 77772 139118 78132
rect 139182 77926 139210 78132
rect 139170 77920 139222 77926
rect 139170 77862 139222 77868
rect 139274 77772 139302 78132
rect 139366 77926 139394 78132
rect 139458 77926 139486 78132
rect 139550 77926 139578 78132
rect 139642 77926 139670 78132
rect 139734 77926 139762 78132
rect 139354 77920 139406 77926
rect 139354 77862 139406 77868
rect 139446 77920 139498 77926
rect 139446 77862 139498 77868
rect 139538 77920 139590 77926
rect 139538 77862 139590 77868
rect 139630 77920 139682 77926
rect 139630 77862 139682 77868
rect 139722 77920 139774 77926
rect 139722 77862 139774 77868
rect 139826 77772 139854 78132
rect 139090 77744 139164 77772
rect 138846 77687 138902 77696
rect 138848 77648 138900 77654
rect 138848 77590 138900 77596
rect 138940 77648 138992 77654
rect 138940 77590 138992 77596
rect 138584 77540 138704 77568
rect 138756 77580 138808 77586
rect 138584 77489 138612 77540
rect 138756 77522 138808 77528
rect 138570 77480 138626 77489
rect 138570 77415 138626 77424
rect 138664 77444 138716 77450
rect 138664 77386 138716 77392
rect 138572 77376 138624 77382
rect 138570 77344 138572 77353
rect 138624 77344 138626 77353
rect 138570 77279 138626 77288
rect 138572 77240 138624 77246
rect 138572 77182 138624 77188
rect 138584 74202 138612 77182
rect 138676 75002 138704 77386
rect 138664 74996 138716 75002
rect 138664 74938 138716 74944
rect 138768 74934 138796 77522
rect 138756 74928 138808 74934
rect 138756 74870 138808 74876
rect 138584 74174 138796 74202
rect 138664 74112 138716 74118
rect 138664 74054 138716 74060
rect 138572 74044 138624 74050
rect 138572 73986 138624 73992
rect 138584 69018 138612 73986
rect 138676 69698 138704 74054
rect 138768 72486 138796 74174
rect 138860 74050 138888 77590
rect 138952 75041 138980 77590
rect 139032 77512 139084 77518
rect 139032 77454 139084 77460
rect 139044 76401 139072 77454
rect 139030 76392 139086 76401
rect 139030 76327 139086 76336
rect 138938 75032 138994 75041
rect 138938 74967 138994 74976
rect 139032 74996 139084 75002
rect 139032 74938 139084 74944
rect 138848 74044 138900 74050
rect 138848 73986 138900 73992
rect 138940 73704 138992 73710
rect 138940 73646 138992 73652
rect 138756 72480 138808 72486
rect 138756 72422 138808 72428
rect 138664 69692 138716 69698
rect 138664 69634 138716 69640
rect 138572 69012 138624 69018
rect 138572 68954 138624 68960
rect 138480 62212 138532 62218
rect 138480 62154 138532 62160
rect 138664 62144 138716 62150
rect 138664 62086 138716 62092
rect 138388 9240 138440 9246
rect 138388 9182 138440 9188
rect 138296 5296 138348 5302
rect 138296 5238 138348 5244
rect 138204 4820 138256 4826
rect 138204 4762 138256 4768
rect 137744 4140 137796 4146
rect 137744 4082 137796 4088
rect 138676 4010 138704 62086
rect 138952 4078 138980 73646
rect 138940 4072 138992 4078
rect 138940 4014 138992 4020
rect 138664 4004 138716 4010
rect 138664 3946 138716 3952
rect 137652 3732 137704 3738
rect 137652 3674 137704 3680
rect 136456 3596 136508 3602
rect 136456 3538 136508 3544
rect 135168 3470 135220 3476
rect 135272 3454 136128 3482
rect 135272 480 135300 3454
rect 136468 480 136496 3538
rect 137664 480 137692 3674
rect 138848 3664 138900 3670
rect 138848 3606 138900 3612
rect 138860 480 138888 3606
rect 139044 3466 139072 74938
rect 139136 73001 139164 77744
rect 139228 77744 139302 77772
rect 139780 77744 139854 77772
rect 139918 77761 139946 78132
rect 139904 77752 139960 77761
rect 139228 75274 139256 77744
rect 139780 77738 139808 77744
rect 139492 77716 139544 77722
rect 139492 77658 139544 77664
rect 139642 77710 139808 77738
rect 139308 77648 139360 77654
rect 139308 77590 139360 77596
rect 139400 77648 139452 77654
rect 139400 77590 139452 77596
rect 139320 76401 139348 77590
rect 139306 76392 139362 76401
rect 139306 76327 139362 76336
rect 139412 75750 139440 77590
rect 139400 75744 139452 75750
rect 139400 75686 139452 75692
rect 139216 75268 139268 75274
rect 139216 75210 139268 75216
rect 139400 74044 139452 74050
rect 139400 73986 139452 73992
rect 139122 72992 139178 73001
rect 139122 72927 139178 72936
rect 139412 24546 139440 73986
rect 139504 25974 139532 77658
rect 139642 77636 139670 77710
rect 139904 77687 139960 77696
rect 140010 77704 140038 78132
rect 140102 77772 140130 78132
rect 140194 77926 140222 78132
rect 140182 77920 140234 77926
rect 140182 77862 140234 77868
rect 140286 77772 140314 78132
rect 140378 77926 140406 78132
rect 140366 77920 140418 77926
rect 140366 77862 140418 77868
rect 140102 77744 140176 77772
rect 140286 77744 140360 77772
rect 140010 77676 140084 77704
rect 139642 77608 139716 77636
rect 139584 77376 139636 77382
rect 139584 77318 139636 77324
rect 139596 77217 139624 77318
rect 139582 77208 139638 77217
rect 139582 77143 139638 77152
rect 139584 73500 139636 73506
rect 139584 73442 139636 73448
rect 139492 25968 139544 25974
rect 139492 25910 139544 25916
rect 139596 25838 139624 73442
rect 139688 25906 139716 77608
rect 139952 77580 140004 77586
rect 139952 77522 140004 77528
rect 139768 77512 139820 77518
rect 139768 77454 139820 77460
rect 139860 77512 139912 77518
rect 139860 77454 139912 77460
rect 139780 46238 139808 77454
rect 139872 75041 139900 77454
rect 139858 75032 139914 75041
rect 139858 74967 139914 74976
rect 139860 74928 139912 74934
rect 139860 74870 139912 74876
rect 139872 63170 139900 74870
rect 139964 74304 139992 77522
rect 140056 74934 140084 77676
rect 140044 74928 140096 74934
rect 140044 74870 140096 74876
rect 139964 74276 140084 74304
rect 139952 74180 140004 74186
rect 139952 74122 140004 74128
rect 139964 64598 139992 74122
rect 140056 67250 140084 74276
rect 140148 73506 140176 77744
rect 140228 77648 140280 77654
rect 140228 77590 140280 77596
rect 140240 74050 140268 77590
rect 140332 74186 140360 77744
rect 140470 77738 140498 78132
rect 140562 77858 140590 78132
rect 140550 77852 140602 77858
rect 140550 77794 140602 77800
rect 140654 77738 140682 78132
rect 140746 77926 140774 78132
rect 140838 77926 140866 78132
rect 140734 77920 140786 77926
rect 140734 77862 140786 77868
rect 140826 77920 140878 77926
rect 140826 77862 140878 77868
rect 140470 77710 140544 77738
rect 140412 77648 140464 77654
rect 140516 77625 140544 77710
rect 140608 77710 140682 77738
rect 140780 77716 140832 77722
rect 140412 77590 140464 77596
rect 140502 77616 140558 77625
rect 140424 75410 140452 77590
rect 140502 77551 140558 77560
rect 140502 77480 140558 77489
rect 140502 77415 140558 77424
rect 140412 75404 140464 75410
rect 140412 75346 140464 75352
rect 140412 75268 140464 75274
rect 140412 75210 140464 75216
rect 140320 74180 140372 74186
rect 140320 74122 140372 74128
rect 140228 74044 140280 74050
rect 140228 73986 140280 73992
rect 140136 73500 140188 73506
rect 140136 73442 140188 73448
rect 140044 67244 140096 67250
rect 140044 67186 140096 67192
rect 139952 64592 140004 64598
rect 139952 64534 140004 64540
rect 139860 63164 139912 63170
rect 139860 63106 139912 63112
rect 140044 62212 140096 62218
rect 140044 62154 140096 62160
rect 139768 46232 139820 46238
rect 139768 46174 139820 46180
rect 139676 25900 139728 25906
rect 139676 25842 139728 25848
rect 139584 25832 139636 25838
rect 139584 25774 139636 25780
rect 139400 24540 139452 24546
rect 139400 24482 139452 24488
rect 140056 12434 140084 62154
rect 140136 57928 140188 57934
rect 140136 57870 140188 57876
rect 139964 12406 140084 12434
rect 139964 3670 139992 12406
rect 140148 3874 140176 57870
rect 140424 26042 140452 75210
rect 140516 71774 140544 77415
rect 140608 75041 140636 77710
rect 140780 77658 140832 77664
rect 140688 77648 140740 77654
rect 140688 77590 140740 77596
rect 140594 75032 140650 75041
rect 140594 74967 140650 74976
rect 140700 74905 140728 77590
rect 140792 74984 140820 77658
rect 140930 77568 140958 78132
rect 141022 77926 141050 78132
rect 141114 77926 141142 78132
rect 141206 77926 141234 78132
rect 141298 77926 141326 78132
rect 141010 77920 141062 77926
rect 141010 77862 141062 77868
rect 141102 77920 141154 77926
rect 141102 77862 141154 77868
rect 141194 77920 141246 77926
rect 141194 77862 141246 77868
rect 141286 77920 141338 77926
rect 141286 77862 141338 77868
rect 141148 77648 141200 77654
rect 140884 77540 140958 77568
rect 141068 77608 141148 77636
rect 140884 75274 140912 77540
rect 140964 77240 141016 77246
rect 140964 77182 141016 77188
rect 140872 75268 140924 75274
rect 140872 75210 140924 75216
rect 140792 74956 140912 74984
rect 140686 74896 140742 74905
rect 140686 74831 140742 74840
rect 140780 74860 140832 74866
rect 140780 74802 140832 74808
rect 140516 71746 140728 71774
rect 140700 71466 140728 71746
rect 140688 71460 140740 71466
rect 140688 71402 140740 71408
rect 140412 26036 140464 26042
rect 140412 25978 140464 25984
rect 140792 6662 140820 74802
rect 140884 74730 140912 74956
rect 140872 74724 140924 74730
rect 140872 74666 140924 74672
rect 140976 74610 141004 77182
rect 140884 74582 141004 74610
rect 140884 17678 140912 74582
rect 140964 73092 141016 73098
rect 140964 73034 141016 73040
rect 140976 27266 141004 73034
rect 141068 27334 141096 77608
rect 141390 77636 141418 78132
rect 141482 77738 141510 78132
rect 141574 77926 141602 78132
rect 141666 77926 141694 78132
rect 141562 77920 141614 77926
rect 141562 77862 141614 77868
rect 141654 77920 141706 77926
rect 141654 77862 141706 77868
rect 141608 77784 141660 77790
rect 141482 77710 141556 77738
rect 141758 77738 141786 78132
rect 141850 77926 141878 78132
rect 141942 77926 141970 78132
rect 141838 77920 141890 77926
rect 141838 77862 141890 77868
rect 141930 77920 141982 77926
rect 141930 77862 141982 77868
rect 141608 77726 141660 77732
rect 141390 77608 141464 77636
rect 141148 77590 141200 77596
rect 141332 77512 141384 77518
rect 141332 77454 141384 77460
rect 141240 77444 141292 77450
rect 141240 77386 141292 77392
rect 141148 77376 141200 77382
rect 141148 77318 141200 77324
rect 141160 75818 141188 77318
rect 141148 75812 141200 75818
rect 141148 75754 141200 75760
rect 141148 70916 141200 70922
rect 141148 70858 141200 70864
rect 141160 28762 141188 70858
rect 141252 34202 141280 77386
rect 141240 34196 141292 34202
rect 141240 34138 141292 34144
rect 141344 33862 141372 77454
rect 141436 74866 141464 77608
rect 141424 74860 141476 74866
rect 141424 74802 141476 74808
rect 141528 73098 141556 77710
rect 141516 73092 141568 73098
rect 141516 73034 141568 73040
rect 141620 71774 141648 77726
rect 141436 71746 141648 71774
rect 141712 77710 141786 77738
rect 141884 77716 141936 77722
rect 141436 64530 141464 71746
rect 141712 70922 141740 77710
rect 142034 77704 142062 78132
rect 141884 77658 141936 77664
rect 141988 77676 142062 77704
rect 141792 77648 141844 77654
rect 141792 77590 141844 77596
rect 141804 71330 141832 77590
rect 141792 71324 141844 71330
rect 141792 71266 141844 71272
rect 141700 70916 141752 70922
rect 141700 70858 141752 70864
rect 141896 70394 141924 77658
rect 141988 74225 142016 77676
rect 142126 77636 142154 78132
rect 142218 77926 142246 78132
rect 142310 77926 142338 78132
rect 142206 77920 142258 77926
rect 142206 77862 142258 77868
rect 142298 77920 142350 77926
rect 142298 77862 142350 77868
rect 142402 77772 142430 78132
rect 142494 77926 142522 78132
rect 142586 77926 142614 78132
rect 142678 77926 142706 78132
rect 142770 77926 142798 78132
rect 142482 77920 142534 77926
rect 142482 77862 142534 77868
rect 142574 77920 142626 77926
rect 142574 77862 142626 77868
rect 142666 77920 142718 77926
rect 142666 77862 142718 77868
rect 142758 77920 142810 77926
rect 142758 77862 142810 77868
rect 142356 77744 142430 77772
rect 142252 77716 142304 77722
rect 142252 77658 142304 77664
rect 142080 77608 142154 77636
rect 142080 74633 142108 77608
rect 142160 77512 142212 77518
rect 142160 77454 142212 77460
rect 142066 74624 142122 74633
rect 142066 74559 142122 74568
rect 141974 74216 142030 74225
rect 141974 74151 142030 74160
rect 141528 70366 141924 70394
rect 141528 67182 141556 70366
rect 141516 67176 141568 67182
rect 141516 67118 141568 67124
rect 141424 64524 141476 64530
rect 141424 64466 141476 64472
rect 141332 33856 141384 33862
rect 141332 33798 141384 33804
rect 141148 28756 141200 28762
rect 141148 28698 141200 28704
rect 141056 27328 141108 27334
rect 141056 27270 141108 27276
rect 140964 27260 141016 27266
rect 140964 27202 141016 27208
rect 140872 17672 140924 17678
rect 140872 17614 140924 17620
rect 140780 6656 140832 6662
rect 140780 6598 140832 6604
rect 142172 6594 142200 77454
rect 142264 76974 142292 77658
rect 142356 77586 142384 77744
rect 142862 77738 142890 78132
rect 142620 77716 142672 77722
rect 142620 77658 142672 77664
rect 142816 77710 142890 77738
rect 142954 77738 142982 78132
rect 143046 77858 143074 78132
rect 143034 77852 143086 77858
rect 143034 77794 143086 77800
rect 143138 77761 143166 78132
rect 143124 77752 143180 77761
rect 142954 77710 143028 77738
rect 142436 77648 142488 77654
rect 142436 77590 142488 77596
rect 142344 77580 142396 77586
rect 142344 77522 142396 77528
rect 142344 77444 142396 77450
rect 142344 77386 142396 77392
rect 142252 76968 142304 76974
rect 142252 76910 142304 76916
rect 142252 74248 142304 74254
rect 142252 74190 142304 74196
rect 142264 28626 142292 74190
rect 142356 74118 142384 77386
rect 142344 74112 142396 74118
rect 142344 74054 142396 74060
rect 142344 70916 142396 70922
rect 142344 70858 142396 70864
rect 142252 28620 142304 28626
rect 142252 28562 142304 28568
rect 142356 28558 142384 70858
rect 142448 28694 142476 77590
rect 142632 77466 142660 77658
rect 142712 77648 142764 77654
rect 142712 77590 142764 77596
rect 142540 77438 142660 77466
rect 142540 34134 142568 77438
rect 142620 77376 142672 77382
rect 142620 77318 142672 77324
rect 142632 60314 142660 77318
rect 142724 74254 142752 77590
rect 142712 74248 142764 74254
rect 142712 74190 142764 74196
rect 142712 74112 142764 74118
rect 142712 74054 142764 74060
rect 142724 65890 142752 74054
rect 142816 70922 142844 77710
rect 142896 77580 142948 77586
rect 142896 77522 142948 77528
rect 142908 71262 142936 77522
rect 143000 71754 143028 77710
rect 143124 77687 143180 77696
rect 143078 77616 143134 77625
rect 143230 77568 143258 78132
rect 143322 77926 143350 78132
rect 143310 77920 143362 77926
rect 143310 77862 143362 77868
rect 143414 77568 143442 78132
rect 143506 77858 143534 78132
rect 143494 77852 143546 77858
rect 143494 77794 143546 77800
rect 143598 77761 143626 78132
rect 143584 77752 143640 77761
rect 143584 77687 143640 77696
rect 143690 77704 143718 78132
rect 143782 77772 143810 78132
rect 143874 77926 143902 78132
rect 143966 77926 143994 78132
rect 144058 77926 144086 78132
rect 143862 77920 143914 77926
rect 143862 77862 143914 77868
rect 143954 77920 144006 77926
rect 143954 77862 144006 77868
rect 144046 77920 144098 77926
rect 144046 77862 144098 77868
rect 144150 77858 144178 78132
rect 144138 77852 144190 77858
rect 144138 77794 144190 77800
rect 143782 77744 143856 77772
rect 143690 77676 143764 77704
rect 143078 77551 143134 77560
rect 143092 73914 143120 77551
rect 143184 77540 143258 77568
rect 143368 77540 143442 77568
rect 143632 77580 143684 77586
rect 143184 74769 143212 77540
rect 143264 77444 143316 77450
rect 143264 77386 143316 77392
rect 143276 74905 143304 77386
rect 143262 74896 143318 74905
rect 143262 74831 143318 74840
rect 143170 74760 143226 74769
rect 143170 74695 143226 74704
rect 143368 74633 143396 77540
rect 143632 77522 143684 77528
rect 143448 77444 143500 77450
rect 143448 77386 143500 77392
rect 143460 74769 143488 77386
rect 143540 77308 143592 77314
rect 143540 77250 143592 77256
rect 143446 74760 143502 74769
rect 143446 74695 143502 74704
rect 143354 74624 143410 74633
rect 143354 74559 143410 74568
rect 143080 73908 143132 73914
rect 143080 73850 143132 73856
rect 143000 71726 143120 71754
rect 142988 71664 143040 71670
rect 142988 71606 143040 71612
rect 142896 71256 142948 71262
rect 142896 71198 142948 71204
rect 142804 70916 142856 70922
rect 142804 70858 142856 70864
rect 142804 69012 142856 69018
rect 142804 68954 142856 68960
rect 142712 65884 142764 65890
rect 142712 65826 142764 65832
rect 142620 60308 142672 60314
rect 142620 60250 142672 60256
rect 142528 34128 142580 34134
rect 142528 34070 142580 34076
rect 142436 28688 142488 28694
rect 142436 28630 142488 28636
rect 142344 28552 142396 28558
rect 142344 28494 142396 28500
rect 142252 20664 142304 20670
rect 142252 20606 142304 20612
rect 142160 6588 142212 6594
rect 142160 6530 142212 6536
rect 141240 4208 141292 4214
rect 141240 4150 141292 4156
rect 140044 3868 140096 3874
rect 140044 3810 140096 3816
rect 140136 3868 140188 3874
rect 140136 3810 140188 3816
rect 139952 3664 140004 3670
rect 139952 3606 140004 3612
rect 139032 3460 139084 3466
rect 139032 3402 139084 3408
rect 140056 480 140084 3810
rect 141252 480 141280 4150
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142264 354 142292 20606
rect 142816 3602 142844 68954
rect 143000 3806 143028 71606
rect 143092 71194 143120 71726
rect 143080 71188 143132 71194
rect 143080 71130 143132 71136
rect 143552 7818 143580 77250
rect 143644 77081 143672 77522
rect 143630 77072 143686 77081
rect 143630 77007 143686 77016
rect 143632 75676 143684 75682
rect 143632 75618 143684 75624
rect 143644 14754 143672 75618
rect 143736 75342 143764 77676
rect 143724 75336 143776 75342
rect 143724 75278 143776 75284
rect 143828 75002 143856 77744
rect 144092 77716 144144 77722
rect 144242 77704 144270 78132
rect 144334 77772 144362 78132
rect 144426 77926 144454 78132
rect 144518 77926 144546 78132
rect 144414 77920 144466 77926
rect 144414 77862 144466 77868
rect 144506 77920 144558 77926
rect 144506 77862 144558 77868
rect 144610 77772 144638 78132
rect 144334 77744 144408 77772
rect 144564 77761 144638 77772
rect 144242 77676 144316 77704
rect 144092 77658 144144 77664
rect 144000 77512 144052 77518
rect 144000 77454 144052 77460
rect 143908 77444 143960 77450
rect 143908 77386 143960 77392
rect 143816 74996 143868 75002
rect 143816 74938 143868 74944
rect 143816 74316 143868 74322
rect 143816 74258 143868 74264
rect 143724 73772 143776 73778
rect 143724 73714 143776 73720
rect 143736 20262 143764 73714
rect 143828 28490 143856 74258
rect 143920 30054 143948 77386
rect 144012 75426 144040 77454
rect 144104 75682 144132 77658
rect 144184 77580 144236 77586
rect 144184 77522 144236 77528
rect 144092 75676 144144 75682
rect 144092 75618 144144 75624
rect 144196 75528 144224 77522
rect 144288 76906 144316 77676
rect 144276 76900 144328 76906
rect 144276 76842 144328 76848
rect 144196 75500 144316 75528
rect 144012 75398 144224 75426
rect 144000 75336 144052 75342
rect 144000 75278 144052 75284
rect 144012 30122 144040 75278
rect 144092 74996 144144 75002
rect 144092 74938 144144 74944
rect 144104 34066 144132 74938
rect 144196 61878 144224 75398
rect 144184 61872 144236 61878
rect 144184 61814 144236 61820
rect 144288 61810 144316 75500
rect 144380 73778 144408 77744
rect 144550 77752 144638 77761
rect 144460 77716 144512 77722
rect 144606 77744 144638 77752
rect 144550 77687 144606 77696
rect 144460 77658 144512 77664
rect 144472 74322 144500 77658
rect 144552 77648 144604 77654
rect 144702 77636 144730 78132
rect 144794 77772 144822 78132
rect 144886 77897 144914 78132
rect 144872 77888 144928 77897
rect 144872 77823 144928 77832
rect 144794 77744 144868 77772
rect 144552 77590 144604 77596
rect 144656 77608 144730 77636
rect 144564 77353 144592 77590
rect 144550 77344 144606 77353
rect 144550 77279 144606 77288
rect 144552 76900 144604 76906
rect 144552 76842 144604 76848
rect 144460 74316 144512 74322
rect 144460 74258 144512 74264
rect 144564 74186 144592 76842
rect 144656 75041 144684 77608
rect 144840 77294 144868 77744
rect 144978 77466 145006 78132
rect 145070 77568 145098 78132
rect 145162 77858 145190 78132
rect 145254 77858 145282 78132
rect 145150 77852 145202 77858
rect 145150 77794 145202 77800
rect 145242 77852 145294 77858
rect 145242 77794 145294 77800
rect 145346 77790 145374 78132
rect 145438 77926 145466 78132
rect 145530 77926 145558 78132
rect 145622 77926 145650 78132
rect 145426 77920 145478 77926
rect 145426 77862 145478 77868
rect 145518 77920 145570 77926
rect 145518 77862 145570 77868
rect 145610 77920 145662 77926
rect 145610 77862 145662 77868
rect 145334 77784 145386 77790
rect 145610 77784 145662 77790
rect 145334 77726 145386 77732
rect 145608 77752 145610 77761
rect 145714 77772 145742 78132
rect 145806 77926 145834 78132
rect 145794 77920 145846 77926
rect 145794 77862 145846 77868
rect 145898 77772 145926 78132
rect 145662 77752 145664 77761
rect 145714 77744 145788 77772
rect 145852 77761 145926 77772
rect 145426 77716 145478 77722
rect 145478 77676 145558 77704
rect 145608 77687 145664 77696
rect 145426 77658 145478 77664
rect 145530 77602 145558 77676
rect 145196 77580 145248 77586
rect 145070 77540 145144 77568
rect 144978 77438 145052 77466
rect 144748 77266 144868 77294
rect 144920 77308 144972 77314
rect 144642 75032 144698 75041
rect 144642 74967 144698 74976
rect 144552 74180 144604 74186
rect 144552 74122 144604 74128
rect 144748 74089 144776 77266
rect 144920 77250 144972 77256
rect 144932 75177 144960 77250
rect 145024 75682 145052 77438
rect 145012 75676 145064 75682
rect 145012 75618 145064 75624
rect 144918 75168 144974 75177
rect 144918 75103 144974 75112
rect 145012 75132 145064 75138
rect 145116 75120 145144 77540
rect 145196 77522 145248 77528
rect 145380 77580 145432 77586
rect 145530 77574 145604 77602
rect 145380 77522 145432 77528
rect 145208 75614 145236 77522
rect 145288 77444 145340 77450
rect 145288 77386 145340 77392
rect 145196 75608 145248 75614
rect 145196 75550 145248 75556
rect 145116 75092 145236 75120
rect 145012 75074 145064 75080
rect 144920 74928 144972 74934
rect 144920 74870 144972 74876
rect 144734 74080 144790 74089
rect 144734 74015 144790 74024
rect 144368 73772 144420 73778
rect 144368 73714 144420 73720
rect 144460 73296 144512 73302
rect 144460 73238 144512 73244
rect 144276 61804 144328 61810
rect 144276 61746 144328 61752
rect 144092 34060 144144 34066
rect 144092 34002 144144 34008
rect 144000 30116 144052 30122
rect 144000 30058 144052 30064
rect 143908 30048 143960 30054
rect 143908 29990 143960 29996
rect 143816 28484 143868 28490
rect 143816 28426 143868 28432
rect 143724 20256 143776 20262
rect 143724 20198 143776 20204
rect 143632 14748 143684 14754
rect 143632 14690 143684 14696
rect 143540 7812 143592 7818
rect 143540 7754 143592 7760
rect 143540 4072 143592 4078
rect 143540 4014 143592 4020
rect 142988 3800 143040 3806
rect 142988 3742 143040 3748
rect 142804 3596 142856 3602
rect 142804 3538 142856 3544
rect 143552 480 143580 4014
rect 144472 3942 144500 73238
rect 144932 20398 144960 74870
rect 145024 27198 145052 75074
rect 145102 75032 145158 75041
rect 145102 74967 145158 74976
rect 145116 28422 145144 74967
rect 145208 29986 145236 75092
rect 145300 74984 145328 77386
rect 145392 75138 145420 77522
rect 145470 77480 145526 77489
rect 145470 77415 145472 77424
rect 145524 77415 145526 77424
rect 145472 77386 145524 77392
rect 145472 77308 145524 77314
rect 145472 77250 145524 77256
rect 145380 75132 145432 75138
rect 145380 75074 145432 75080
rect 145300 74956 145420 74984
rect 145288 74860 145340 74866
rect 145288 74802 145340 74808
rect 145300 33930 145328 74802
rect 145392 33998 145420 74956
rect 145484 74934 145512 77250
rect 145472 74928 145524 74934
rect 145472 74870 145524 74876
rect 145472 74792 145524 74798
rect 145472 74734 145524 74740
rect 145484 35630 145512 74734
rect 145576 63102 145604 77574
rect 145656 77512 145708 77518
rect 145656 77454 145708 77460
rect 145668 64462 145696 77454
rect 145760 74866 145788 77744
rect 145838 77752 145926 77761
rect 145894 77744 145926 77752
rect 145838 77687 145894 77696
rect 145990 77704 146018 78132
rect 146082 77926 146110 78132
rect 146070 77920 146122 77926
rect 146070 77862 146122 77868
rect 146174 77704 146202 78132
rect 146266 77761 146294 78132
rect 146358 77858 146386 78132
rect 146450 77858 146478 78132
rect 146346 77852 146398 77858
rect 146346 77794 146398 77800
rect 146438 77852 146490 77858
rect 146438 77794 146490 77800
rect 145990 77676 146064 77704
rect 145838 77616 145894 77625
rect 145838 77551 145840 77560
rect 145892 77551 145894 77560
rect 145840 77522 145892 77528
rect 145930 77480 145986 77489
rect 145840 77444 145892 77450
rect 145930 77415 145986 77424
rect 145840 77386 145892 77392
rect 145852 76265 145880 77386
rect 145838 76256 145894 76265
rect 145838 76191 145894 76200
rect 145748 74860 145800 74866
rect 145748 74802 145800 74808
rect 145944 74118 145972 77415
rect 146036 74798 146064 77676
rect 146128 77676 146202 77704
rect 146252 77752 146308 77761
rect 146252 77687 146308 77696
rect 146128 76401 146156 77676
rect 146298 77616 146354 77625
rect 146220 77574 146298 77602
rect 146114 76392 146170 76401
rect 146114 76327 146170 76336
rect 146024 74792 146076 74798
rect 146024 74734 146076 74740
rect 145932 74112 145984 74118
rect 145932 74054 145984 74060
rect 146220 71233 146248 77574
rect 146542 77568 146570 78132
rect 146634 77636 146662 78132
rect 146726 77926 146754 78132
rect 146714 77920 146766 77926
rect 146714 77862 146766 77868
rect 146818 77772 146846 78132
rect 146772 77744 146846 77772
rect 146910 77761 146938 78132
rect 147002 77790 147030 78132
rect 146990 77784 147042 77790
rect 146896 77752 146952 77761
rect 146634 77625 146708 77636
rect 146634 77616 146722 77625
rect 146634 77608 146666 77616
rect 146298 77551 146354 77560
rect 146496 77540 146570 77568
rect 146666 77551 146722 77560
rect 146392 77512 146444 77518
rect 146392 77454 146444 77460
rect 146300 77444 146352 77450
rect 146300 77386 146352 77392
rect 146312 76498 146340 77386
rect 146300 76492 146352 76498
rect 146300 76434 146352 76440
rect 146300 76356 146352 76362
rect 146300 76298 146352 76304
rect 146206 71224 146262 71233
rect 146206 71159 146262 71168
rect 145656 64456 145708 64462
rect 145656 64398 145708 64404
rect 145564 63096 145616 63102
rect 145564 63038 145616 63044
rect 145472 35624 145524 35630
rect 145472 35566 145524 35572
rect 145380 33992 145432 33998
rect 145380 33934 145432 33940
rect 145288 33924 145340 33930
rect 145288 33866 145340 33872
rect 145196 29980 145248 29986
rect 145196 29922 145248 29928
rect 145104 28416 145156 28422
rect 145104 28358 145156 28364
rect 145012 27192 145064 27198
rect 145012 27134 145064 27140
rect 144920 20392 144972 20398
rect 144920 20334 144972 20340
rect 144920 9240 144972 9246
rect 144920 9182 144972 9188
rect 144736 4140 144788 4146
rect 144736 4082 144788 4088
rect 144460 3936 144512 3942
rect 144460 3878 144512 3884
rect 144748 480 144776 4082
rect 144932 3738 144960 9182
rect 146312 6526 146340 76298
rect 146404 76158 146432 77454
rect 146392 76152 146444 76158
rect 146392 76094 146444 76100
rect 146392 73976 146444 73982
rect 146392 73918 146444 73924
rect 146404 7750 146432 73918
rect 146496 20330 146524 77540
rect 146668 77512 146720 77518
rect 146574 77480 146630 77489
rect 146668 77454 146720 77460
rect 146574 77415 146630 77424
rect 146588 76226 146616 77415
rect 146576 76220 146628 76226
rect 146576 76162 146628 76168
rect 146576 76084 146628 76090
rect 146576 76026 146628 76032
rect 146588 73794 146616 76026
rect 146680 73982 146708 77454
rect 146772 76242 146800 77744
rect 146990 77726 147042 77732
rect 146896 77687 146952 77696
rect 147094 77704 147122 78132
rect 147186 77926 147214 78132
rect 147278 77926 147306 78132
rect 147370 77926 147398 78132
rect 147462 77926 147490 78132
rect 147554 77926 147582 78132
rect 147646 77926 147674 78132
rect 147738 77926 147766 78132
rect 147174 77920 147226 77926
rect 147174 77862 147226 77868
rect 147266 77920 147318 77926
rect 147266 77862 147318 77868
rect 147358 77920 147410 77926
rect 147358 77862 147410 77868
rect 147450 77920 147502 77926
rect 147450 77862 147502 77868
rect 147542 77920 147594 77926
rect 147542 77862 147594 77868
rect 147634 77920 147686 77926
rect 147634 77862 147686 77868
rect 147726 77920 147778 77926
rect 147726 77862 147778 77868
rect 147220 77784 147272 77790
rect 147220 77726 147272 77732
rect 147680 77784 147732 77790
rect 147830 77772 147858 78132
rect 147680 77726 147732 77732
rect 147784 77744 147858 77772
rect 147094 77676 147168 77704
rect 146852 77648 146904 77654
rect 146852 77590 146904 77596
rect 147034 77616 147090 77625
rect 146864 76362 146892 77590
rect 146944 77580 146996 77586
rect 147034 77551 147090 77560
rect 146944 77522 146996 77528
rect 146956 76906 146984 77522
rect 146944 76900 146996 76906
rect 146944 76842 146996 76848
rect 146852 76356 146904 76362
rect 146852 76298 146904 76304
rect 146772 76214 146984 76242
rect 146760 76152 146812 76158
rect 146760 76094 146812 76100
rect 146668 73976 146720 73982
rect 146668 73918 146720 73924
rect 146588 73766 146708 73794
rect 146576 73432 146628 73438
rect 146576 73374 146628 73380
rect 146588 25770 146616 73374
rect 146680 27130 146708 73766
rect 146772 29918 146800 76094
rect 146852 70780 146904 70786
rect 146852 70722 146904 70728
rect 146864 35494 146892 70722
rect 146956 35562 146984 76214
rect 147048 61742 147076 77551
rect 147140 70786 147168 77676
rect 147232 73438 147260 77726
rect 147312 77716 147364 77722
rect 147312 77658 147364 77664
rect 147404 77716 147456 77722
rect 147404 77658 147456 77664
rect 147324 76809 147352 77658
rect 147310 76800 147366 76809
rect 147310 76735 147366 76744
rect 147312 76220 147364 76226
rect 147312 76162 147364 76168
rect 147220 73432 147272 73438
rect 147220 73374 147272 73380
rect 147128 70780 147180 70786
rect 147128 70722 147180 70728
rect 147324 69014 147352 76162
rect 147416 73545 147444 77658
rect 147496 77648 147548 77654
rect 147496 77590 147548 77596
rect 147508 74338 147536 77590
rect 147588 77240 147640 77246
rect 147588 77182 147640 77188
rect 147600 76838 147628 77182
rect 147588 76832 147640 76838
rect 147588 76774 147640 76780
rect 147692 76158 147720 77726
rect 147680 76152 147732 76158
rect 147680 76094 147732 76100
rect 147680 75064 147732 75070
rect 147680 75006 147732 75012
rect 147692 74610 147720 75006
rect 147784 74780 147812 77744
rect 147922 77704 147950 78132
rect 148014 77926 148042 78132
rect 148002 77920 148054 77926
rect 148002 77862 148054 77868
rect 148106 77704 148134 78132
rect 147876 77676 147950 77704
rect 148060 77676 148134 77704
rect 147876 74934 147904 77676
rect 147956 77580 148008 77586
rect 147956 77522 148008 77528
rect 147968 75002 147996 77522
rect 147956 74996 148008 75002
rect 147956 74938 148008 74944
rect 147864 74928 147916 74934
rect 147864 74870 147916 74876
rect 147784 74752 147996 74780
rect 147692 74582 147812 74610
rect 147508 74310 147628 74338
rect 147496 74248 147548 74254
rect 147496 74190 147548 74196
rect 147508 73914 147536 74190
rect 147600 73953 147628 74310
rect 147680 74316 147732 74322
rect 147680 74258 147732 74264
rect 147586 73944 147642 73953
rect 147496 73908 147548 73914
rect 147586 73879 147642 73888
rect 147496 73850 147548 73856
rect 147402 73536 147458 73545
rect 147402 73471 147458 73480
rect 147140 68986 147352 69014
rect 147140 64394 147168 68986
rect 147128 64388 147180 64394
rect 147128 64330 147180 64336
rect 147036 61736 147088 61742
rect 147036 61678 147088 61684
rect 146944 35556 146996 35562
rect 146944 35498 146996 35504
rect 146852 35488 146904 35494
rect 146852 35430 146904 35436
rect 146760 29912 146812 29918
rect 146760 29854 146812 29860
rect 146668 27124 146720 27130
rect 146668 27066 146720 27072
rect 146576 25764 146628 25770
rect 146576 25706 146628 25712
rect 146484 20324 146536 20330
rect 146484 20266 146536 20272
rect 146392 7744 146444 7750
rect 146392 7686 146444 7692
rect 147692 7682 147720 74258
rect 147784 13598 147812 74582
rect 147864 71120 147916 71126
rect 147864 71062 147916 71068
rect 147876 16182 147904 71062
rect 147968 29850 147996 74752
rect 147956 29844 148008 29850
rect 147956 29786 148008 29792
rect 148060 29782 148088 77676
rect 148198 77636 148226 78132
rect 148290 77926 148318 78132
rect 148382 77926 148410 78132
rect 148474 77926 148502 78132
rect 148566 77926 148594 78132
rect 148278 77920 148330 77926
rect 148278 77862 148330 77868
rect 148370 77920 148422 77926
rect 148370 77862 148422 77868
rect 148462 77920 148514 77926
rect 148462 77862 148514 77868
rect 148554 77920 148606 77926
rect 148554 77862 148606 77868
rect 148324 77784 148376 77790
rect 148658 77772 148686 78132
rect 148750 77926 148778 78132
rect 148842 77926 148870 78132
rect 148934 77926 148962 78132
rect 149026 77926 149054 78132
rect 148738 77920 148790 77926
rect 148738 77862 148790 77868
rect 148830 77920 148882 77926
rect 148830 77862 148882 77868
rect 148922 77920 148974 77926
rect 148922 77862 148974 77868
rect 149014 77920 149066 77926
rect 149014 77862 149066 77868
rect 149118 77772 149146 78132
rect 149210 77926 149238 78132
rect 149302 77926 149330 78132
rect 149394 77926 149422 78132
rect 149486 77926 149514 78132
rect 149198 77920 149250 77926
rect 149198 77862 149250 77868
rect 149290 77920 149342 77926
rect 149290 77862 149342 77868
rect 149382 77920 149434 77926
rect 149382 77862 149434 77868
rect 149474 77920 149526 77926
rect 149474 77862 149526 77868
rect 149244 77784 149296 77790
rect 148376 77744 148456 77772
rect 148658 77761 148732 77772
rect 148658 77752 148746 77761
rect 148658 77744 148690 77752
rect 148324 77726 148376 77732
rect 148152 77608 148226 77636
rect 148324 77648 148376 77654
rect 148152 75070 148180 77608
rect 148324 77590 148376 77596
rect 148232 77444 148284 77450
rect 148232 77386 148284 77392
rect 148140 75064 148192 75070
rect 148140 75006 148192 75012
rect 148140 74928 148192 74934
rect 148140 74870 148192 74876
rect 148152 35426 148180 74870
rect 148244 71126 148272 77386
rect 148232 71120 148284 71126
rect 148232 71062 148284 71068
rect 148232 70780 148284 70786
rect 148232 70722 148284 70728
rect 148244 54602 148272 70722
rect 148336 60246 148364 77590
rect 148428 74322 148456 77744
rect 149118 77744 149192 77772
rect 148690 77687 148746 77696
rect 148784 77716 148836 77722
rect 148784 77658 148836 77664
rect 148876 77716 148928 77722
rect 148876 77658 148928 77664
rect 148968 77716 149020 77722
rect 148968 77658 149020 77664
rect 148598 77616 148654 77625
rect 148598 77551 148654 77560
rect 148692 77580 148744 77586
rect 148508 77376 148560 77382
rect 148508 77318 148560 77324
rect 148416 74316 148468 74322
rect 148416 74258 148468 74264
rect 148520 70786 148548 77318
rect 148612 76022 148640 77551
rect 148692 77522 148744 77528
rect 148600 76016 148652 76022
rect 148600 75958 148652 75964
rect 148600 75404 148652 75410
rect 148600 75346 148652 75352
rect 148508 70780 148560 70786
rect 148508 70722 148560 70728
rect 148612 70394 148640 75346
rect 148704 70530 148732 77522
rect 148796 75041 148824 77658
rect 148888 75721 148916 77658
rect 148874 75712 148930 75721
rect 148874 75647 148930 75656
rect 148782 75032 148838 75041
rect 148782 74967 148838 74976
rect 148980 74633 149008 77658
rect 149058 77344 149114 77353
rect 149058 77279 149060 77288
rect 149112 77279 149114 77288
rect 149060 77250 149112 77256
rect 149164 77246 149192 77744
rect 149244 77726 149296 77732
rect 149152 77240 149204 77246
rect 149152 77182 149204 77188
rect 149152 75540 149204 75546
rect 149152 75482 149204 75488
rect 148966 74624 149022 74633
rect 148966 74559 149022 74568
rect 148704 70502 149100 70530
rect 148612 70366 149008 70394
rect 148980 68610 149008 70366
rect 149072 69737 149100 70502
rect 149058 69728 149114 69737
rect 149058 69663 149114 69672
rect 149060 69624 149112 69630
rect 149060 69566 149112 69572
rect 148968 68604 149020 68610
rect 148968 68546 149020 68552
rect 148324 60240 148376 60246
rect 148324 60182 148376 60188
rect 148232 54596 148284 54602
rect 148232 54538 148284 54544
rect 148140 35420 148192 35426
rect 148140 35362 148192 35368
rect 148048 29776 148100 29782
rect 148048 29718 148100 29724
rect 147864 16176 147916 16182
rect 147864 16118 147916 16124
rect 147772 13592 147824 13598
rect 147772 13534 147824 13540
rect 149072 9246 149100 69566
rect 149060 9240 149112 9246
rect 149060 9182 149112 9188
rect 149164 9178 149192 75482
rect 149256 73438 149284 77726
rect 149336 77716 149388 77722
rect 149336 77658 149388 77664
rect 149428 77716 149480 77722
rect 149428 77658 149480 77664
rect 149348 77489 149376 77658
rect 149334 77480 149390 77489
rect 149334 77415 149390 77424
rect 149336 77376 149388 77382
rect 149336 77318 149388 77324
rect 149244 73432 149296 73438
rect 149244 73374 149296 73380
rect 149244 73296 149296 73302
rect 149244 73238 149296 73244
rect 149256 10742 149284 73238
rect 149348 31550 149376 77318
rect 149336 31544 149388 31550
rect 149336 31486 149388 31492
rect 149440 31482 149468 77658
rect 149578 77602 149606 78132
rect 149670 77790 149698 78132
rect 149762 77926 149790 78132
rect 149854 77926 149882 78132
rect 149946 77926 149974 78132
rect 149750 77920 149802 77926
rect 149750 77862 149802 77868
rect 149842 77920 149894 77926
rect 149842 77862 149894 77868
rect 149934 77920 149986 77926
rect 149934 77862 149986 77868
rect 149658 77784 149710 77790
rect 149658 77726 149710 77732
rect 149796 77784 149848 77790
rect 149796 77726 149848 77732
rect 149888 77784 149940 77790
rect 150038 77772 150066 78132
rect 150130 77926 150158 78132
rect 150118 77920 150170 77926
rect 150118 77862 150170 77868
rect 150038 77744 150112 77772
rect 149888 77726 149940 77732
rect 149532 77574 149606 77602
rect 149704 77648 149756 77654
rect 149704 77590 149756 77596
rect 149532 35358 149560 77574
rect 149612 77512 149664 77518
rect 149612 77454 149664 77460
rect 149624 75138 149652 77454
rect 149612 75132 149664 75138
rect 149612 75074 149664 75080
rect 149612 71596 149664 71602
rect 149612 71538 149664 71544
rect 149624 53106 149652 71538
rect 149716 60178 149744 77590
rect 149808 75290 149836 77726
rect 149900 75546 149928 77726
rect 149980 77580 150032 77586
rect 149980 77522 150032 77528
rect 149992 75721 150020 77522
rect 149978 75712 150034 75721
rect 149978 75647 150034 75656
rect 149888 75540 149940 75546
rect 149888 75482 149940 75488
rect 149808 75262 149928 75290
rect 149796 75132 149848 75138
rect 149796 75074 149848 75080
rect 149808 69630 149836 75074
rect 149900 69970 149928 75262
rect 150084 73302 150112 77744
rect 150222 77738 150250 78132
rect 150314 77926 150342 78132
rect 150406 77926 150434 78132
rect 150498 77926 150526 78132
rect 150590 77926 150618 78132
rect 150302 77920 150354 77926
rect 150302 77862 150354 77868
rect 150394 77920 150446 77926
rect 150394 77862 150446 77868
rect 150486 77920 150538 77926
rect 150486 77862 150538 77868
rect 150578 77920 150630 77926
rect 150578 77862 150630 77868
rect 150348 77784 150400 77790
rect 150222 77710 150296 77738
rect 150682 77772 150710 78132
rect 150348 77726 150400 77732
rect 150636 77744 150710 77772
rect 150164 77648 150216 77654
rect 150164 77590 150216 77596
rect 150176 76265 150204 77590
rect 150162 76256 150218 76265
rect 150162 76191 150218 76200
rect 150164 76152 150216 76158
rect 150164 76094 150216 76100
rect 150072 73296 150124 73302
rect 150072 73238 150124 73244
rect 149888 69964 149940 69970
rect 149888 69906 149940 69912
rect 150176 69873 150204 76094
rect 150268 71602 150296 77710
rect 150256 71596 150308 71602
rect 150256 71538 150308 71544
rect 150162 69864 150218 69873
rect 150162 69799 150218 69808
rect 149980 69692 150032 69698
rect 149980 69634 150032 69640
rect 149796 69624 149848 69630
rect 149796 69566 149848 69572
rect 149704 60172 149756 60178
rect 149704 60114 149756 60120
rect 149612 53100 149664 53106
rect 149612 53042 149664 53048
rect 149520 35352 149572 35358
rect 149520 35294 149572 35300
rect 149428 31476 149480 31482
rect 149428 31418 149480 31424
rect 149244 10736 149296 10742
rect 149244 10678 149296 10684
rect 149152 9172 149204 9178
rect 149152 9114 149204 9120
rect 147680 7676 147732 7682
rect 147680 7618 147732 7624
rect 146300 6520 146352 6526
rect 146300 6462 146352 6468
rect 148324 5160 148376 5166
rect 148324 5102 148376 5108
rect 145932 4004 145984 4010
rect 145932 3946 145984 3952
rect 144920 3732 144972 3738
rect 144920 3674 144972 3680
rect 145944 480 145972 3946
rect 147128 3528 147180 3534
rect 147128 3470 147180 3476
rect 147140 480 147168 3470
rect 148336 480 148364 5102
rect 149520 3868 149572 3874
rect 149520 3810 149572 3816
rect 149532 480 149560 3810
rect 149992 3738 150020 69634
rect 150360 69601 150388 77726
rect 150532 77716 150584 77722
rect 150532 77658 150584 77664
rect 150438 77344 150494 77353
rect 150438 77279 150494 77288
rect 150452 75614 150480 77279
rect 150440 75608 150492 75614
rect 150440 75550 150492 75556
rect 150544 75546 150572 77658
rect 150532 75540 150584 75546
rect 150532 75482 150584 75488
rect 150440 75064 150492 75070
rect 150440 75006 150492 75012
rect 150346 69592 150402 69601
rect 150346 69527 150402 69536
rect 150452 69014 150480 75006
rect 150452 68986 150572 69014
rect 150544 10674 150572 68986
rect 150636 18970 150664 77744
rect 150774 77704 150802 78132
rect 150728 77676 150802 77704
rect 150728 75614 150756 77676
rect 150866 77636 150894 78132
rect 150958 77897 150986 78132
rect 151050 77926 151078 78132
rect 151142 77926 151170 78132
rect 151038 77920 151090 77926
rect 150944 77888 151000 77897
rect 151038 77862 151090 77868
rect 151130 77920 151182 77926
rect 151130 77862 151182 77868
rect 150944 77823 151000 77832
rect 151234 77772 151262 78132
rect 151326 77926 151354 78132
rect 151314 77920 151366 77926
rect 151314 77862 151366 77868
rect 151418 77772 151446 78132
rect 151510 77926 151538 78132
rect 151498 77920 151550 77926
rect 151498 77862 151550 77868
rect 151602 77772 151630 78132
rect 151694 77897 151722 78132
rect 151786 77926 151814 78132
rect 151878 77926 151906 78132
rect 151774 77920 151826 77926
rect 151680 77888 151736 77897
rect 151774 77862 151826 77868
rect 151866 77920 151918 77926
rect 151866 77862 151918 77868
rect 151680 77823 151736 77832
rect 151082 77752 151138 77761
rect 150992 77716 151044 77722
rect 151234 77744 151308 77772
rect 151082 77687 151138 77696
rect 150992 77658 151044 77664
rect 150820 77608 150894 77636
rect 150716 75608 150768 75614
rect 150716 75550 150768 75556
rect 150716 72616 150768 72622
rect 150716 72558 150768 72564
rect 150728 23186 150756 72558
rect 150820 24478 150848 77608
rect 150900 75540 150952 75546
rect 150900 75482 150952 75488
rect 150912 31414 150940 75482
rect 151004 75070 151032 77658
rect 151096 75698 151124 77687
rect 151176 77648 151228 77654
rect 151176 77590 151228 77596
rect 151188 75857 151216 77590
rect 151174 75848 151230 75857
rect 151174 75783 151230 75792
rect 151096 75670 151216 75698
rect 151084 75608 151136 75614
rect 151084 75550 151136 75556
rect 150992 75064 151044 75070
rect 150992 75006 151044 75012
rect 150992 70508 151044 70514
rect 150992 70450 151044 70456
rect 151004 61674 151032 70450
rect 151096 64326 151124 75550
rect 151188 69902 151216 75670
rect 151280 72622 151308 77744
rect 151372 77744 151446 77772
rect 151556 77744 151630 77772
rect 151728 77784 151780 77790
rect 151372 77704 151400 77744
rect 151372 77676 151492 77704
rect 151360 77580 151412 77586
rect 151360 77522 151412 77528
rect 151268 72616 151320 72622
rect 151268 72558 151320 72564
rect 151372 70514 151400 77522
rect 151464 72146 151492 77676
rect 151556 75721 151584 77744
rect 151970 77738 151998 78132
rect 152062 77897 152090 78132
rect 152154 77926 152182 78132
rect 152142 77920 152194 77926
rect 152048 77888 152104 77897
rect 152142 77862 152194 77868
rect 152048 77823 152104 77832
rect 152246 77738 152274 78132
rect 152338 77897 152366 78132
rect 152430 77926 152458 78132
rect 152522 77926 152550 78132
rect 152418 77920 152470 77926
rect 152324 77888 152380 77897
rect 152418 77862 152470 77868
rect 152510 77920 152562 77926
rect 152614 77897 152642 78132
rect 152706 77926 152734 78132
rect 152694 77920 152746 77926
rect 152510 77862 152562 77868
rect 152600 77888 152656 77897
rect 152324 77823 152380 77832
rect 152798 77897 152826 78132
rect 152890 77926 152918 78132
rect 152982 77926 153010 78132
rect 153074 77926 153102 78132
rect 152878 77920 152930 77926
rect 152694 77862 152746 77868
rect 152784 77888 152840 77897
rect 152600 77823 152656 77832
rect 152878 77862 152930 77868
rect 152970 77920 153022 77926
rect 152970 77862 153022 77868
rect 153062 77920 153114 77926
rect 153062 77862 153114 77868
rect 152784 77823 152840 77832
rect 151728 77726 151780 77732
rect 151740 77294 151768 77726
rect 151820 77716 151872 77722
rect 151820 77658 151872 77664
rect 151924 77710 151998 77738
rect 152108 77710 152274 77738
rect 152738 77752 152794 77761
rect 152464 77716 152516 77722
rect 151648 77266 151768 77294
rect 151542 75712 151598 75721
rect 151542 75647 151598 75656
rect 151542 75576 151598 75585
rect 151542 75511 151598 75520
rect 151452 72140 151504 72146
rect 151452 72082 151504 72088
rect 151360 70508 151412 70514
rect 151360 70450 151412 70456
rect 151176 69896 151228 69902
rect 151176 69838 151228 69844
rect 151084 64320 151136 64326
rect 151084 64262 151136 64268
rect 150992 61668 151044 61674
rect 150992 61610 151044 61616
rect 150900 31408 150952 31414
rect 150900 31350 150952 31356
rect 150808 24472 150860 24478
rect 150808 24414 150860 24420
rect 150716 23180 150768 23186
rect 150716 23122 150768 23128
rect 150624 18964 150676 18970
rect 150624 18906 150676 18912
rect 150532 10668 150584 10674
rect 150532 10610 150584 10616
rect 150624 5364 150676 5370
rect 150624 5306 150676 5312
rect 149980 3732 150032 3738
rect 149980 3674 150032 3680
rect 150636 480 150664 5306
rect 151556 5234 151584 75511
rect 151648 73154 151676 77266
rect 151832 75138 151860 77658
rect 151820 75132 151872 75138
rect 151820 75074 151872 75080
rect 151924 74984 151952 77710
rect 152004 77512 152056 77518
rect 152004 77454 152056 77460
rect 152016 76838 152044 77454
rect 152004 76832 152056 76838
rect 152004 76774 152056 76780
rect 151924 74956 152044 74984
rect 151912 73772 151964 73778
rect 151912 73714 151964 73720
rect 151648 73126 151768 73154
rect 151740 72865 151768 73126
rect 151726 72856 151782 72865
rect 151726 72791 151782 72800
rect 151820 70508 151872 70514
rect 151820 70450 151872 70456
rect 151832 10606 151860 70450
rect 151924 11966 151952 73714
rect 152016 13530 152044 74956
rect 152108 14686 152136 77710
rect 152738 77687 152794 77696
rect 152832 77716 152884 77722
rect 152464 77658 152516 77664
rect 152188 77648 152240 77654
rect 152188 77590 152240 77596
rect 152200 75698 152228 77590
rect 152280 77580 152332 77586
rect 152280 77522 152332 77528
rect 152292 75857 152320 77522
rect 152372 77308 152424 77314
rect 152372 77250 152424 77256
rect 152384 76634 152412 77250
rect 152372 76628 152424 76634
rect 152372 76570 152424 76576
rect 152278 75848 152334 75857
rect 152278 75783 152334 75792
rect 152200 75670 152412 75698
rect 152278 75576 152334 75585
rect 152278 75511 152334 75520
rect 152188 73364 152240 73370
rect 152188 73306 152240 73312
rect 152200 25702 152228 73306
rect 152292 55894 152320 75511
rect 152384 62966 152412 75670
rect 152476 70514 152504 77658
rect 152556 77648 152608 77654
rect 152556 77590 152608 77596
rect 152568 73370 152596 77590
rect 152648 77580 152700 77586
rect 152648 77522 152700 77528
rect 152660 73778 152688 77522
rect 152752 75290 152780 77687
rect 152832 77658 152884 77664
rect 152924 77716 152976 77722
rect 153166 77704 153194 78132
rect 153258 77926 153286 78132
rect 153246 77920 153298 77926
rect 153246 77862 153298 77868
rect 153350 77772 153378 78132
rect 153442 77897 153470 78132
rect 153428 77888 153484 77897
rect 153428 77823 153484 77832
rect 152924 77658 152976 77664
rect 153120 77676 153194 77704
rect 153304 77744 153378 77772
rect 152844 76129 152872 77658
rect 152830 76120 152886 76129
rect 152830 76055 152886 76064
rect 152830 75984 152886 75993
rect 152830 75919 152832 75928
rect 152884 75919 152886 75928
rect 152832 75890 152884 75896
rect 152936 75721 152964 77658
rect 153120 77602 153148 77676
rect 153074 77574 153148 77602
rect 153198 77616 153254 77625
rect 153074 77466 153102 77574
rect 153198 77551 153200 77560
rect 153252 77551 153254 77560
rect 153200 77522 153252 77528
rect 153074 77438 153148 77466
rect 153120 76158 153148 77438
rect 153198 76800 153254 76809
rect 153198 76735 153254 76744
rect 153108 76152 153160 76158
rect 153108 76094 153160 76100
rect 152922 75712 152978 75721
rect 152922 75647 152978 75656
rect 152924 75540 152976 75546
rect 152924 75482 152976 75488
rect 152752 75262 152872 75290
rect 152740 75200 152792 75206
rect 152740 75142 152792 75148
rect 152648 73772 152700 73778
rect 152648 73714 152700 73720
rect 152648 73432 152700 73438
rect 152648 73374 152700 73380
rect 152556 73364 152608 73370
rect 152556 73306 152608 73312
rect 152464 70508 152516 70514
rect 152464 70450 152516 70456
rect 152660 70038 152688 73374
rect 152752 70394 152780 75142
rect 152844 73506 152872 75262
rect 152832 73500 152884 73506
rect 152832 73442 152884 73448
rect 152936 72690 152964 75482
rect 153108 75268 153160 75274
rect 153108 75210 153160 75216
rect 153120 74322 153148 75210
rect 153108 74316 153160 74322
rect 153108 74258 153160 74264
rect 152924 72684 152976 72690
rect 152924 72626 152976 72632
rect 152752 70366 152872 70394
rect 152648 70032 152700 70038
rect 152648 69974 152700 69980
rect 152372 62960 152424 62966
rect 152372 62902 152424 62908
rect 152280 55888 152332 55894
rect 152280 55830 152332 55836
rect 152188 25696 152240 25702
rect 152188 25638 152240 25644
rect 152096 14680 152148 14686
rect 152096 14622 152148 14628
rect 152004 13524 152056 13530
rect 152004 13466 152056 13472
rect 151912 11960 151964 11966
rect 151912 11902 151964 11908
rect 151820 10600 151872 10606
rect 151820 10542 151872 10548
rect 151544 5228 151596 5234
rect 151544 5170 151596 5176
rect 151820 5092 151872 5098
rect 151820 5034 151872 5040
rect 151832 480 151860 5034
rect 152844 3194 152872 70366
rect 153212 5166 153240 76735
rect 153304 75410 153332 77744
rect 153534 77738 153562 78132
rect 153488 77710 153562 77738
rect 153384 77512 153436 77518
rect 153384 77454 153436 77460
rect 153292 75404 153344 75410
rect 153292 75346 153344 75352
rect 153290 75304 153346 75313
rect 153290 75239 153346 75248
rect 153304 9110 153332 75239
rect 153396 11762 153424 77454
rect 153488 75886 153516 77710
rect 153626 77636 153654 78132
rect 153718 77897 153746 78132
rect 153704 77888 153760 77897
rect 153810 77858 153838 78132
rect 153902 77926 153930 78132
rect 153890 77920 153942 77926
rect 153890 77862 153942 77868
rect 153704 77823 153760 77832
rect 153798 77852 153850 77858
rect 153798 77794 153850 77800
rect 153994 77772 154022 78132
rect 154086 77897 154114 78132
rect 154072 77888 154128 77897
rect 154178 77858 154206 78132
rect 154270 77858 154298 78132
rect 154072 77823 154128 77832
rect 154166 77852 154218 77858
rect 154166 77794 154218 77800
rect 154258 77852 154310 77858
rect 154258 77794 154310 77800
rect 153994 77744 154068 77772
rect 153752 77716 153804 77722
rect 153752 77658 153804 77664
rect 153580 77608 153654 77636
rect 153476 75880 153528 75886
rect 153476 75822 153528 75828
rect 153476 75608 153528 75614
rect 153476 75550 153528 75556
rect 153488 11830 153516 75550
rect 153580 11898 153608 77608
rect 153658 76256 153714 76265
rect 153658 76191 153714 76200
rect 153672 13462 153700 76191
rect 153764 75614 153792 77658
rect 153936 77648 153988 77654
rect 153936 77590 153988 77596
rect 153842 77208 153898 77217
rect 153842 77143 153898 77152
rect 153856 75614 153884 77143
rect 153948 75970 153976 77590
rect 154040 76401 154068 77744
rect 154362 77738 154390 78132
rect 154120 77716 154172 77722
rect 154120 77658 154172 77664
rect 154316 77710 154390 77738
rect 154132 76809 154160 77658
rect 154210 77616 154266 77625
rect 154210 77551 154266 77560
rect 154118 76800 154174 76809
rect 154118 76735 154174 76744
rect 154026 76392 154082 76401
rect 154026 76327 154082 76336
rect 153948 75942 154068 75970
rect 153936 75880 153988 75886
rect 153936 75822 153988 75828
rect 153752 75608 153804 75614
rect 153752 75550 153804 75556
rect 153844 75608 153896 75614
rect 153844 75550 153896 75556
rect 153752 75404 153804 75410
rect 153752 75346 153804 75352
rect 153764 27062 153792 75346
rect 153844 75200 153896 75206
rect 153844 75142 153896 75148
rect 153856 60110 153884 75142
rect 153948 61606 153976 75822
rect 154040 75206 154068 75942
rect 154120 75948 154172 75954
rect 154120 75890 154172 75896
rect 154028 75200 154080 75206
rect 154028 75142 154080 75148
rect 154026 75032 154082 75041
rect 154026 74967 154082 74976
rect 154040 69766 154068 74967
rect 154132 71398 154160 75890
rect 154224 75857 154252 77551
rect 154210 75848 154266 75857
rect 154210 75783 154266 75792
rect 154316 75721 154344 77710
rect 154454 77602 154482 78132
rect 154546 77897 154574 78132
rect 154532 77888 154588 77897
rect 154532 77823 154588 77832
rect 154638 77772 154666 78132
rect 154592 77744 154666 77772
rect 154454 77574 154528 77602
rect 154396 77512 154448 77518
rect 154396 77454 154448 77460
rect 154302 75712 154358 75721
rect 154302 75647 154358 75656
rect 154408 75274 154436 77454
rect 154500 75585 154528 77574
rect 154486 75576 154542 75585
rect 154486 75511 154542 75520
rect 154396 75268 154448 75274
rect 154396 75210 154448 75216
rect 154488 75132 154540 75138
rect 154488 75074 154540 75080
rect 154212 72140 154264 72146
rect 154212 72082 154264 72088
rect 154120 71392 154172 71398
rect 154120 71334 154172 71340
rect 154028 69760 154080 69766
rect 154028 69702 154080 69708
rect 154224 65822 154252 72082
rect 154500 69834 154528 75074
rect 154592 74730 154620 77744
rect 154730 77466 154758 78132
rect 154822 77926 154850 78132
rect 154810 77920 154862 77926
rect 154810 77862 154862 77868
rect 154914 77772 154942 78132
rect 155006 77897 155034 78132
rect 154992 77888 155048 77897
rect 154992 77823 155048 77832
rect 155098 77772 155126 78132
rect 154868 77744 154942 77772
rect 155052 77744 155126 77772
rect 154730 77438 154804 77466
rect 154672 77376 154724 77382
rect 154672 77318 154724 77324
rect 154684 76702 154712 77318
rect 154672 76696 154724 76702
rect 154672 76638 154724 76644
rect 154672 75880 154724 75886
rect 154672 75822 154724 75828
rect 154580 74724 154632 74730
rect 154580 74666 154632 74672
rect 154684 73154 154712 75822
rect 154776 75698 154804 77438
rect 154868 77382 154896 77744
rect 154948 77648 155000 77654
rect 154948 77590 155000 77596
rect 154856 77376 154908 77382
rect 154856 77318 154908 77324
rect 154854 77072 154910 77081
rect 154854 77007 154910 77016
rect 154868 75857 154896 77007
rect 154854 75848 154910 75857
rect 154854 75783 154910 75792
rect 154776 75670 154896 75698
rect 154762 75576 154818 75585
rect 154762 75511 154818 75520
rect 154592 73126 154712 73154
rect 154488 69828 154540 69834
rect 154488 69770 154540 69776
rect 154212 65816 154264 65822
rect 154212 65758 154264 65764
rect 153936 61600 153988 61606
rect 153936 61542 153988 61548
rect 153844 60104 153896 60110
rect 153844 60046 153896 60052
rect 153752 27056 153804 27062
rect 153752 26998 153804 27004
rect 153660 13456 153712 13462
rect 153660 13398 153712 13404
rect 154592 13394 154620 73126
rect 154672 71868 154724 71874
rect 154672 71810 154724 71816
rect 154684 14618 154712 71810
rect 154776 16114 154804 75511
rect 154868 29714 154896 75670
rect 154960 75546 154988 77590
rect 154948 75540 155000 75546
rect 154948 75482 155000 75488
rect 154948 72548 155000 72554
rect 154948 72490 155000 72496
rect 154960 31346 154988 72490
rect 155052 35290 155080 77744
rect 155190 77704 155218 78132
rect 155282 77926 155310 78132
rect 155374 77926 155402 78132
rect 155466 77926 155494 78132
rect 155270 77920 155322 77926
rect 155270 77862 155322 77868
rect 155362 77920 155414 77926
rect 155362 77862 155414 77868
rect 155454 77920 155506 77926
rect 155454 77862 155506 77868
rect 155558 77772 155586 78132
rect 155512 77744 155586 77772
rect 155650 77772 155678 78132
rect 155742 77926 155770 78132
rect 155834 77926 155862 78132
rect 155926 77931 155954 78132
rect 155730 77920 155782 77926
rect 155730 77862 155782 77868
rect 155822 77920 155874 77926
rect 155822 77862 155874 77868
rect 155912 77922 155968 77931
rect 155912 77857 155968 77866
rect 155868 77784 155920 77790
rect 155650 77744 155816 77772
rect 155144 77676 155218 77704
rect 155408 77716 155460 77722
rect 155144 75886 155172 77676
rect 155408 77658 155460 77664
rect 155224 77580 155276 77586
rect 155224 77522 155276 77528
rect 155132 75880 155184 75886
rect 155132 75822 155184 75828
rect 155132 75608 155184 75614
rect 155132 75550 155184 75556
rect 155040 35284 155092 35290
rect 155040 35226 155092 35232
rect 155144 35222 155172 75550
rect 155236 75138 155264 77522
rect 155314 77480 155370 77489
rect 155314 77415 155370 77424
rect 155328 76838 155356 77415
rect 155316 76832 155368 76838
rect 155316 76774 155368 76780
rect 155316 76696 155368 76702
rect 155316 76638 155368 76644
rect 155224 75132 155276 75138
rect 155224 75074 155276 75080
rect 155224 74996 155276 75002
rect 155224 74938 155276 74944
rect 155236 74866 155264 74938
rect 155224 74860 155276 74866
rect 155224 74802 155276 74808
rect 155224 74724 155276 74730
rect 155224 74666 155276 74672
rect 155236 57390 155264 74666
rect 155328 62898 155356 76638
rect 155420 71874 155448 77658
rect 155512 72554 155540 77744
rect 155592 77648 155644 77654
rect 155592 77590 155644 77596
rect 155604 77294 155632 77590
rect 155604 77266 155724 77294
rect 155696 76809 155724 77266
rect 155682 76800 155738 76809
rect 155682 76735 155738 76744
rect 155684 76696 155736 76702
rect 155684 76638 155736 76644
rect 155592 76016 155644 76022
rect 155592 75958 155644 75964
rect 155604 73778 155632 75958
rect 155696 75478 155724 76638
rect 155788 75614 155816 77744
rect 156018 77772 156046 78132
rect 156110 77926 156138 78132
rect 156202 77931 156230 78132
rect 156098 77920 156150 77926
rect 156098 77862 156150 77868
rect 156188 77922 156244 77931
rect 156188 77857 156244 77866
rect 156294 77772 156322 78132
rect 156386 77926 156414 78132
rect 156478 77926 156506 78132
rect 156570 77926 156598 78132
rect 156374 77920 156426 77926
rect 156374 77862 156426 77868
rect 156466 77920 156518 77926
rect 156466 77862 156518 77868
rect 156558 77920 156610 77926
rect 156558 77862 156610 77868
rect 156018 77744 156092 77772
rect 155868 77726 155920 77732
rect 155776 75608 155828 75614
rect 155776 75550 155828 75556
rect 155684 75472 155736 75478
rect 155684 75414 155736 75420
rect 155592 73772 155644 73778
rect 155592 73714 155644 73720
rect 155880 73154 155908 77726
rect 155958 77616 156014 77625
rect 155958 77551 156014 77560
rect 155972 75970 156000 77551
rect 156064 76294 156092 77744
rect 156156 77744 156322 77772
rect 156420 77784 156472 77790
rect 156156 76702 156184 77744
rect 156662 77772 156690 78132
rect 156754 77926 156782 78132
rect 156846 77926 156874 78132
rect 156742 77920 156794 77926
rect 156742 77862 156794 77868
rect 156834 77920 156886 77926
rect 156834 77862 156886 77868
rect 156788 77784 156840 77790
rect 156662 77744 156736 77772
rect 156420 77726 156472 77732
rect 156236 77648 156288 77654
rect 156236 77590 156288 77596
rect 156144 76696 156196 76702
rect 156144 76638 156196 76644
rect 156144 76560 156196 76566
rect 156144 76502 156196 76508
rect 156052 76288 156104 76294
rect 156052 76230 156104 76236
rect 155972 75942 156092 75970
rect 155960 75880 156012 75886
rect 156064 75857 156092 75942
rect 155960 75822 156012 75828
rect 156050 75848 156106 75857
rect 155788 73126 155908 73154
rect 155788 72865 155816 73126
rect 155774 72856 155830 72865
rect 155774 72791 155830 72800
rect 155500 72548 155552 72554
rect 155500 72490 155552 72496
rect 155408 71868 155460 71874
rect 155408 71810 155460 71816
rect 155316 62892 155368 62898
rect 155316 62834 155368 62840
rect 155224 57384 155276 57390
rect 155224 57326 155276 57332
rect 155132 35216 155184 35222
rect 155132 35158 155184 35164
rect 154948 31340 155000 31346
rect 154948 31282 155000 31288
rect 154856 29708 154908 29714
rect 154856 29650 154908 29656
rect 154764 16108 154816 16114
rect 154764 16050 154816 16056
rect 154672 14612 154724 14618
rect 154672 14554 154724 14560
rect 154580 13388 154632 13394
rect 154580 13330 154632 13336
rect 153568 11892 153620 11898
rect 153568 11834 153620 11840
rect 153476 11824 153528 11830
rect 153476 11766 153528 11772
rect 153384 11756 153436 11762
rect 153384 11698 153436 11704
rect 153292 9104 153344 9110
rect 153292 9046 153344 9052
rect 155972 6458 156000 75822
rect 156050 75783 156106 75792
rect 156050 75712 156106 75721
rect 156050 75647 156106 75656
rect 155960 6452 156012 6458
rect 155960 6394 156012 6400
rect 156064 6390 156092 75647
rect 156156 13258 156184 76502
rect 156248 13326 156276 77590
rect 156326 77072 156382 77081
rect 156326 77007 156382 77016
rect 156340 75886 156368 77007
rect 156432 76430 156460 77726
rect 156512 77648 156564 77654
rect 156708 77625 156736 77744
rect 156788 77726 156840 77732
rect 156512 77590 156564 77596
rect 156694 77616 156750 77625
rect 156420 76424 156472 76430
rect 156420 76366 156472 76372
rect 156420 76288 156472 76294
rect 156420 76230 156472 76236
rect 156328 75880 156380 75886
rect 156328 75822 156380 75828
rect 156432 75698 156460 76230
rect 156340 75670 156460 75698
rect 156340 14482 156368 75670
rect 156420 75472 156472 75478
rect 156420 75414 156472 75420
rect 156432 16046 156460 75414
rect 156524 50522 156552 77590
rect 156604 77580 156656 77586
rect 156694 77551 156750 77560
rect 156604 77522 156656 77528
rect 156616 75562 156644 77522
rect 156696 77308 156748 77314
rect 156696 77250 156748 77256
rect 156708 75886 156736 77250
rect 156800 76566 156828 77726
rect 156938 77704 156966 78132
rect 157030 77772 157058 78132
rect 157122 77931 157150 78132
rect 157108 77922 157164 77931
rect 157108 77857 157164 77866
rect 157214 77772 157242 78132
rect 157306 77926 157334 78132
rect 157294 77920 157346 77926
rect 157398 77897 157426 78132
rect 157490 77926 157518 78132
rect 157582 77926 157610 78132
rect 157674 77926 157702 78132
rect 157766 77931 157794 78132
rect 157478 77920 157530 77926
rect 157294 77862 157346 77868
rect 157384 77888 157440 77897
rect 157478 77862 157530 77868
rect 157570 77920 157622 77926
rect 157570 77862 157622 77868
rect 157662 77920 157714 77926
rect 157662 77862 157714 77868
rect 157752 77922 157808 77931
rect 157858 77926 157886 78132
rect 157950 77926 157978 78132
rect 157752 77857 157808 77866
rect 157846 77920 157898 77926
rect 157846 77862 157898 77868
rect 157938 77920 157990 77926
rect 157938 77862 157990 77868
rect 157384 77823 157440 77832
rect 157524 77784 157576 77790
rect 157030 77744 157104 77772
rect 157214 77761 157288 77772
rect 157214 77752 157302 77761
rect 157214 77744 157246 77752
rect 156938 77676 157012 77704
rect 156984 77586 157012 77676
rect 156880 77580 156932 77586
rect 156880 77522 156932 77528
rect 156972 77580 157024 77586
rect 156972 77522 157024 77528
rect 156788 76560 156840 76566
rect 156788 76502 156840 76508
rect 156788 76424 156840 76430
rect 156788 76366 156840 76372
rect 156696 75880 156748 75886
rect 156696 75822 156748 75828
rect 156616 75534 156736 75562
rect 156604 75472 156656 75478
rect 156604 75414 156656 75420
rect 156616 54534 156644 75414
rect 156708 75206 156736 75534
rect 156696 75200 156748 75206
rect 156696 75142 156748 75148
rect 156800 71774 156828 76366
rect 156892 75478 156920 77522
rect 156972 77444 157024 77450
rect 156972 77386 157024 77392
rect 156880 75472 156932 75478
rect 156880 75414 156932 75420
rect 156984 73154 157012 77386
rect 157076 75449 157104 77744
rect 157430 77752 157486 77761
rect 157246 77687 157302 77696
rect 157340 77716 157392 77722
rect 157708 77784 157760 77790
rect 157524 77726 157576 77732
rect 157628 77732 157708 77738
rect 158042 77772 158070 78132
rect 157628 77726 157760 77732
rect 157890 77752 157946 77761
rect 157430 77687 157486 77696
rect 157340 77658 157392 77664
rect 157156 77648 157208 77654
rect 157156 77590 157208 77596
rect 157168 75954 157196 77590
rect 157248 77580 157300 77586
rect 157248 77522 157300 77528
rect 157156 75948 157208 75954
rect 157156 75890 157208 75896
rect 157260 75698 157288 77522
rect 157352 75914 157380 77658
rect 157444 76022 157472 77687
rect 157536 76702 157564 77726
rect 157628 77710 157748 77726
rect 157524 76696 157576 76702
rect 157524 76638 157576 76644
rect 157432 76016 157484 76022
rect 157432 75958 157484 75964
rect 157524 75948 157576 75954
rect 157352 75886 157472 75914
rect 157524 75890 157576 75896
rect 157444 75721 157472 75886
rect 157168 75670 157288 75698
rect 157430 75712 157486 75721
rect 157062 75440 157118 75449
rect 157062 75375 157118 75384
rect 156708 71746 156828 71774
rect 156892 73126 157012 73154
rect 156892 71774 156920 73126
rect 157168 72729 157196 75670
rect 157430 75647 157486 75656
rect 157340 75608 157392 75614
rect 157340 75550 157392 75556
rect 157248 75132 157300 75138
rect 157248 75074 157300 75080
rect 157260 73642 157288 75074
rect 157248 73636 157300 73642
rect 157248 73578 157300 73584
rect 157154 72720 157210 72729
rect 157154 72655 157210 72664
rect 156892 71746 157196 71774
rect 156708 67114 156736 71746
rect 157168 70394 157196 71746
rect 156800 70366 157196 70394
rect 156800 69698 156828 70366
rect 156788 69692 156840 69698
rect 156788 69634 156840 69640
rect 156696 67108 156748 67114
rect 156696 67050 156748 67056
rect 156604 54528 156656 54534
rect 156604 54470 156656 54476
rect 156512 50516 156564 50522
rect 156512 50458 156564 50464
rect 156420 16040 156472 16046
rect 156420 15982 156472 15988
rect 156328 14476 156380 14482
rect 156328 14418 156380 14424
rect 156236 13320 156288 13326
rect 156236 13262 156288 13268
rect 156144 13252 156196 13258
rect 156144 13194 156196 13200
rect 156052 6384 156104 6390
rect 156052 6326 156104 6332
rect 153200 5160 153252 5166
rect 153200 5102 153252 5108
rect 157352 5098 157380 75550
rect 157432 75540 157484 75546
rect 157432 75482 157484 75488
rect 157444 9042 157472 75482
rect 157536 13190 157564 75890
rect 157628 75342 157656 77710
rect 157890 77687 157946 77696
rect 157996 77744 158070 77772
rect 158134 77772 158162 78132
rect 158226 77926 158254 78132
rect 158318 77926 158346 78132
rect 158214 77920 158266 77926
rect 158214 77862 158266 77868
rect 158306 77920 158358 77926
rect 158306 77862 158358 77868
rect 158410 77772 158438 78132
rect 158502 77897 158530 78132
rect 158488 77888 158544 77897
rect 158488 77823 158544 77832
rect 158594 77772 158622 78132
rect 158686 77897 158714 78132
rect 158672 77888 158728 77897
rect 158672 77823 158728 77832
rect 158778 77772 158806 78132
rect 158870 77926 158898 78132
rect 158962 77926 158990 78132
rect 159054 77926 159082 78132
rect 159146 77926 159174 78132
rect 158858 77920 158910 77926
rect 158858 77862 158910 77868
rect 158950 77920 159002 77926
rect 158950 77862 159002 77868
rect 159042 77920 159094 77926
rect 159042 77862 159094 77868
rect 159134 77920 159186 77926
rect 159134 77862 159186 77868
rect 158134 77744 158208 77772
rect 158410 77744 158484 77772
rect 158548 77761 158622 77772
rect 157708 77648 157760 77654
rect 157708 77590 157760 77596
rect 157800 77648 157852 77654
rect 157800 77590 157852 77596
rect 157616 75336 157668 75342
rect 157616 75278 157668 75284
rect 157616 75200 157668 75206
rect 157616 75142 157668 75148
rect 157628 15978 157656 75142
rect 157720 23118 157748 77590
rect 157812 60042 157840 77590
rect 157904 75614 157932 77687
rect 157892 75608 157944 75614
rect 157892 75550 157944 75556
rect 157996 75546 158024 77744
rect 158076 77512 158128 77518
rect 158076 77454 158128 77460
rect 157984 75540 158036 75546
rect 157984 75482 158036 75488
rect 157892 75336 157944 75342
rect 157892 75278 157944 75284
rect 157904 62830 157932 75278
rect 158088 75206 158116 77454
rect 158180 77294 158208 77744
rect 158260 77716 158312 77722
rect 158260 77658 158312 77664
rect 158272 77625 158300 77658
rect 158258 77616 158314 77625
rect 158456 77602 158484 77744
rect 158534 77752 158622 77761
rect 158590 77744 158622 77752
rect 158732 77744 158806 77772
rect 159238 77761 159266 78132
rect 159330 77858 159358 78132
rect 159422 77858 159450 78132
rect 159318 77852 159370 77858
rect 159318 77794 159370 77800
rect 159410 77852 159462 77858
rect 159410 77794 159462 77800
rect 159224 77752 159280 77761
rect 158534 77687 158590 77696
rect 158732 77602 158760 77744
rect 159224 77687 159280 77696
rect 158258 77551 158314 77560
rect 158364 77574 158484 77602
rect 158640 77574 158760 77602
rect 158812 77648 158864 77654
rect 158812 77590 158864 77596
rect 158996 77648 159048 77654
rect 158996 77590 159048 77596
rect 159088 77648 159140 77654
rect 159514 77602 159542 78132
rect 159606 77926 159634 78132
rect 159594 77920 159646 77926
rect 159594 77862 159646 77868
rect 159698 77772 159726 78132
rect 159790 77926 159818 78132
rect 159882 77926 159910 78132
rect 159974 77926 160002 78132
rect 160066 77926 160094 78132
rect 160158 77926 160186 78132
rect 159778 77920 159830 77926
rect 159778 77862 159830 77868
rect 159870 77920 159922 77926
rect 159870 77862 159922 77868
rect 159962 77920 160014 77926
rect 159962 77862 160014 77868
rect 160054 77920 160106 77926
rect 160054 77862 160106 77868
rect 160146 77920 160198 77926
rect 160146 77862 160198 77868
rect 159698 77761 159772 77772
rect 159698 77752 159786 77761
rect 159698 77744 159730 77752
rect 160250 77738 160278 78132
rect 160342 77926 160370 78132
rect 160330 77920 160382 77926
rect 160330 77862 160382 77868
rect 159730 77687 159786 77696
rect 160204 77710 160278 77738
rect 159088 77590 159140 77596
rect 158180 77266 158300 77294
rect 158076 75200 158128 75206
rect 158076 75142 158128 75148
rect 158272 75070 158300 77266
rect 158364 76129 158392 77574
rect 158444 77512 158496 77518
rect 158496 77472 158576 77500
rect 158444 77454 158496 77460
rect 158444 77308 158496 77314
rect 158444 77250 158496 77256
rect 158350 76120 158406 76129
rect 158350 76055 158406 76064
rect 158352 76016 158404 76022
rect 158352 75958 158404 75964
rect 158260 75064 158312 75070
rect 158260 75006 158312 75012
rect 158364 73154 158392 75958
rect 158456 75614 158484 77250
rect 158548 77081 158576 77472
rect 158534 77072 158590 77081
rect 158534 77007 158590 77016
rect 158640 76770 158668 77574
rect 158628 76764 158680 76770
rect 158628 76706 158680 76712
rect 158720 76696 158772 76702
rect 158720 76638 158772 76644
rect 158536 76152 158588 76158
rect 158536 76094 158588 76100
rect 158444 75608 158496 75614
rect 158444 75550 158496 75556
rect 158548 75410 158576 76094
rect 158732 75546 158760 76638
rect 158720 75540 158772 75546
rect 158720 75482 158772 75488
rect 158536 75404 158588 75410
rect 158536 75346 158588 75352
rect 158824 74984 158852 77590
rect 158904 77580 158956 77586
rect 158904 77522 158956 77528
rect 158916 75177 158944 77522
rect 158902 75168 158958 75177
rect 158902 75103 158958 75112
rect 157996 73126 158392 73154
rect 158732 74956 158852 74984
rect 158904 74996 158956 75002
rect 157996 65754 158024 73126
rect 158352 72684 158404 72690
rect 158352 72626 158404 72632
rect 157984 65748 158036 65754
rect 157984 65690 158036 65696
rect 157892 62824 157944 62830
rect 157892 62766 157944 62772
rect 157800 60036 157852 60042
rect 157800 59978 157852 59984
rect 157708 23112 157760 23118
rect 157708 23054 157760 23060
rect 158364 21826 158392 72626
rect 158352 21820 158404 21826
rect 158352 21762 158404 21768
rect 157616 15972 157668 15978
rect 157616 15914 157668 15920
rect 157524 13184 157576 13190
rect 157524 13126 157576 13132
rect 158732 10470 158760 74956
rect 158904 74938 158956 74944
rect 158812 74792 158864 74798
rect 158812 74734 158864 74740
rect 158824 17542 158852 74734
rect 158916 17610 158944 74938
rect 159008 21690 159036 77590
rect 159100 73914 159128 77590
rect 159180 77580 159232 77586
rect 159180 77522 159232 77528
rect 159468 77574 159542 77602
rect 159640 77648 159692 77654
rect 159640 77590 159692 77596
rect 159916 77648 159968 77654
rect 159916 77590 159968 77596
rect 160008 77648 160060 77654
rect 160008 77590 160060 77596
rect 160100 77648 160152 77654
rect 160100 77590 160152 77596
rect 159192 76090 159220 77522
rect 159272 77512 159324 77518
rect 159272 77454 159324 77460
rect 159180 76084 159232 76090
rect 159180 76026 159232 76032
rect 159180 75948 159232 75954
rect 159180 75890 159232 75896
rect 159088 73908 159140 73914
rect 159088 73850 159140 73856
rect 159088 72004 159140 72010
rect 159088 71946 159140 71952
rect 158996 21684 159048 21690
rect 158996 21626 159048 21632
rect 159100 21622 159128 71946
rect 159192 31278 159220 75890
rect 159284 75002 159312 77454
rect 159364 77376 159416 77382
rect 159364 77318 159416 77324
rect 159376 75954 159404 77318
rect 159364 75948 159416 75954
rect 159364 75890 159416 75896
rect 159364 75608 159416 75614
rect 159364 75550 159416 75556
rect 159272 74996 159324 75002
rect 159272 74938 159324 74944
rect 159272 73908 159324 73914
rect 159272 73850 159324 73856
rect 159284 61538 159312 73850
rect 159376 64190 159404 75550
rect 159468 72010 159496 77574
rect 159546 77480 159602 77489
rect 159546 77415 159602 77424
rect 159560 77081 159588 77415
rect 159546 77072 159602 77081
rect 159546 77007 159602 77016
rect 159548 76220 159600 76226
rect 159548 76162 159600 76168
rect 159560 74798 159588 76162
rect 159548 74792 159600 74798
rect 159548 74734 159600 74740
rect 159652 74633 159680 77590
rect 159928 76226 159956 77590
rect 159916 76220 159968 76226
rect 159916 76162 159968 76168
rect 159916 76084 159968 76090
rect 159916 76026 159968 76032
rect 159638 74624 159694 74633
rect 159638 74559 159694 74568
rect 159928 72758 159956 76026
rect 160020 75041 160048 77590
rect 160112 76566 160140 77590
rect 160100 76560 160152 76566
rect 160100 76502 160152 76508
rect 160100 76084 160152 76090
rect 160100 76026 160152 76032
rect 160006 75032 160062 75041
rect 160006 74967 160062 74976
rect 160112 74934 160140 76026
rect 160100 74928 160152 74934
rect 160100 74870 160152 74876
rect 160204 74780 160232 77710
rect 160434 77704 160462 78132
rect 160526 77926 160554 78132
rect 160514 77920 160566 77926
rect 160514 77862 160566 77868
rect 160618 77858 160646 78132
rect 160606 77852 160658 77858
rect 160606 77794 160658 77800
rect 160710 77761 160738 78132
rect 160802 77772 160830 78132
rect 160894 77926 160922 78132
rect 160986 77926 161014 78132
rect 160882 77920 160934 77926
rect 160882 77862 160934 77868
rect 160974 77920 161026 77926
rect 160974 77862 161026 77868
rect 160388 77676 160462 77704
rect 160696 77752 160752 77761
rect 160802 77744 160876 77772
rect 160696 77687 160752 77696
rect 160284 77580 160336 77586
rect 160284 77522 160336 77528
rect 160296 75614 160324 77522
rect 160284 75608 160336 75614
rect 160284 75550 160336 75556
rect 160284 75472 160336 75478
rect 160284 75414 160336 75420
rect 160112 74752 160232 74780
rect 159916 72752 159968 72758
rect 159916 72694 159968 72700
rect 159456 72004 159508 72010
rect 159456 71946 159508 71952
rect 159364 64184 159416 64190
rect 159364 64126 159416 64132
rect 159272 61532 159324 61538
rect 159272 61474 159324 61480
rect 159180 31272 159232 31278
rect 159180 31214 159232 31220
rect 159088 21616 159140 21622
rect 159088 21558 159140 21564
rect 158904 17604 158956 17610
rect 158904 17546 158956 17552
rect 158812 17536 158864 17542
rect 158812 17478 158864 17484
rect 158902 16416 158958 16425
rect 158902 16351 158958 16360
rect 158720 10464 158772 10470
rect 158720 10406 158772 10412
rect 157432 9036 157484 9042
rect 157432 8978 157484 8984
rect 157340 5092 157392 5098
rect 157340 5034 157392 5040
rect 154212 4956 154264 4962
rect 154212 4898 154264 4904
rect 153016 3936 153068 3942
rect 153016 3878 153068 3884
rect 152832 3188 152884 3194
rect 152832 3130 152884 3136
rect 153028 480 153056 3878
rect 154224 480 154252 4898
rect 157800 4888 157852 4894
rect 157800 4830 157852 4836
rect 155408 3800 155460 3806
rect 155408 3742 155460 3748
rect 155420 480 155448 3742
rect 156604 3188 156656 3194
rect 156604 3130 156656 3136
rect 156616 480 156644 3130
rect 157812 480 157840 4830
rect 158916 480 158944 16351
rect 160112 6322 160140 74752
rect 160192 74044 160244 74050
rect 160192 73986 160244 73992
rect 160204 17338 160232 73986
rect 160296 17474 160324 75414
rect 160388 75206 160416 77676
rect 160560 77648 160612 77654
rect 160466 77616 160522 77625
rect 160560 77590 160612 77596
rect 160744 77648 160796 77654
rect 160744 77590 160796 77596
rect 160466 77551 160522 77560
rect 160480 76158 160508 77551
rect 160468 76152 160520 76158
rect 160468 76094 160520 76100
rect 160468 75608 160520 75614
rect 160468 75550 160520 75556
rect 160376 75200 160428 75206
rect 160376 75142 160428 75148
rect 160376 74792 160428 74798
rect 160480 74780 160508 75550
rect 160572 75478 160600 77590
rect 160652 77580 160704 77586
rect 160652 77522 160704 77528
rect 160664 75614 160692 77522
rect 160652 75608 160704 75614
rect 160756 75585 160784 77590
rect 160652 75550 160704 75556
rect 160742 75576 160798 75585
rect 160742 75511 160798 75520
rect 160560 75472 160612 75478
rect 160560 75414 160612 75420
rect 160560 75336 160612 75342
rect 160560 75278 160612 75284
rect 160572 74934 160600 75278
rect 160652 75200 160704 75206
rect 160652 75142 160704 75148
rect 160560 74928 160612 74934
rect 160560 74870 160612 74876
rect 160480 74752 160600 74780
rect 160376 74734 160428 74740
rect 160284 17468 160336 17474
rect 160284 17410 160336 17416
rect 160192 17332 160244 17338
rect 160192 17274 160244 17280
rect 160388 17270 160416 74734
rect 160466 74488 160522 74497
rect 160466 74423 160522 74432
rect 160480 17406 160508 74423
rect 160572 26994 160600 74752
rect 160664 58750 160692 75142
rect 160848 74050 160876 77744
rect 161078 77738 161106 78132
rect 161032 77727 161106 77738
rect 160928 77716 160980 77722
rect 160928 77658 160980 77664
rect 161018 77718 161106 77727
rect 161074 77710 161106 77718
rect 160940 74644 160968 77658
rect 161018 77653 161074 77662
rect 161170 77636 161198 78132
rect 161262 77858 161290 78132
rect 161354 77858 161382 78132
rect 161446 77858 161474 78132
rect 161250 77852 161302 77858
rect 161250 77794 161302 77800
rect 161342 77852 161394 77858
rect 161342 77794 161394 77800
rect 161434 77852 161486 77858
rect 161434 77794 161486 77800
rect 161538 77772 161566 78132
rect 161630 77926 161658 78132
rect 161722 77926 161750 78132
rect 161814 77926 161842 78132
rect 161618 77920 161670 77926
rect 161618 77862 161670 77868
rect 161710 77920 161762 77926
rect 161710 77862 161762 77868
rect 161802 77920 161854 77926
rect 161802 77862 161854 77868
rect 161538 77744 161612 77772
rect 161296 77716 161348 77722
rect 161296 77658 161348 77664
rect 161388 77716 161440 77722
rect 161388 77658 161440 77664
rect 161124 77608 161198 77636
rect 161020 77580 161072 77586
rect 161020 77522 161072 77528
rect 161032 74798 161060 77522
rect 161124 75206 161152 77608
rect 161204 77512 161256 77518
rect 161204 77454 161256 77460
rect 161216 76634 161244 77454
rect 161204 76628 161256 76634
rect 161204 76570 161256 76576
rect 161308 75585 161336 77658
rect 161400 75993 161428 77658
rect 161478 77616 161534 77625
rect 161478 77551 161534 77560
rect 161386 75984 161442 75993
rect 161386 75919 161442 75928
rect 161294 75576 161350 75585
rect 161294 75511 161350 75520
rect 161296 75472 161348 75478
rect 161296 75414 161348 75420
rect 161112 75200 161164 75206
rect 161112 75142 161164 75148
rect 161020 74792 161072 74798
rect 161020 74734 161072 74740
rect 160940 74616 161244 74644
rect 160836 74044 160888 74050
rect 160836 73986 160888 73992
rect 161020 73500 161072 73506
rect 161020 73442 161072 73448
rect 161032 63034 161060 73442
rect 161216 72622 161244 74616
rect 161308 73506 161336 75414
rect 161388 74928 161440 74934
rect 161388 74870 161440 74876
rect 161296 73500 161348 73506
rect 161296 73442 161348 73448
rect 161204 72616 161256 72622
rect 161204 72558 161256 72564
rect 161400 71126 161428 74870
rect 161388 71120 161440 71126
rect 161388 71062 161440 71068
rect 161020 63028 161072 63034
rect 161020 62970 161072 62976
rect 160652 58744 160704 58750
rect 160652 58686 160704 58692
rect 160560 26988 160612 26994
rect 160560 26930 160612 26936
rect 160468 17400 160520 17406
rect 160468 17342 160520 17348
rect 160376 17264 160428 17270
rect 160376 17206 160428 17212
rect 161492 7614 161520 77551
rect 161584 77314 161612 77744
rect 161906 77704 161934 78132
rect 161998 77926 162026 78132
rect 161986 77920 162038 77926
rect 161986 77862 162038 77868
rect 162090 77858 162118 78132
rect 162182 77926 162210 78132
rect 162170 77920 162222 77926
rect 162170 77862 162222 77868
rect 162078 77852 162130 77858
rect 162078 77794 162130 77800
rect 162274 77772 162302 78132
rect 162366 77897 162394 78132
rect 162458 77926 162486 78132
rect 162446 77920 162498 77926
rect 162352 77888 162408 77897
rect 162446 77862 162498 77868
rect 162352 77823 162408 77832
rect 162550 77772 162578 78132
rect 162642 77926 162670 78132
rect 162734 77931 162762 78132
rect 162630 77920 162682 77926
rect 162630 77862 162682 77868
rect 162720 77922 162776 77931
rect 162826 77926 162854 78132
rect 162918 77926 162946 78132
rect 163010 77926 163038 78132
rect 162720 77857 162776 77866
rect 162814 77920 162866 77926
rect 162814 77862 162866 77868
rect 162906 77920 162958 77926
rect 162906 77862 162958 77868
rect 162998 77920 163050 77926
rect 163102 77897 163130 78132
rect 162998 77862 163050 77868
rect 163088 77888 163144 77897
rect 163088 77823 163144 77832
rect 162274 77744 162440 77772
rect 162550 77761 162624 77772
rect 162550 77752 162638 77761
rect 162550 77744 162582 77752
rect 162412 77738 162440 77744
rect 161860 77676 161934 77704
rect 162032 77716 162084 77722
rect 161756 77580 161808 77586
rect 161756 77522 161808 77528
rect 161664 77512 161716 77518
rect 161664 77454 161716 77460
rect 161572 77308 161624 77314
rect 161572 77250 161624 77256
rect 161572 76356 161624 76362
rect 161572 76298 161624 76304
rect 161584 76022 161612 76298
rect 161572 76016 161624 76022
rect 161572 75958 161624 75964
rect 161676 75914 161704 77454
rect 161768 76129 161796 77522
rect 161754 76120 161810 76129
rect 161754 76055 161810 76064
rect 161756 76016 161808 76022
rect 161756 75958 161808 75964
rect 161584 75886 161704 75914
rect 161584 18834 161612 75886
rect 161664 75336 161716 75342
rect 161664 75278 161716 75284
rect 161676 26926 161704 75278
rect 161768 28354 161796 75958
rect 161860 29646 161888 77676
rect 162032 77658 162084 77664
rect 162124 77716 162176 77722
rect 162412 77710 162486 77738
rect 162124 77658 162176 77664
rect 161940 77580 161992 77586
rect 161940 77522 161992 77528
rect 161952 76362 161980 77522
rect 161940 76356 161992 76362
rect 161940 76298 161992 76304
rect 161940 76220 161992 76226
rect 161940 76162 161992 76168
rect 161952 75886 161980 76162
rect 161940 75880 161992 75886
rect 161940 75822 161992 75828
rect 161940 75404 161992 75410
rect 161940 75346 161992 75352
rect 161952 73710 161980 75346
rect 161940 73704 161992 73710
rect 161940 73646 161992 73652
rect 162044 64874 162072 77658
rect 162136 76106 162164 77658
rect 162308 77648 162360 77654
rect 162458 77602 162486 77710
rect 162582 77687 162638 77696
rect 162308 77590 162360 77596
rect 162216 77444 162268 77450
rect 162216 77386 162268 77392
rect 162228 76702 162256 77386
rect 162216 76696 162268 76702
rect 162216 76638 162268 76644
rect 162136 76078 162256 76106
rect 162124 75948 162176 75954
rect 162124 75890 162176 75896
rect 162136 74866 162164 75890
rect 162228 75342 162256 76078
rect 162320 75426 162348 77590
rect 162412 77574 162486 77602
rect 162860 77648 162912 77654
rect 163194 77636 163222 78132
rect 163286 77772 163314 78132
rect 163378 77926 163406 78132
rect 163366 77920 163418 77926
rect 163470 77897 163498 78132
rect 163562 77926 163590 78132
rect 163654 77926 163682 78132
rect 163746 77926 163774 78132
rect 163838 77926 163866 78132
rect 163930 77926 163958 78132
rect 164022 77931 164050 78132
rect 163550 77920 163602 77926
rect 163366 77862 163418 77868
rect 163456 77888 163512 77897
rect 163550 77862 163602 77868
rect 163642 77920 163694 77926
rect 163642 77862 163694 77868
rect 163734 77920 163786 77926
rect 163734 77862 163786 77868
rect 163826 77920 163878 77926
rect 163826 77862 163878 77868
rect 163918 77920 163970 77926
rect 163918 77862 163970 77868
rect 164008 77922 164064 77931
rect 164008 77857 164064 77866
rect 163456 77823 163512 77832
rect 163412 77784 163464 77790
rect 163286 77744 163360 77772
rect 162860 77590 162912 77596
rect 163148 77608 163222 77636
rect 162768 77580 162820 77586
rect 162412 75546 162440 77574
rect 162768 77522 162820 77528
rect 162492 77512 162544 77518
rect 162492 77454 162544 77460
rect 162504 76265 162532 77454
rect 162584 77444 162636 77450
rect 162584 77386 162636 77392
rect 162596 76401 162624 77386
rect 162676 76832 162728 76838
rect 162674 76800 162676 76809
rect 162728 76800 162730 76809
rect 162674 76735 162730 76744
rect 162582 76392 162638 76401
rect 162582 76327 162638 76336
rect 162490 76256 162546 76265
rect 162490 76191 162546 76200
rect 162400 75540 162452 75546
rect 162400 75482 162452 75488
rect 162320 75398 162716 75426
rect 162216 75336 162268 75342
rect 162216 75278 162268 75284
rect 162400 75268 162452 75274
rect 162400 75210 162452 75216
rect 162124 74860 162176 74866
rect 162124 74802 162176 74808
rect 162412 73828 162440 75210
rect 161952 64846 162072 64874
rect 162228 73800 162440 73828
rect 161952 50454 161980 64846
rect 162228 64258 162256 73800
rect 162308 73704 162360 73710
rect 162308 73646 162360 73652
rect 162216 64252 162268 64258
rect 162216 64194 162268 64200
rect 162320 58818 162348 73646
rect 162688 72826 162716 75398
rect 162780 75274 162808 77522
rect 162768 75268 162820 75274
rect 162768 75210 162820 75216
rect 162872 74866 162900 77590
rect 162952 77512 163004 77518
rect 162950 77480 162952 77489
rect 163004 77480 163006 77489
rect 162950 77415 163006 77424
rect 162952 77240 163004 77246
rect 162952 77182 163004 77188
rect 163042 77208 163098 77217
rect 162964 76362 162992 77182
rect 163042 77143 163098 77152
rect 163056 76430 163084 77143
rect 163044 76424 163096 76430
rect 163044 76366 163096 76372
rect 162952 76356 163004 76362
rect 162952 76298 163004 76304
rect 162952 75472 163004 75478
rect 162952 75414 163004 75420
rect 162860 74860 162912 74866
rect 162860 74802 162912 74808
rect 162860 74656 162912 74662
rect 162860 74598 162912 74604
rect 162676 72820 162728 72826
rect 162676 72762 162728 72768
rect 162308 58812 162360 58818
rect 162308 58754 162360 58760
rect 161940 50448 161992 50454
rect 161940 50390 161992 50396
rect 161848 29640 161900 29646
rect 161848 29582 161900 29588
rect 161756 28348 161808 28354
rect 161756 28290 161808 28296
rect 161664 26920 161716 26926
rect 161664 26862 161716 26868
rect 161572 18828 161624 18834
rect 161572 18770 161624 18776
rect 161480 7608 161532 7614
rect 161480 7550 161532 7556
rect 160100 6316 160152 6322
rect 160100 6258 160152 6264
rect 162872 4962 162900 74598
rect 162964 6254 162992 75414
rect 163148 75342 163176 77608
rect 163332 77294 163360 77744
rect 163412 77726 163464 77732
rect 163964 77784 164016 77790
rect 164114 77772 164142 78132
rect 164206 77897 164234 78132
rect 164298 77926 164326 78132
rect 164286 77920 164338 77926
rect 164192 77888 164248 77897
rect 164286 77862 164338 77868
rect 164192 77823 164248 77832
rect 163964 77726 164016 77732
rect 164068 77744 164142 77772
rect 164390 77772 164418 78132
rect 164482 77926 164510 78132
rect 164574 77926 164602 78132
rect 164470 77920 164522 77926
rect 164470 77862 164522 77868
rect 164562 77920 164614 77926
rect 164562 77862 164614 77868
rect 164390 77744 164464 77772
rect 163240 77266 163360 77294
rect 163136 75336 163188 75342
rect 163136 75278 163188 75284
rect 163240 75188 163268 77266
rect 163424 76072 163452 77726
rect 163688 77716 163740 77722
rect 163688 77658 163740 77664
rect 163780 77716 163832 77722
rect 163780 77658 163832 77664
rect 163504 77648 163556 77654
rect 163504 77590 163556 77596
rect 163148 75160 163268 75188
rect 163332 76044 163452 76072
rect 163044 73364 163096 73370
rect 163044 73306 163096 73312
rect 163056 8974 163084 73306
rect 163148 20126 163176 75160
rect 163228 74996 163280 75002
rect 163228 74938 163280 74944
rect 163136 20120 163188 20126
rect 163136 20062 163188 20068
rect 163240 20058 163268 74938
rect 163332 32570 163360 76044
rect 163410 75984 163466 75993
rect 163410 75919 163466 75928
rect 163424 50386 163452 75919
rect 163516 75002 163544 77590
rect 163596 77580 163648 77586
rect 163596 77522 163648 77528
rect 163608 77246 163636 77522
rect 163596 77240 163648 77246
rect 163596 77182 163648 77188
rect 163594 75576 163650 75585
rect 163594 75511 163650 75520
rect 163504 74996 163556 75002
rect 163504 74938 163556 74944
rect 163504 74860 163556 74866
rect 163504 74802 163556 74808
rect 163516 58682 163544 74802
rect 163608 68542 163636 75511
rect 163700 74662 163728 77658
rect 163688 74656 163740 74662
rect 163688 74598 163740 74604
rect 163792 73370 163820 77658
rect 163872 77648 163924 77654
rect 163872 77590 163924 77596
rect 163884 75818 163912 77590
rect 163872 75812 163924 75818
rect 163872 75754 163924 75760
rect 163976 75478 164004 77726
rect 164068 76265 164096 77744
rect 164332 77648 164384 77654
rect 164436 77625 164464 77744
rect 164516 77716 164568 77722
rect 164516 77658 164568 77664
rect 164332 77590 164384 77596
rect 164422 77616 164478 77625
rect 164148 77580 164200 77586
rect 164148 77522 164200 77528
rect 164054 76256 164110 76265
rect 164054 76191 164110 76200
rect 164056 75812 164108 75818
rect 164056 75754 164108 75760
rect 163964 75472 164016 75478
rect 163964 75414 164016 75420
rect 163964 75268 164016 75274
rect 163964 75210 164016 75216
rect 163780 73364 163832 73370
rect 163780 73306 163832 73312
rect 163870 73128 163926 73137
rect 163870 73063 163926 73072
rect 163884 72690 163912 73063
rect 163872 72684 163924 72690
rect 163872 72626 163924 72632
rect 163780 72344 163832 72350
rect 163780 72286 163832 72292
rect 163596 68536 163648 68542
rect 163596 68478 163648 68484
rect 163504 58676 163556 58682
rect 163504 58618 163556 58624
rect 163412 50380 163464 50386
rect 163412 50322 163464 50328
rect 163320 32564 163372 32570
rect 163320 32506 163372 32512
rect 163228 20052 163280 20058
rect 163228 19994 163280 20000
rect 163044 8968 163096 8974
rect 163044 8910 163096 8916
rect 162952 6248 163004 6254
rect 162952 6190 163004 6196
rect 162860 4956 162912 4962
rect 162860 4898 162912 4904
rect 160098 4856 160154 4865
rect 160098 4791 160154 4800
rect 162492 4820 162544 4826
rect 160112 480 160140 4791
rect 162492 4762 162544 4768
rect 161294 3360 161350 3369
rect 161294 3295 161350 3304
rect 161308 480 161336 3295
rect 162504 480 162532 4762
rect 163688 3732 163740 3738
rect 163688 3674 163740 3680
rect 163700 480 163728 3674
rect 163792 3534 163820 72286
rect 163976 71806 164004 75210
rect 164068 72554 164096 75754
rect 164160 75478 164188 77522
rect 164238 77480 164294 77489
rect 164238 77415 164294 77424
rect 164252 76498 164280 77415
rect 164344 76566 164372 77590
rect 164422 77551 164478 77560
rect 164424 77512 164476 77518
rect 164424 77454 164476 77460
rect 164332 76560 164384 76566
rect 164332 76502 164384 76508
rect 164240 76492 164292 76498
rect 164240 76434 164292 76440
rect 164436 75698 164464 77454
rect 164344 75670 164464 75698
rect 164528 75682 164556 77658
rect 164666 77636 164694 78132
rect 164758 77738 164786 78132
rect 164850 77931 164878 78132
rect 164836 77922 164892 77931
rect 164942 77926 164970 78132
rect 165034 77926 165062 78132
rect 165126 77926 165154 78132
rect 165218 77926 165246 78132
rect 164836 77857 164892 77866
rect 164930 77920 164982 77926
rect 164930 77862 164982 77868
rect 165022 77920 165074 77926
rect 165022 77862 165074 77868
rect 165114 77920 165166 77926
rect 165114 77862 165166 77868
rect 165206 77920 165258 77926
rect 165310 77897 165338 78132
rect 165206 77862 165258 77868
rect 165296 77888 165352 77897
rect 165296 77823 165352 77832
rect 164758 77710 164924 77738
rect 164666 77608 164832 77636
rect 164700 77512 164752 77518
rect 164700 77454 164752 77460
rect 164516 75676 164568 75682
rect 164148 75472 164200 75478
rect 164148 75414 164200 75420
rect 164240 75404 164292 75410
rect 164240 75346 164292 75352
rect 164056 72548 164108 72554
rect 164056 72490 164108 72496
rect 163964 71800 164016 71806
rect 163964 71742 164016 71748
rect 164252 10402 164280 75346
rect 164344 13122 164372 75670
rect 164516 75618 164568 75624
rect 164608 75472 164660 75478
rect 164608 75414 164660 75420
rect 164514 75304 164570 75313
rect 164514 75239 164570 75248
rect 164424 75132 164476 75138
rect 164424 75074 164476 75080
rect 164436 74866 164464 75074
rect 164424 74860 164476 74866
rect 164424 74802 164476 74808
rect 164424 74724 164476 74730
rect 164424 74666 164476 74672
rect 164436 15910 164464 74666
rect 164528 19990 164556 75239
rect 164620 25634 164648 75414
rect 164608 25628 164660 25634
rect 164608 25570 164660 25576
rect 164712 25566 164740 77454
rect 164804 75410 164832 77608
rect 164896 77586 164924 77710
rect 165068 77716 165120 77722
rect 165068 77658 165120 77664
rect 165160 77716 165212 77722
rect 165160 77658 165212 77664
rect 164884 77580 164936 77586
rect 164884 77522 164936 77528
rect 164976 77580 165028 77586
rect 164976 77522 165028 77528
rect 164882 77480 164938 77489
rect 164882 77415 164938 77424
rect 164896 75886 164924 77415
rect 164884 75880 164936 75886
rect 164884 75822 164936 75828
rect 164792 75404 164844 75410
rect 164792 75346 164844 75352
rect 164988 75290 165016 77522
rect 164804 75262 165016 75290
rect 164804 31210 164832 75262
rect 164974 75168 165030 75177
rect 164884 75132 164936 75138
rect 165080 75138 165108 77658
rect 164974 75103 165030 75112
rect 165068 75132 165120 75138
rect 164884 75074 164936 75080
rect 164896 57322 164924 75074
rect 164988 68406 165016 75103
rect 165068 75074 165120 75080
rect 165172 74730 165200 77658
rect 165252 77648 165304 77654
rect 165402 77636 165430 78132
rect 165494 77931 165522 78132
rect 165480 77922 165536 77931
rect 165480 77857 165536 77866
rect 165586 77858 165614 78132
rect 165574 77852 165626 77858
rect 165574 77794 165626 77800
rect 165678 77738 165706 78132
rect 165252 77590 165304 77596
rect 165356 77608 165430 77636
rect 165632 77710 165706 77738
rect 165264 74798 165292 77590
rect 165356 77081 165384 77608
rect 165436 77376 165488 77382
rect 165436 77318 165488 77324
rect 165342 77072 165398 77081
rect 165342 77007 165398 77016
rect 165344 76492 165396 76498
rect 165344 76434 165396 76440
rect 165252 74792 165304 74798
rect 165252 74734 165304 74740
rect 165160 74724 165212 74730
rect 165160 74666 165212 74672
rect 165356 72593 165384 76434
rect 165448 75410 165476 77318
rect 165528 76832 165580 76838
rect 165526 76800 165528 76809
rect 165580 76800 165582 76809
rect 165526 76735 165582 76744
rect 165528 75676 165580 75682
rect 165528 75618 165580 75624
rect 165436 75404 165488 75410
rect 165436 75346 165488 75352
rect 165342 72584 165398 72593
rect 165342 72519 165398 72528
rect 165540 68474 165568 75618
rect 165632 74662 165660 77710
rect 165770 77636 165798 78132
rect 165862 77897 165890 78132
rect 165954 77926 165982 78132
rect 165942 77920 165994 77926
rect 165848 77888 165904 77897
rect 165942 77862 165994 77868
rect 165848 77823 165904 77832
rect 165896 77784 165948 77790
rect 166046 77772 166074 78132
rect 166138 77926 166166 78132
rect 166230 77926 166258 78132
rect 166126 77920 166178 77926
rect 166126 77862 166178 77868
rect 166218 77920 166270 77926
rect 166218 77862 166270 77868
rect 166046 77744 166212 77772
rect 165896 77726 165948 77732
rect 165724 77608 165798 77636
rect 165908 77636 165936 77726
rect 166080 77648 166132 77654
rect 165908 77608 166028 77636
rect 165620 74656 165672 74662
rect 165620 74598 165672 74604
rect 165724 73710 165752 77608
rect 165894 77480 165950 77489
rect 165894 77415 165950 77424
rect 165804 77376 165856 77382
rect 165804 77318 165856 77324
rect 165816 76226 165844 77318
rect 165804 76220 165856 76226
rect 165804 76162 165856 76168
rect 165804 76016 165856 76022
rect 165804 75958 165856 75964
rect 165816 75750 165844 75958
rect 165804 75744 165856 75750
rect 165804 75686 165856 75692
rect 165804 74724 165856 74730
rect 165804 74666 165856 74672
rect 165712 73704 165764 73710
rect 165712 73646 165764 73652
rect 165620 73568 165672 73574
rect 165620 73510 165672 73516
rect 165710 73536 165766 73545
rect 165528 68468 165580 68474
rect 165528 68410 165580 68416
rect 164976 68400 165028 68406
rect 164976 68342 165028 68348
rect 164884 57316 164936 57322
rect 164884 57258 164936 57264
rect 164792 31204 164844 31210
rect 164792 31146 164844 31152
rect 164700 25560 164752 25566
rect 164700 25502 164752 25508
rect 165632 21418 165660 73510
rect 165710 73471 165766 73480
rect 165724 21554 165752 73471
rect 165712 21548 165764 21554
rect 165712 21490 165764 21496
rect 165816 21486 165844 74666
rect 165908 28286 165936 77415
rect 166000 31074 166028 77608
rect 166184 77625 166212 77744
rect 166322 77636 166350 78132
rect 166414 77772 166442 78132
rect 166506 77926 166534 78132
rect 166598 77926 166626 78132
rect 166690 77926 166718 78132
rect 166494 77920 166546 77926
rect 166494 77862 166546 77868
rect 166586 77920 166638 77926
rect 166586 77862 166638 77868
rect 166678 77920 166730 77926
rect 166678 77862 166730 77868
rect 166782 77772 166810 78132
rect 166414 77744 166488 77772
rect 166080 77590 166132 77596
rect 166170 77616 166226 77625
rect 166092 75177 166120 77590
rect 166170 77551 166226 77560
rect 166276 77608 166350 77636
rect 166078 75168 166134 75177
rect 166078 75103 166134 75112
rect 166276 74730 166304 77608
rect 166356 77512 166408 77518
rect 166460 77489 166488 77744
rect 166736 77744 166810 77772
rect 166874 77772 166902 78132
rect 166966 77897 166994 78132
rect 166952 77888 167008 77897
rect 166952 77823 167008 77832
rect 166874 77744 166948 77772
rect 166540 77716 166592 77722
rect 166540 77658 166592 77664
rect 166632 77716 166684 77722
rect 166632 77658 166684 77664
rect 166356 77454 166408 77460
rect 166446 77480 166502 77489
rect 166264 74724 166316 74730
rect 166264 74666 166316 74672
rect 166264 73704 166316 73710
rect 166264 73646 166316 73652
rect 166172 73432 166224 73438
rect 166172 73374 166224 73380
rect 166078 70952 166134 70961
rect 166078 70887 166134 70896
rect 166092 31142 166120 70887
rect 166184 57254 166212 73374
rect 166276 61470 166304 73646
rect 166368 67046 166396 77454
rect 166446 77415 166502 77424
rect 166552 76820 166580 77658
rect 166644 77081 166672 77658
rect 166630 77072 166686 77081
rect 166630 77007 166686 77016
rect 166552 76792 166672 76820
rect 166644 73574 166672 76792
rect 166736 76265 166764 77744
rect 166816 77648 166868 77654
rect 166920 77625 166948 77744
rect 167058 77704 167086 78132
rect 167150 77772 167178 78132
rect 167242 77897 167270 78132
rect 167228 77888 167284 77897
rect 167228 77823 167284 77832
rect 167334 77772 167362 78132
rect 167150 77744 167224 77772
rect 167058 77676 167132 77704
rect 166816 77590 166868 77596
rect 166906 77616 166962 77625
rect 166722 76256 166778 76265
rect 166722 76191 166778 76200
rect 166722 76120 166778 76129
rect 166722 76055 166778 76064
rect 166736 73778 166764 76055
rect 166724 73772 166776 73778
rect 166724 73714 166776 73720
rect 166632 73568 166684 73574
rect 166632 73510 166684 73516
rect 166828 73438 166856 77590
rect 166906 77551 166962 77560
rect 166908 77512 166960 77518
rect 166908 77454 166960 77460
rect 166998 77480 167054 77489
rect 166920 77081 166948 77454
rect 166998 77415 167054 77424
rect 166906 77072 166962 77081
rect 166906 77007 166962 77016
rect 166906 76800 166962 76809
rect 167012 76770 167040 77415
rect 167104 77217 167132 77676
rect 167090 77208 167146 77217
rect 167090 77143 167146 77152
rect 167090 77072 167146 77081
rect 167090 77007 167146 77016
rect 166906 76735 166962 76744
rect 167000 76764 167052 76770
rect 166920 75914 166948 76735
rect 167000 76706 167052 76712
rect 166920 75886 167040 75914
rect 166906 75848 166962 75857
rect 166906 75783 166962 75792
rect 166920 73914 166948 75783
rect 167012 74534 167040 75886
rect 167104 75664 167132 77007
rect 167196 76344 167224 77744
rect 167288 77744 167362 77772
rect 167426 77772 167454 78132
rect 167518 77931 167546 78132
rect 167504 77922 167560 77931
rect 167504 77857 167560 77866
rect 167610 77772 167638 78132
rect 167702 77926 167730 78132
rect 167794 77926 167822 78132
rect 167690 77920 167742 77926
rect 167690 77862 167742 77868
rect 167782 77920 167834 77926
rect 167782 77862 167834 77868
rect 167886 77772 167914 78132
rect 167426 77744 167500 77772
rect 167288 76498 167316 77744
rect 167472 76922 167500 77744
rect 167564 77744 167638 77772
rect 167840 77744 167914 77772
rect 167978 77772 168006 78132
rect 168070 77897 168098 78132
rect 168162 77926 168190 78132
rect 168150 77920 168202 77926
rect 168056 77888 168112 77897
rect 168150 77862 168202 77868
rect 168056 77823 168112 77832
rect 168104 77784 168156 77790
rect 167978 77744 168052 77772
rect 167564 77568 167592 77744
rect 167736 77716 167788 77722
rect 167736 77658 167788 77664
rect 167564 77540 167684 77568
rect 167552 77444 167604 77450
rect 167552 77386 167604 77392
rect 167564 77353 167592 77386
rect 167550 77344 167606 77353
rect 167550 77279 167606 77288
rect 167472 76894 167592 76922
rect 167276 76492 167328 76498
rect 167276 76434 167328 76440
rect 167196 76316 167408 76344
rect 167274 76256 167330 76265
rect 167274 76191 167330 76200
rect 167104 75636 167224 75664
rect 167012 74506 167132 74534
rect 167000 74452 167052 74458
rect 167000 74394 167052 74400
rect 167012 74361 167040 74394
rect 166998 74352 167054 74361
rect 166998 74287 167054 74296
rect 166998 74216 167054 74225
rect 166998 74151 167054 74160
rect 166908 73908 166960 73914
rect 166908 73850 166960 73856
rect 167012 73817 167040 74151
rect 166998 73808 167054 73817
rect 166998 73743 167054 73752
rect 166816 73432 166868 73438
rect 166816 73374 166868 73380
rect 166356 67040 166408 67046
rect 166356 66982 166408 66988
rect 166264 61464 166316 61470
rect 166264 61406 166316 61412
rect 166172 57248 166224 57254
rect 166172 57190 166224 57196
rect 166080 31136 166132 31142
rect 166080 31078 166132 31084
rect 165988 31068 166040 31074
rect 165988 31010 166040 31016
rect 165896 28280 165948 28286
rect 165896 28222 165948 28228
rect 165804 21480 165856 21486
rect 165804 21422 165856 21428
rect 165620 21412 165672 21418
rect 165620 21354 165672 21360
rect 164516 19984 164568 19990
rect 164516 19926 164568 19932
rect 164424 15904 164476 15910
rect 164424 15846 164476 15852
rect 164332 13116 164384 13122
rect 164332 13058 164384 13064
rect 164240 10396 164292 10402
rect 164240 10338 164292 10344
rect 167104 10334 167132 74506
rect 167196 22914 167224 75636
rect 167288 22982 167316 76191
rect 167380 23050 167408 76316
rect 167564 76265 167592 76894
rect 167550 76256 167606 76265
rect 167550 76191 167606 76200
rect 167552 76152 167604 76158
rect 167552 76094 167604 76100
rect 167460 75676 167512 75682
rect 167460 75618 167512 75624
rect 167472 32502 167500 75618
rect 167564 75070 167592 76094
rect 167552 75064 167604 75070
rect 167552 75006 167604 75012
rect 167552 74928 167604 74934
rect 167552 74870 167604 74876
rect 167564 65618 167592 74870
rect 167656 65686 167684 77540
rect 167748 75682 167776 77658
rect 167736 75676 167788 75682
rect 167736 75618 167788 75624
rect 167840 74934 167868 77744
rect 168024 77294 168052 77744
rect 168254 77738 168282 78132
rect 168346 77926 168374 78132
rect 168438 77926 168466 78132
rect 168334 77920 168386 77926
rect 168334 77862 168386 77868
rect 168426 77920 168478 77926
rect 168426 77862 168478 77868
rect 168530 77772 168558 78132
rect 168622 77897 168650 78132
rect 168608 77888 168664 77897
rect 168608 77823 168664 77832
rect 168530 77744 168604 77772
rect 168104 77726 168156 77732
rect 167932 77266 168052 77294
rect 167932 75834 167960 77266
rect 168010 77208 168066 77217
rect 168010 77143 168066 77152
rect 168024 76158 168052 77143
rect 168116 76809 168144 77726
rect 168208 77710 168282 77738
rect 168102 76800 168158 76809
rect 168102 76735 168158 76744
rect 168104 76492 168156 76498
rect 168104 76434 168156 76440
rect 168012 76152 168064 76158
rect 168012 76094 168064 76100
rect 167932 75806 168052 75834
rect 167920 75744 167972 75750
rect 167920 75686 167972 75692
rect 167828 74928 167880 74934
rect 167828 74870 167880 74876
rect 167826 74760 167882 74769
rect 167826 74695 167882 74704
rect 167840 72486 167868 74695
rect 167828 72480 167880 72486
rect 167828 72422 167880 72428
rect 167932 70394 167960 75686
rect 167748 70366 167960 70394
rect 168024 70394 168052 75806
rect 168116 75750 168144 76434
rect 168208 75857 168236 77710
rect 168288 77648 168340 77654
rect 168576 77625 168604 77744
rect 168714 77704 168742 78132
rect 168668 77676 168742 77704
rect 168806 77704 168834 78132
rect 168898 77858 168926 78132
rect 168990 77926 169018 78132
rect 168978 77920 169030 77926
rect 168978 77862 169030 77868
rect 168886 77852 168938 77858
rect 168886 77794 168938 77800
rect 169082 77772 169110 78132
rect 169174 77897 169202 78132
rect 169160 77888 169216 77897
rect 169160 77823 169216 77832
rect 169036 77744 169110 77772
rect 168806 77676 168880 77704
rect 168288 77590 168340 77596
rect 168378 77616 168434 77625
rect 168300 76401 168328 77590
rect 168378 77551 168434 77560
rect 168562 77616 168618 77625
rect 168562 77551 168618 77560
rect 168286 76392 168342 76401
rect 168286 76327 168342 76336
rect 168194 75848 168250 75857
rect 168194 75783 168250 75792
rect 168104 75744 168156 75750
rect 168104 75686 168156 75692
rect 168288 74452 168340 74458
rect 168288 74394 168340 74400
rect 168300 73642 168328 74394
rect 168392 73846 168420 77551
rect 168564 77512 168616 77518
rect 168564 77454 168616 77460
rect 168470 76392 168526 76401
rect 168470 76327 168526 76336
rect 168380 73840 168432 73846
rect 168380 73782 168432 73788
rect 168288 73636 168340 73642
rect 168288 73578 168340 73584
rect 168380 72344 168432 72350
rect 168380 72286 168432 72292
rect 168024 70366 168236 70394
rect 167748 66978 167776 70366
rect 167736 66972 167788 66978
rect 167736 66914 167788 66920
rect 167644 65680 167696 65686
rect 167644 65622 167696 65628
rect 167552 65612 167604 65618
rect 167552 65554 167604 65560
rect 167460 32496 167512 32502
rect 167460 32438 167512 32444
rect 167368 23044 167420 23050
rect 167368 22986 167420 22992
rect 167276 22976 167328 22982
rect 167276 22918 167328 22924
rect 167184 22908 167236 22914
rect 167184 22850 167236 22856
rect 167092 10328 167144 10334
rect 167092 10270 167144 10276
rect 167184 5024 167236 5030
rect 167184 4966 167236 4972
rect 166080 3596 166132 3602
rect 166080 3538 166132 3544
rect 163780 3528 163832 3534
rect 163780 3470 163832 3476
rect 164884 3528 164936 3534
rect 164884 3470 164936 3476
rect 164896 480 164924 3470
rect 166092 480 166120 3538
rect 167196 480 167224 4966
rect 168208 4894 168236 70366
rect 168392 6186 168420 72286
rect 168484 18766 168512 76327
rect 168576 74594 168604 77454
rect 168668 76770 168696 77676
rect 168656 76764 168708 76770
rect 168656 76706 168708 76712
rect 168748 76560 168800 76566
rect 168748 76502 168800 76508
rect 168656 76492 168708 76498
rect 168656 76434 168708 76440
rect 168564 74588 168616 74594
rect 168564 74530 168616 74536
rect 168564 74384 168616 74390
rect 168564 74326 168616 74332
rect 168472 18760 168524 18766
rect 168472 18702 168524 18708
rect 168576 18698 168604 74326
rect 168668 73154 168696 76434
rect 168760 75274 168788 76502
rect 168748 75268 168800 75274
rect 168748 75210 168800 75216
rect 168668 73126 168788 73154
rect 168656 72412 168708 72418
rect 168656 72354 168708 72360
rect 168564 18692 168616 18698
rect 168564 18634 168616 18640
rect 168668 18630 168696 72354
rect 168760 72282 168788 73126
rect 168748 72276 168800 72282
rect 168748 72218 168800 72224
rect 168748 72140 168800 72146
rect 168748 72082 168800 72088
rect 168760 24206 168788 72082
rect 168852 24274 168880 77676
rect 168932 77648 168984 77654
rect 168932 77590 168984 77596
rect 168944 74390 168972 77590
rect 169036 75818 169064 77744
rect 169266 77704 169294 78132
rect 169358 77897 169386 78132
rect 169344 77888 169400 77897
rect 169344 77823 169400 77832
rect 169450 77704 169478 78132
rect 169542 77897 169570 78132
rect 169634 77926 169662 78132
rect 169622 77920 169674 77926
rect 169528 77888 169584 77897
rect 169622 77862 169674 77868
rect 169726 77858 169754 78132
rect 169528 77823 169584 77832
rect 169714 77852 169766 77858
rect 169714 77794 169766 77800
rect 169818 77738 169846 78132
rect 169220 77676 169294 77704
rect 169404 77676 169478 77704
rect 169576 77716 169628 77722
rect 169114 77616 169170 77625
rect 169114 77551 169170 77560
rect 169024 75812 169076 75818
rect 169024 75754 169076 75760
rect 169024 75676 169076 75682
rect 169024 75618 169076 75624
rect 168932 74384 168984 74390
rect 168932 74326 168984 74332
rect 168932 73840 168984 73846
rect 168932 73782 168984 73788
rect 168944 24342 168972 73782
rect 169036 68338 169064 75618
rect 169128 72418 169156 77551
rect 169116 72412 169168 72418
rect 169116 72354 169168 72360
rect 169220 72350 169248 77676
rect 169298 77616 169354 77625
rect 169298 77551 169354 77560
rect 169208 72344 169260 72350
rect 169208 72286 169260 72292
rect 169116 72276 169168 72282
rect 169116 72218 169168 72224
rect 169128 71058 169156 72218
rect 169312 72146 169340 77551
rect 169404 76498 169432 77676
rect 169576 77658 169628 77664
rect 169668 77716 169720 77722
rect 169668 77658 169720 77664
rect 169772 77710 169846 77738
rect 169482 77616 169538 77625
rect 169482 77551 169538 77560
rect 169392 76492 169444 76498
rect 169392 76434 169444 76440
rect 169392 76152 169444 76158
rect 169392 76094 169444 76100
rect 169404 75206 169432 76094
rect 169496 75682 169524 77551
rect 169484 75676 169536 75682
rect 169484 75618 169536 75624
rect 169392 75200 169444 75206
rect 169392 75142 169444 75148
rect 169392 74452 169444 74458
rect 169392 74394 169444 74400
rect 169404 74361 169432 74394
rect 169390 74352 169446 74361
rect 169390 74287 169446 74296
rect 169588 73681 169616 77658
rect 169680 76401 169708 77658
rect 169666 76392 169722 76401
rect 169666 76327 169722 76336
rect 169668 75812 169720 75818
rect 169668 75754 169720 75760
rect 169680 73710 169708 75754
rect 169772 74390 169800 77710
rect 169910 77636 169938 78132
rect 170002 77926 170030 78132
rect 169990 77920 170042 77926
rect 170094 77897 170122 78132
rect 169990 77862 170042 77868
rect 170080 77888 170136 77897
rect 170080 77823 170136 77832
rect 170186 77772 170214 78132
rect 170278 77931 170306 78132
rect 170264 77922 170320 77931
rect 170370 77926 170398 78132
rect 170264 77857 170320 77866
rect 170358 77920 170410 77926
rect 170358 77862 170410 77868
rect 170140 77744 170214 77772
rect 170312 77784 170364 77790
rect 169990 77716 170042 77722
rect 169990 77658 170042 77664
rect 169864 77608 169938 77636
rect 169760 74384 169812 74390
rect 169760 74326 169812 74332
rect 169760 73840 169812 73846
rect 169760 73782 169812 73788
rect 169668 73704 169720 73710
rect 169574 73672 169630 73681
rect 169668 73646 169720 73652
rect 169574 73607 169630 73616
rect 169300 72140 169352 72146
rect 169300 72082 169352 72088
rect 169116 71052 169168 71058
rect 169116 70994 169168 71000
rect 169024 68332 169076 68338
rect 169024 68274 169076 68280
rect 168932 24336 168984 24342
rect 168932 24278 168984 24284
rect 168840 24268 168892 24274
rect 168840 24210 168892 24216
rect 168748 24200 168800 24206
rect 168748 24142 168800 24148
rect 168656 18624 168708 18630
rect 168656 18566 168708 18572
rect 168380 6180 168432 6186
rect 168380 6122 168432 6128
rect 168196 4888 168248 4894
rect 168196 4830 168248 4836
rect 169772 4826 169800 73782
rect 169864 22846 169892 77608
rect 170002 77296 170030 77658
rect 170002 77268 170076 77296
rect 169944 75676 169996 75682
rect 169944 75618 169996 75624
rect 169956 24138 169984 75618
rect 170048 32434 170076 77268
rect 170140 75682 170168 77744
rect 170462 77761 170490 78132
rect 170312 77726 170364 77732
rect 170448 77752 170504 77761
rect 170324 77246 170352 77726
rect 170448 77687 170504 77696
rect 170404 77648 170456 77654
rect 170404 77590 170456 77596
rect 170312 77240 170364 77246
rect 170312 77182 170364 77188
rect 170416 76566 170444 77590
rect 170554 77466 170582 78132
rect 170646 77897 170674 78132
rect 170738 77926 170766 78132
rect 170726 77920 170778 77926
rect 170632 77888 170688 77897
rect 170726 77862 170778 77868
rect 170632 77823 170688 77832
rect 170680 77784 170732 77790
rect 170830 77772 170858 78132
rect 170680 77726 170732 77732
rect 170784 77744 170858 77772
rect 170554 77438 170628 77466
rect 170404 76560 170456 76566
rect 170404 76502 170456 76508
rect 170600 75721 170628 77438
rect 170310 75712 170366 75721
rect 170128 75676 170180 75682
rect 170310 75647 170366 75656
rect 170586 75712 170642 75721
rect 170586 75647 170642 75656
rect 170128 75618 170180 75624
rect 170218 75032 170274 75041
rect 170218 74967 170274 74976
rect 170128 74928 170180 74934
rect 170128 74870 170180 74876
rect 170140 33114 170168 74870
rect 170232 33794 170260 74967
rect 170324 61402 170352 75647
rect 170404 75132 170456 75138
rect 170404 75074 170456 75080
rect 170416 74730 170444 75074
rect 170496 74792 170548 74798
rect 170496 74734 170548 74740
rect 170404 74724 170456 74730
rect 170404 74666 170456 74672
rect 170404 74384 170456 74390
rect 170404 74326 170456 74332
rect 170416 65550 170444 74326
rect 170508 72457 170536 74734
rect 170692 73846 170720 77726
rect 170784 76922 170812 77744
rect 170922 77636 170950 78132
rect 171014 77897 171042 78132
rect 171000 77888 171056 77897
rect 171106 77858 171134 78132
rect 171198 77926 171226 78132
rect 171290 77926 171318 78132
rect 171382 77926 171410 78132
rect 171186 77920 171238 77926
rect 171186 77862 171238 77868
rect 171278 77920 171330 77926
rect 171278 77862 171330 77868
rect 171370 77920 171422 77926
rect 171370 77862 171422 77868
rect 171000 77823 171056 77832
rect 171094 77852 171146 77858
rect 171094 77794 171146 77800
rect 171474 77772 171502 78132
rect 171428 77744 171502 77772
rect 171566 77772 171594 78132
rect 171658 77897 171686 78132
rect 171750 77926 171778 78132
rect 171738 77920 171790 77926
rect 171644 77888 171700 77897
rect 171738 77862 171790 77868
rect 171644 77823 171700 77832
rect 171566 77744 171640 77772
rect 171428 77704 171456 77744
rect 171336 77676 171456 77704
rect 170922 77608 170996 77636
rect 170784 76894 170904 76922
rect 170772 76764 170824 76770
rect 170772 76706 170824 76712
rect 170784 74769 170812 76706
rect 170770 74760 170826 74769
rect 170770 74695 170826 74704
rect 170772 74588 170824 74594
rect 170772 74530 170824 74536
rect 170680 73840 170732 73846
rect 170680 73782 170732 73788
rect 170494 72448 170550 72457
rect 170494 72383 170550 72392
rect 170680 71800 170732 71806
rect 170680 71742 170732 71748
rect 170404 65544 170456 65550
rect 170404 65486 170456 65492
rect 170312 61396 170364 61402
rect 170312 61338 170364 61344
rect 170220 33788 170272 33794
rect 170220 33730 170272 33736
rect 170128 33108 170180 33114
rect 170128 33050 170180 33056
rect 170036 32428 170088 32434
rect 170036 32370 170088 32376
rect 169944 24132 169996 24138
rect 169944 24074 169996 24080
rect 169852 22840 169904 22846
rect 169852 22782 169904 22788
rect 170692 5030 170720 71742
rect 170784 66910 170812 74530
rect 170876 73273 170904 76894
rect 170968 74934 170996 77608
rect 171138 77344 171194 77353
rect 171138 77279 171194 77288
rect 171152 76770 171180 77279
rect 171140 76764 171192 76770
rect 171140 76706 171192 76712
rect 171336 76634 171364 77676
rect 171508 77580 171560 77586
rect 171508 77522 171560 77528
rect 171520 77353 171548 77522
rect 171506 77344 171562 77353
rect 171506 77279 171562 77288
rect 171612 77081 171640 77744
rect 171842 77738 171870 78132
rect 171934 77926 171962 78132
rect 172026 77926 172054 78132
rect 171922 77920 171974 77926
rect 171922 77862 171974 77868
rect 172014 77920 172066 77926
rect 172014 77862 172066 77868
rect 171842 77710 171916 77738
rect 172118 77722 172146 78132
rect 172210 77897 172238 78132
rect 172196 77888 172252 77897
rect 172196 77823 172252 77832
rect 172302 77738 172330 78132
rect 172394 77931 172422 78132
rect 172380 77922 172436 77931
rect 172380 77857 172436 77866
rect 172486 77738 172514 78132
rect 171692 77648 171744 77654
rect 171692 77590 171744 77596
rect 171784 77648 171836 77654
rect 171784 77590 171836 77596
rect 171704 77246 171732 77590
rect 171692 77240 171744 77246
rect 171692 77182 171744 77188
rect 171598 77072 171654 77081
rect 171598 77007 171654 77016
rect 171796 76809 171824 77590
rect 171782 76800 171838 76809
rect 171782 76735 171838 76744
rect 171048 76628 171100 76634
rect 171048 76570 171100 76576
rect 171324 76628 171376 76634
rect 171324 76570 171376 76576
rect 170956 74928 171008 74934
rect 170956 74870 171008 74876
rect 170862 73264 170918 73273
rect 170862 73199 170918 73208
rect 171060 71602 171088 76570
rect 171140 76220 171192 76226
rect 171140 76162 171192 76168
rect 171152 74526 171180 76162
rect 171784 74928 171836 74934
rect 171784 74870 171836 74876
rect 171508 74656 171560 74662
rect 171508 74598 171560 74604
rect 171690 74624 171746 74633
rect 171140 74520 171192 74526
rect 171140 74462 171192 74468
rect 171048 71596 171100 71602
rect 171048 71538 171100 71544
rect 170772 66904 170824 66910
rect 170772 66846 170824 66852
rect 171520 42090 171548 74598
rect 171690 74559 171746 74568
rect 171508 42084 171560 42090
rect 171508 42026 171560 42032
rect 171704 24410 171732 74559
rect 171796 71738 171824 74870
rect 171888 74798 171916 77710
rect 171968 77716 172020 77722
rect 171968 77658 172020 77664
rect 172106 77716 172158 77722
rect 172302 77710 172376 77738
rect 172106 77658 172158 77664
rect 171980 77489 172008 77658
rect 172244 77648 172296 77654
rect 172164 77596 172244 77602
rect 172164 77590 172296 77596
rect 172060 77580 172112 77586
rect 172060 77522 172112 77528
rect 172164 77574 172284 77590
rect 171966 77480 172022 77489
rect 172072 77450 172100 77522
rect 172164 77489 172192 77574
rect 172150 77480 172206 77489
rect 171966 77415 172022 77424
rect 172060 77444 172112 77450
rect 172150 77415 172206 77424
rect 172244 77444 172296 77450
rect 172060 77386 172112 77392
rect 172244 77386 172296 77392
rect 172058 77344 172114 77353
rect 172058 77279 172114 77288
rect 171968 77172 172020 77178
rect 171968 77114 172020 77120
rect 171980 76498 172008 77114
rect 171968 76492 172020 76498
rect 171968 76434 172020 76440
rect 172072 76430 172100 77279
rect 172060 76424 172112 76430
rect 172060 76366 172112 76372
rect 172256 76362 172284 77386
rect 172348 76430 172376 77710
rect 172440 77710 172514 77738
rect 172440 77489 172468 77710
rect 172578 77636 172606 78132
rect 172670 77704 172698 78132
rect 172762 77897 172790 78132
rect 172748 77888 172804 77897
rect 172748 77823 172804 77832
rect 172854 77738 172882 78132
rect 172808 77710 172882 77738
rect 172946 77738 172974 78132
rect 173038 77926 173066 78132
rect 173026 77920 173078 77926
rect 173026 77862 173078 77868
rect 173130 77738 173158 78132
rect 172946 77710 173020 77738
rect 172670 77676 172744 77704
rect 172578 77608 172652 77636
rect 172426 77480 172482 77489
rect 172426 77415 172482 77424
rect 172336 76424 172388 76430
rect 172336 76366 172388 76372
rect 172244 76356 172296 76362
rect 172244 76298 172296 76304
rect 172624 75818 172652 77608
rect 172716 76226 172744 77676
rect 172704 76220 172756 76226
rect 172704 76162 172756 76168
rect 172612 75812 172664 75818
rect 172612 75754 172664 75760
rect 172334 75440 172390 75449
rect 172334 75375 172390 75384
rect 172244 74860 172296 74866
rect 172244 74802 172296 74808
rect 171876 74792 171928 74798
rect 171876 74734 171928 74740
rect 171966 73808 172022 73817
rect 171876 73772 171928 73778
rect 171966 73743 172022 73752
rect 171876 73714 171928 73720
rect 171784 71732 171836 71738
rect 171784 71674 171836 71680
rect 171784 71596 171836 71602
rect 171784 71538 171836 71544
rect 171692 24404 171744 24410
rect 171692 24346 171744 24352
rect 170680 5024 170732 5030
rect 170680 4966 170732 4972
rect 169760 4820 169812 4826
rect 169760 4762 169812 4768
rect 171796 3738 171824 71538
rect 171784 3732 171836 3738
rect 171784 3674 171836 3680
rect 171888 3670 171916 73714
rect 171980 5386 172008 73743
rect 172060 72820 172112 72826
rect 172060 72762 172112 72768
rect 172072 5522 172100 72762
rect 172150 70000 172206 70009
rect 172150 69935 172206 69944
rect 172164 6914 172192 69935
rect 172256 10538 172284 74802
rect 172348 14550 172376 75375
rect 172808 74534 172836 77710
rect 172992 77353 173020 77710
rect 173084 77710 173158 77738
rect 172978 77344 173034 77353
rect 172978 77279 173034 77288
rect 173084 76401 173112 77710
rect 173222 77636 173250 78132
rect 173176 77608 173250 77636
rect 173314 77636 173342 78132
rect 173406 77738 173434 78132
rect 173498 77897 173526 78132
rect 173484 77888 173540 77897
rect 173484 77823 173540 77832
rect 173590 77772 173618 78132
rect 173682 77926 173710 78132
rect 173774 77926 173802 78132
rect 173670 77920 173722 77926
rect 173670 77862 173722 77868
rect 173762 77920 173814 77926
rect 173866 77897 173894 78132
rect 173762 77862 173814 77868
rect 173852 77888 173908 77897
rect 173852 77823 173908 77832
rect 173958 77772 173986 78132
rect 173544 77744 173618 77772
rect 173912 77744 173986 77772
rect 173406 77710 173480 77738
rect 173314 77625 173388 77636
rect 173314 77616 173402 77625
rect 173314 77608 173346 77616
rect 173176 76537 173204 77608
rect 173346 77551 173402 77560
rect 173452 76673 173480 77710
rect 173544 76945 173572 77744
rect 173624 77648 173676 77654
rect 173622 77616 173624 77625
rect 173676 77616 173678 77625
rect 173622 77551 173678 77560
rect 173530 76936 173586 76945
rect 173530 76871 173586 76880
rect 173438 76664 173494 76673
rect 173438 76599 173494 76608
rect 173162 76528 173218 76537
rect 173912 76498 173940 77744
rect 174050 77636 174078 78132
rect 174142 77738 174170 78132
rect 174234 77874 174262 78132
rect 174358 77888 174414 77897
rect 174234 77846 174308 77874
rect 174142 77710 174216 77738
rect 174004 77608 174078 77636
rect 174004 77110 174032 77608
rect 173992 77104 174044 77110
rect 173992 77046 174044 77052
rect 174188 77042 174216 77710
rect 174176 77036 174228 77042
rect 174176 76978 174228 76984
rect 173162 76463 173218 76472
rect 173900 76492 173952 76498
rect 173900 76434 173952 76440
rect 173070 76392 173126 76401
rect 173070 76327 173126 76336
rect 172978 76256 173034 76265
rect 172978 76191 173034 76200
rect 172716 74506 172836 74534
rect 172716 73642 172744 74506
rect 172992 74458 173020 76191
rect 173164 75744 173216 75750
rect 173164 75686 173216 75692
rect 172980 74452 173032 74458
rect 172980 74394 173032 74400
rect 172704 73636 172756 73642
rect 172704 73578 172756 73584
rect 172428 73500 172480 73506
rect 172428 73442 172480 73448
rect 172440 18902 172468 73442
rect 172518 65512 172574 65521
rect 172518 65447 172574 65456
rect 172428 18896 172480 18902
rect 172428 18838 172480 18844
rect 172532 16574 172560 65447
rect 172532 16546 172744 16574
rect 172336 14544 172388 14550
rect 172336 14486 172388 14492
rect 172244 10532 172296 10538
rect 172244 10474 172296 10480
rect 172164 6886 172284 6914
rect 172072 5494 172192 5522
rect 171980 5358 172100 5386
rect 171968 5296 172020 5302
rect 171968 5238 172020 5244
rect 169576 3664 169628 3670
rect 169576 3606 169628 3612
rect 171876 3664 171928 3670
rect 171876 3606 171928 3612
rect 168380 3324 168432 3330
rect 168380 3266 168432 3272
rect 168392 480 168420 3266
rect 169588 480 169616 3606
rect 170772 3392 170824 3398
rect 170772 3334 170824 3340
rect 170784 480 170812 3334
rect 171980 480 172008 5238
rect 172072 3806 172100 5358
rect 172060 3800 172112 3806
rect 172060 3742 172112 3748
rect 172164 3602 172192 5494
rect 172152 3596 172204 3602
rect 172152 3538 172204 3544
rect 172256 3534 172284 6886
rect 172244 3528 172296 3534
rect 172244 3470 172296 3476
rect 142406 354 142518 480
rect 142264 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 173176 3126 173204 75686
rect 173440 75064 173492 75070
rect 173440 75006 173492 75012
rect 173348 74996 173400 75002
rect 173348 74938 173400 74944
rect 173254 70408 173310 70417
rect 173254 70343 173310 70352
rect 173268 3466 173296 70343
rect 173360 20194 173388 74938
rect 173452 21758 173480 75006
rect 173898 72992 173954 73001
rect 173898 72927 173954 72936
rect 173440 21752 173492 21758
rect 173440 21694 173492 21700
rect 173348 20188 173400 20194
rect 173348 20130 173400 20136
rect 173256 3460 173308 3466
rect 173256 3402 173308 3408
rect 173164 3120 173216 3126
rect 173164 3062 173216 3068
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173912 354 173940 72927
rect 174280 72418 174308 77846
rect 174358 77823 174414 77832
rect 174372 76294 174400 77823
rect 174360 76288 174412 76294
rect 174360 76230 174412 76236
rect 174268 72412 174320 72418
rect 174268 72354 174320 72360
rect 174464 67634 174492 78254
rect 174556 77926 174584 78610
rect 178972 78577 179000 79290
rect 178958 78568 179014 78577
rect 178958 78503 179014 78512
rect 175924 78464 175976 78470
rect 174818 78432 174874 78441
rect 175924 78406 175976 78412
rect 174818 78367 174874 78376
rect 174636 78328 174688 78334
rect 174636 78270 174688 78276
rect 174648 77994 174676 78270
rect 174728 78260 174780 78266
rect 174728 78202 174780 78208
rect 174636 77988 174688 77994
rect 174636 77930 174688 77936
rect 174544 77920 174596 77926
rect 174544 77862 174596 77868
rect 174542 75576 174598 75585
rect 174740 75546 174768 78202
rect 174832 78198 174860 78367
rect 174820 78192 174872 78198
rect 174820 78134 174872 78140
rect 175646 77752 175702 77761
rect 175646 77687 175702 77696
rect 175830 77752 175886 77761
rect 175936 77722 175964 78406
rect 180076 78130 180104 191830
rect 180156 151836 180208 151842
rect 180156 151778 180208 151784
rect 180168 78441 180196 151778
rect 180812 122777 180840 231066
rect 180984 213988 181036 213994
rect 180984 213930 181036 213936
rect 180890 135416 180946 135425
rect 180890 135351 180946 135360
rect 180798 122768 180854 122777
rect 180798 122703 180854 122712
rect 180248 111852 180300 111858
rect 180248 111794 180300 111800
rect 180154 78432 180210 78441
rect 180154 78367 180210 78376
rect 180064 78124 180116 78130
rect 180064 78066 180116 78072
rect 176290 77888 176346 77897
rect 176108 77852 176160 77858
rect 176290 77823 176346 77832
rect 176108 77794 176160 77800
rect 175830 77687 175832 77696
rect 174542 75511 174598 75520
rect 174728 75540 174780 75546
rect 174372 67606 174492 67634
rect 174372 23254 174400 67606
rect 174556 32638 174584 75511
rect 174728 75482 174780 75488
rect 175660 74769 175688 77687
rect 175884 77687 175886 77696
rect 175924 77716 175976 77722
rect 175832 77658 175884 77664
rect 175924 77658 175976 77664
rect 175830 77616 175886 77625
rect 175830 77551 175832 77560
rect 175884 77551 175886 77560
rect 175924 77580 175976 77586
rect 175832 77522 175884 77528
rect 175924 77522 175976 77528
rect 175830 77480 175886 77489
rect 175830 77415 175886 77424
rect 175844 76430 175872 77415
rect 175936 76770 175964 77522
rect 175924 76764 175976 76770
rect 175924 76706 175976 76712
rect 176120 76634 176148 77794
rect 176304 77081 176332 77823
rect 178406 77208 178462 77217
rect 180260 77178 180288 111794
rect 180340 99408 180392 99414
rect 180340 99350 180392 99356
rect 180352 78742 180380 99350
rect 180340 78736 180392 78742
rect 180340 78678 180392 78684
rect 178406 77143 178462 77152
rect 180248 77172 180300 77178
rect 176290 77072 176346 77081
rect 176290 77007 176346 77016
rect 178420 76770 178448 77143
rect 180248 77114 180300 77120
rect 178408 76764 178460 76770
rect 178408 76706 178460 76712
rect 176108 76628 176160 76634
rect 176108 76570 176160 76576
rect 176200 76628 176252 76634
rect 176200 76570 176252 76576
rect 175832 76424 175884 76430
rect 175832 76366 175884 76372
rect 176212 76129 176240 76570
rect 176198 76120 176254 76129
rect 176198 76055 176254 76064
rect 175646 74760 175702 74769
rect 175646 74695 175702 74704
rect 174636 72412 174688 72418
rect 174636 72354 174688 72360
rect 174648 45558 174676 72354
rect 175278 63064 175334 63073
rect 175278 62999 175334 63008
rect 174636 45552 174688 45558
rect 174636 45494 174688 45500
rect 174544 32632 174596 32638
rect 174544 32574 174596 32580
rect 174360 23248 174412 23254
rect 174360 23190 174412 23196
rect 175292 16574 175320 62999
rect 180800 46232 180852 46238
rect 180800 46174 180852 46180
rect 176658 33960 176714 33969
rect 176658 33895 176714 33904
rect 175292 16546 175504 16574
rect 175476 480 175504 16546
rect 176672 11694 176700 33895
rect 176752 26036 176804 26042
rect 176752 25978 176804 25984
rect 176660 11688 176712 11694
rect 176660 11630 176712 11636
rect 176764 6914 176792 25978
rect 179420 25968 179472 25974
rect 179420 25910 179472 25916
rect 179432 16574 179460 25910
rect 180812 16574 180840 46174
rect 180904 33046 180932 135351
rect 180996 129713 181024 213930
rect 189724 205692 189776 205698
rect 189724 205634 189776 205640
rect 188344 165640 188396 165646
rect 188344 165582 188396 165588
rect 182364 163600 182416 163606
rect 182364 163542 182416 163548
rect 182272 142928 182324 142934
rect 182272 142870 182324 142876
rect 181076 141704 181128 141710
rect 181076 141646 181128 141652
rect 180982 129704 181038 129713
rect 180982 129639 181038 129648
rect 181088 115297 181116 141646
rect 181168 137964 181220 137970
rect 181168 137906 181220 137912
rect 181074 115288 181130 115297
rect 181074 115223 181130 115232
rect 181180 113121 181208 137906
rect 182180 136672 182232 136678
rect 182180 136614 182232 136620
rect 182192 133249 182220 136614
rect 182178 133240 182234 133249
rect 182178 133175 182234 133184
rect 182284 124137 182312 142870
rect 182376 128353 182404 163542
rect 182916 163532 182968 163538
rect 182916 163474 182968 163480
rect 182732 143064 182784 143070
rect 182732 143006 182784 143012
rect 182640 141636 182692 141642
rect 182640 141578 182692 141584
rect 182456 138916 182508 138922
rect 182456 138858 182508 138864
rect 182362 128344 182418 128353
rect 182362 128279 182418 128288
rect 182270 124128 182326 124137
rect 182270 124063 182326 124072
rect 181166 113112 181222 113121
rect 181166 113047 181222 113056
rect 182468 110401 182496 138858
rect 182548 138780 182600 138786
rect 182548 138722 182600 138728
rect 182560 116793 182588 138722
rect 182652 119785 182680 141578
rect 182744 125361 182772 143006
rect 182824 142996 182876 143002
rect 182824 142938 182876 142944
rect 182730 125352 182786 125361
rect 182730 125287 182786 125296
rect 182836 121281 182864 142938
rect 182928 126993 182956 163474
rect 183006 133920 183062 133929
rect 183006 133855 183062 133864
rect 182914 126984 182970 126993
rect 182914 126919 182970 126928
rect 182822 121272 182878 121281
rect 182822 121207 182878 121216
rect 182638 119776 182694 119785
rect 182638 119711 182694 119720
rect 182546 116784 182602 116793
rect 182546 116719 182602 116728
rect 182454 110392 182510 110401
rect 182454 110327 182510 110336
rect 182824 100700 182876 100706
rect 182824 100642 182876 100648
rect 182836 100201 182864 100642
rect 182822 100192 182878 100201
rect 182822 100127 182878 100136
rect 182824 99340 182876 99346
rect 182824 99282 182876 99288
rect 182836 98841 182864 99282
rect 182822 98832 182878 98841
rect 182822 98767 182878 98776
rect 182272 89684 182324 89690
rect 182272 89626 182324 89632
rect 182284 89457 182312 89626
rect 182270 89448 182326 89457
rect 182270 89383 182326 89392
rect 182272 85604 182324 85610
rect 182272 85546 182324 85552
rect 182180 85536 182232 85542
rect 182180 85478 182232 85484
rect 182192 85105 182220 85478
rect 182178 85096 182234 85105
rect 182178 85031 182234 85040
rect 182284 83881 182312 85546
rect 182270 83872 182326 83881
rect 182270 83807 182326 83816
rect 182822 81560 182878 81569
rect 182822 81495 182878 81504
rect 181442 77888 181498 77897
rect 181442 77823 181498 77832
rect 181456 77489 181484 77823
rect 181442 77480 181498 77489
rect 181442 77415 181498 77424
rect 182180 67244 182232 67250
rect 182180 67186 182232 67192
rect 180892 33040 180944 33046
rect 180892 32982 180944 32988
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 177856 11688 177908 11694
rect 177856 11630 177908 11636
rect 176672 6886 176792 6914
rect 176672 480 176700 6886
rect 177868 480 177896 11630
rect 179052 3120 179104 3126
rect 179052 3062 179104 3068
rect 179064 480 179092 3062
rect 180260 480 180288 16546
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 173134 -960 173246 326
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 67186
rect 182836 46918 182864 81495
rect 183020 74934 183048 133855
rect 184204 125656 184256 125662
rect 184204 125598 184256 125604
rect 183468 108996 183520 109002
rect 183468 108938 183520 108944
rect 183480 108905 183508 108938
rect 183466 108896 183522 108905
rect 183466 108831 183522 108840
rect 183468 107636 183520 107642
rect 183468 107578 183520 107584
rect 183480 107409 183508 107578
rect 183466 107400 183522 107409
rect 183466 107335 183522 107344
rect 183468 106276 183520 106282
rect 183468 106218 183520 106224
rect 183480 106049 183508 106218
rect 183466 106040 183522 106049
rect 183466 105975 183522 105984
rect 183468 104848 183520 104854
rect 183468 104790 183520 104796
rect 183480 104553 183508 104790
rect 183466 104544 183522 104553
rect 183466 104479 183522 104488
rect 183468 103488 183520 103494
rect 183468 103430 183520 103436
rect 183480 103057 183508 103430
rect 183466 103048 183522 103057
rect 183466 102983 183522 102992
rect 183468 102128 183520 102134
rect 183468 102070 183520 102076
rect 183480 101697 183508 102070
rect 183466 101688 183522 101697
rect 183466 101623 183522 101632
rect 183468 97980 183520 97986
rect 183468 97922 183520 97928
rect 183480 97345 183508 97922
rect 183466 97336 183522 97345
rect 183466 97271 183522 97280
rect 183468 95192 183520 95198
rect 183466 95160 183468 95169
rect 183520 95160 183522 95169
rect 183466 95095 183522 95104
rect 183468 93832 183520 93838
rect 183466 93800 183468 93809
rect 183520 93800 183522 93809
rect 183466 93735 183522 93744
rect 183468 92472 183520 92478
rect 183468 92414 183520 92420
rect 183480 92313 183508 92414
rect 183466 92304 183522 92313
rect 183466 92239 183522 92248
rect 183468 91044 183520 91050
rect 183468 90986 183520 90992
rect 183480 90953 183508 90986
rect 183466 90944 183522 90953
rect 183466 90879 183522 90888
rect 183468 88188 183520 88194
rect 183468 88130 183520 88136
rect 183480 88097 183508 88130
rect 183466 88088 183522 88097
rect 183466 88023 183522 88032
rect 183468 86896 183520 86902
rect 183468 86838 183520 86844
rect 183480 86601 183508 86838
rect 183466 86592 183522 86601
rect 183466 86527 183522 86536
rect 184216 85542 184244 125598
rect 188356 86902 188384 165582
rect 189736 88194 189764 205634
rect 207032 198014 207060 230588
rect 236012 230574 236578 230602
rect 207020 198008 207072 198014
rect 207020 197950 207072 197956
rect 236012 196654 236040 230574
rect 266556 228478 266584 230588
rect 266544 228472 266596 228478
rect 266544 228414 266596 228420
rect 236644 228404 236696 228410
rect 236644 228346 236696 228352
rect 236656 196722 236684 228346
rect 296732 199442 296760 230588
rect 327092 228478 327120 230588
rect 356072 230574 356546 230602
rect 297364 228472 297416 228478
rect 297364 228414 297416 228420
rect 327080 228472 327132 228478
rect 327080 228414 327132 228420
rect 296720 199436 296772 199442
rect 296720 199378 296772 199384
rect 236644 196716 236696 196722
rect 236644 196658 236696 196664
rect 236000 196648 236052 196654
rect 236000 196590 236052 196596
rect 297376 195906 297404 228414
rect 356072 195974 356100 230574
rect 385696 220862 385724 231066
rect 386524 228410 386552 230588
rect 386512 228404 386564 228410
rect 386512 228346 386564 228352
rect 391204 227724 391256 227730
rect 391204 227666 391256 227672
rect 389824 223100 389876 223106
rect 389824 223042 389876 223048
rect 378048 220856 378100 220862
rect 378048 220798 378100 220804
rect 385684 220856 385736 220862
rect 385684 220798 385736 220804
rect 378060 215966 378088 220798
rect 367744 215960 367796 215966
rect 367744 215902 367796 215908
rect 378048 215960 378100 215966
rect 378048 215902 378100 215908
rect 367756 206310 367784 215902
rect 378784 210452 378836 210458
rect 378784 210394 378836 210400
rect 356704 206304 356756 206310
rect 356704 206246 356756 206252
rect 367744 206304 367796 206310
rect 367744 206246 367796 206252
rect 356060 195968 356112 195974
rect 356060 195910 356112 195916
rect 297364 195900 297416 195906
rect 297364 195842 297416 195848
rect 356716 174622 356744 206246
rect 371240 186992 371292 186998
rect 371240 186934 371292 186940
rect 371252 183938 371280 186934
rect 369124 183932 369176 183938
rect 369124 183874 369176 183880
rect 371240 183932 371292 183938
rect 371240 183874 371292 183880
rect 350540 174616 350592 174622
rect 350540 174558 350592 174564
rect 356704 174616 356756 174622
rect 356704 174558 356756 174564
rect 350552 172378 350580 174558
rect 348424 172372 348476 172378
rect 348424 172314 348476 172320
rect 350540 172372 350592 172378
rect 350540 172314 350592 172320
rect 339868 147008 339920 147014
rect 339868 146950 339920 146956
rect 339880 144362 339908 146950
rect 336004 144356 336056 144362
rect 336004 144298 336056 144304
rect 339868 144356 339920 144362
rect 339868 144298 339920 144304
rect 336016 142186 336044 144298
rect 348436 144294 348464 172314
rect 366732 157752 366784 157758
rect 366732 157694 366784 157700
rect 359464 156732 359516 156738
rect 359464 156674 359516 156680
rect 353944 156664 353996 156670
rect 353944 156606 353996 156612
rect 353956 147014 353984 156606
rect 353944 147008 353996 147014
rect 353944 146950 353996 146956
rect 343640 144288 343692 144294
rect 343640 144230 343692 144236
rect 348424 144288 348476 144294
rect 348424 144230 348476 144236
rect 330944 142180 330996 142186
rect 330944 142122 330996 142128
rect 336004 142180 336056 142186
rect 336004 142122 336056 142128
rect 326344 141636 326396 141642
rect 326344 141578 326396 141584
rect 320180 138780 320232 138786
rect 320180 138722 320232 138728
rect 320192 137018 320220 138722
rect 318248 137012 318300 137018
rect 318248 136954 318300 136960
rect 320180 137012 320232 137018
rect 320180 136954 320232 136960
rect 318260 135930 318288 136954
rect 306748 135924 306800 135930
rect 306748 135866 306800 135872
rect 318248 135924 318300 135930
rect 318248 135866 318300 135872
rect 306760 133958 306788 135866
rect 305000 133952 305052 133958
rect 305000 133894 305052 133900
rect 306748 133952 306800 133958
rect 306748 133894 306800 133900
rect 305012 128382 305040 133894
rect 300768 128376 300820 128382
rect 300768 128318 300820 128324
rect 305000 128376 305052 128382
rect 305000 128318 305052 128324
rect 300780 123486 300808 128318
rect 326356 126274 326384 141578
rect 330956 138786 330984 142122
rect 343652 141642 343680 144230
rect 343640 141636 343692 141642
rect 343640 141578 343692 141584
rect 330944 138780 330996 138786
rect 330944 138722 330996 138728
rect 359476 137290 359504 156674
rect 366744 156670 366772 157694
rect 369136 156738 369164 183874
rect 378796 172582 378824 210394
rect 389836 186998 389864 223042
rect 391216 212226 391244 227666
rect 389916 212220 389968 212226
rect 389916 212162 389968 212168
rect 391204 212220 391256 212226
rect 391204 212162 391256 212168
rect 389824 186992 389876 186998
rect 389824 186934 389876 186940
rect 389928 186386 389956 212162
rect 387800 186380 387852 186386
rect 387800 186322 387852 186328
rect 389916 186380 389968 186386
rect 389916 186322 389968 186328
rect 387812 183598 387840 186322
rect 387800 183592 387852 183598
rect 387800 183534 387852 183540
rect 385040 183524 385092 183530
rect 385040 183466 385092 183472
rect 385052 179450 385080 183466
rect 384304 179444 384356 179450
rect 384304 179386 384356 179392
rect 385040 179444 385092 179450
rect 385040 179386 385092 179392
rect 378784 172576 378836 172582
rect 378784 172518 378836 172524
rect 376116 172508 376168 172514
rect 376116 172450 376168 172456
rect 376024 170400 376076 170406
rect 376024 170342 376076 170348
rect 374000 162852 374052 162858
rect 374000 162794 374052 162800
rect 374012 158794 374040 162794
rect 373920 158766 374040 158794
rect 373920 157758 373948 158766
rect 373908 157752 373960 157758
rect 373908 157694 373960 157700
rect 376036 157418 376064 170342
rect 376128 162858 376156 172450
rect 384316 170406 384344 179386
rect 384304 170400 384356 170406
rect 384304 170342 384356 170348
rect 376116 162852 376168 162858
rect 376116 162794 376168 162800
rect 375012 157412 375064 157418
rect 375012 157354 375064 157360
rect 376024 157412 376076 157418
rect 376024 157354 376076 157360
rect 369124 156732 369176 156738
rect 369124 156674 369176 156680
rect 366732 156664 366784 156670
rect 366732 156606 366784 156612
rect 375024 153270 375052 157354
rect 373356 153264 373408 153270
rect 373356 153206 373408 153212
rect 375012 153264 375064 153270
rect 375012 153206 375064 153212
rect 373368 146266 373396 153206
rect 371884 146260 371936 146266
rect 371884 146202 371936 146208
rect 373356 146260 373408 146266
rect 373356 146202 373408 146208
rect 371896 140826 371924 146202
rect 369860 140820 369912 140826
rect 369860 140762 369912 140768
rect 371884 140820 371936 140826
rect 371884 140762 371936 140768
rect 369872 137358 369900 140762
rect 366364 137352 366416 137358
rect 366364 137294 366416 137300
rect 369860 137352 369912 137358
rect 369860 137294 369912 137300
rect 359464 137284 359516 137290
rect 359464 137226 359516 137232
rect 366376 129946 366404 137294
rect 361948 129940 362000 129946
rect 361948 129882 362000 129888
rect 366364 129940 366416 129946
rect 366364 129882 366416 129888
rect 314660 126268 314712 126274
rect 314660 126210 314712 126216
rect 326344 126268 326396 126274
rect 326344 126210 326396 126216
rect 314672 123962 314700 126210
rect 312176 123956 312228 123962
rect 312176 123898 312228 123904
rect 314660 123956 314712 123962
rect 314660 123898 314712 123904
rect 295248 123480 295300 123486
rect 295248 123422 295300 123428
rect 300768 123480 300820 123486
rect 300768 123422 300820 123428
rect 295260 117434 295288 123422
rect 312188 117570 312216 123898
rect 361960 123690 361988 129882
rect 360936 123684 360988 123690
rect 360936 123626 360988 123632
rect 361948 123684 362000 123690
rect 361948 123626 362000 123632
rect 360948 117570 360976 123626
rect 307024 117564 307076 117570
rect 307024 117506 307076 117512
rect 312176 117564 312228 117570
rect 312176 117506 312228 117512
rect 358820 117564 358872 117570
rect 358820 117506 358872 117512
rect 360936 117564 360988 117570
rect 360936 117506 360988 117512
rect 292580 117428 292632 117434
rect 292580 117370 292632 117376
rect 295248 117428 295300 117434
rect 295248 117370 295300 117376
rect 292592 114306 292620 117370
rect 291108 114300 291160 114306
rect 291108 114242 291160 114248
rect 292580 114300 292632 114306
rect 292580 114242 292632 114248
rect 291120 107710 291148 114242
rect 307036 111110 307064 117506
rect 358832 115938 358860 117506
rect 354680 115932 354732 115938
rect 354680 115874 354732 115880
rect 358820 115932 358872 115938
rect 358820 115874 358872 115880
rect 354692 113234 354720 115874
rect 354600 113206 354720 113234
rect 303620 111104 303672 111110
rect 303620 111046 303672 111052
rect 307024 111104 307076 111110
rect 307024 111046 307076 111052
rect 291108 107704 291160 107710
rect 291108 107646 291160 107652
rect 303632 105602 303660 111046
rect 354600 109002 354628 113206
rect 354588 108996 354640 109002
rect 354588 108938 354640 108944
rect 291844 105596 291896 105602
rect 291844 105538 291896 105544
rect 303620 105596 303672 105602
rect 303620 105538 303672 105544
rect 189724 88188 189776 88194
rect 189724 88130 189776 88136
rect 291856 87650 291884 105538
rect 284944 87644 284996 87650
rect 284944 87586 284996 87592
rect 291844 87644 291896 87650
rect 291844 87586 291896 87592
rect 188344 86896 188396 86902
rect 188344 86838 188396 86844
rect 184204 85536 184256 85542
rect 184204 85478 184256 85484
rect 183466 80200 183522 80209
rect 183466 80135 183522 80144
rect 183480 80102 183508 80135
rect 183468 80096 183520 80102
rect 183468 80038 183520 80044
rect 231860 77716 231912 77722
rect 231860 77658 231912 77664
rect 200120 77648 200172 77654
rect 200120 77590 200172 77596
rect 195980 76084 196032 76090
rect 195980 76026 196032 76032
rect 183008 74928 183060 74934
rect 183008 74870 183060 74876
rect 184940 71460 184992 71466
rect 184940 71402 184992 71408
rect 182824 46912 182876 46918
rect 182824 46854 182876 46860
rect 183560 25900 183612 25906
rect 183560 25842 183612 25848
rect 183572 16574 183600 25842
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 184952 480 184980 71402
rect 190460 68604 190512 68610
rect 190460 68546 190512 68552
rect 189080 64592 189132 64598
rect 189080 64534 189132 64540
rect 185032 63164 185084 63170
rect 185032 63106 185084 63112
rect 185044 16574 185072 63106
rect 186320 25832 186372 25838
rect 186320 25774 186372 25780
rect 186332 16574 186360 25774
rect 187700 24540 187752 24546
rect 187700 24482 187752 24488
rect 187712 16574 187740 24482
rect 189092 16574 189120 64534
rect 185044 16546 186176 16574
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 189092 16546 189304 16574
rect 186148 480 186176 16546
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189276 354 189304 16546
rect 189694 354 189806 480
rect 189276 326 189806 354
rect 190472 354 190500 68546
rect 193218 62928 193274 62937
rect 193218 62863 193274 62872
rect 191838 18728 191894 18737
rect 191838 18663 191894 18672
rect 191852 16574 191880 18663
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 480 193260 62863
rect 194598 57352 194654 57361
rect 194598 57287 194654 57296
rect 193310 27024 193366 27033
rect 193310 26959 193366 26968
rect 193324 16574 193352 26959
rect 194612 16574 194640 57287
rect 195992 16574 196020 76026
rect 197360 74316 197412 74322
rect 197360 74258 197412 74264
rect 197372 16574 197400 74258
rect 198740 34196 198792 34202
rect 198740 34138 198792 34144
rect 193324 16546 194456 16574
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 194428 480 194456 16546
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 34138
rect 200132 16574 200160 77590
rect 213920 76968 213972 76974
rect 213920 76910 213972 76916
rect 211804 71392 211856 71398
rect 211804 71334 211856 71340
rect 209780 71324 209832 71330
rect 209780 71266 209832 71272
rect 207020 64524 207072 64530
rect 207020 64466 207072 64472
rect 201500 33856 201552 33862
rect 201500 33798 201552 33804
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 11694 201540 33798
rect 201592 27328 201644 27334
rect 201592 27270 201644 27276
rect 201500 11688 201552 11694
rect 201500 11630 201552 11636
rect 201604 6914 201632 27270
rect 204260 27260 204312 27266
rect 204260 27202 204312 27208
rect 204272 16574 204300 27202
rect 205640 17672 205692 17678
rect 205640 17614 205692 17620
rect 205652 16574 205680 17614
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 202696 11688 202748 11694
rect 202696 11630 202748 11636
rect 201512 6886 201632 6914
rect 201512 480 201540 6886
rect 202708 480 202736 11630
rect 203892 6656 203944 6662
rect 203892 6598 203944 6604
rect 203904 480 203932 6598
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 64466
rect 208400 28756 208452 28762
rect 208400 28698 208452 28704
rect 208412 16574 208440 28698
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209792 480 209820 71266
rect 209872 67176 209924 67182
rect 209872 67118 209924 67124
rect 209884 16574 209912 67118
rect 209884 16546 211016 16574
rect 210988 480 211016 16546
rect 211816 3874 211844 71334
rect 213932 16574 213960 76910
rect 215944 74724 215996 74730
rect 215944 74666 215996 74672
rect 215956 33862 215984 74666
rect 226340 74248 226392 74254
rect 226340 74190 226392 74196
rect 216680 71256 216732 71262
rect 216680 71198 216732 71204
rect 215944 33856 215996 33862
rect 215944 33798 215996 33804
rect 215300 28688 215352 28694
rect 215300 28630 215352 28636
rect 213932 16546 214512 16574
rect 213366 12200 213422 12209
rect 213366 12135 213422 12144
rect 211804 3868 211856 3874
rect 211804 3810 211856 3816
rect 212172 3800 212224 3806
rect 212172 3742 212224 3748
rect 212184 480 212212 3742
rect 213380 480 213408 12135
rect 214484 480 214512 16546
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 28630
rect 216692 16574 216720 71198
rect 223580 71188 223632 71194
rect 223580 71130 223632 71136
rect 218060 65884 218112 65890
rect 218060 65826 218112 65832
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 480 218100 65826
rect 220820 60308 220872 60314
rect 220820 60250 220872 60256
rect 219440 34128 219492 34134
rect 219440 34070 219492 34076
rect 218152 28620 218204 28626
rect 218152 28562 218204 28568
rect 218164 16574 218192 28562
rect 219452 16574 219480 34070
rect 220832 16574 220860 60250
rect 222200 28552 222252 28558
rect 222200 28494 222252 28500
rect 222212 16574 222240 28494
rect 218164 16546 219296 16574
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 219268 480 219296 16546
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222764 480 222792 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 71130
rect 225144 6588 225196 6594
rect 225144 6530 225196 6536
rect 225156 480 225184 6530
rect 226352 480 226380 74190
rect 230478 71496 230534 71505
rect 230478 71431 230534 71440
rect 226430 33824 226486 33833
rect 226430 33759 226486 33768
rect 226444 16574 226472 33759
rect 229098 28248 229154 28257
rect 229098 28183 229154 28192
rect 229112 16574 229140 28183
rect 230492 16574 230520 71431
rect 226444 16546 227576 16574
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 227548 480 227576 16546
rect 228730 6216 228786 6225
rect 228730 6151 228786 6160
rect 228744 480 228772 6151
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 77658
rect 284300 77580 284352 77586
rect 284300 77522 284352 77528
rect 252560 77512 252612 77518
rect 252560 77454 252612 77460
rect 249800 76016 249852 76022
rect 249800 75958 249852 75964
rect 242164 75608 242216 75614
rect 242164 75550 242216 75556
rect 240140 74180 240192 74186
rect 240140 74122 240192 74128
rect 234620 61872 234672 61878
rect 234620 61814 234672 61820
rect 233240 30116 233292 30122
rect 233240 30058 233292 30064
rect 233252 16574 233280 30058
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 11694 234660 61814
rect 238760 61804 238812 61810
rect 238760 61746 238812 61752
rect 234712 34060 234764 34066
rect 234712 34002 234764 34008
rect 234620 11688 234672 11694
rect 234620 11630 234672 11636
rect 234724 6914 234752 34002
rect 236000 30048 236052 30054
rect 236000 29990 236052 29996
rect 236012 16574 236040 29990
rect 238772 16574 238800 61746
rect 236012 16546 236592 16574
rect 238772 16546 239352 16574
rect 235816 11688 235868 11694
rect 235816 11630 235868 11636
rect 234632 6886 234752 6914
rect 234632 480 234660 6886
rect 235828 480 235856 11630
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 237656 14748 237708 14754
rect 237656 14690 237708 14696
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 14690
rect 239324 480 239352 16546
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 74122
rect 242176 20262 242204 75550
rect 247038 74080 247094 74089
rect 247038 74015 247094 74024
rect 244278 71360 244334 71369
rect 244278 71295 244334 71304
rect 242900 28484 242952 28490
rect 242900 28426 242952 28432
rect 241520 20256 241572 20262
rect 241520 20198 241572 20204
rect 242164 20256 242216 20262
rect 242164 20198 242216 20204
rect 241532 16574 241560 20198
rect 241532 16546 241744 16574
rect 241716 480 241744 16546
rect 242912 3874 242940 28426
rect 244292 16574 244320 71295
rect 245658 57216 245714 57225
rect 245658 57151 245714 57160
rect 245672 16574 245700 57151
rect 247052 16574 247080 74015
rect 248418 20088 248474 20097
rect 248418 20023 248474 20032
rect 244292 16546 245240 16574
rect 245672 16546 245976 16574
rect 247052 16546 247632 16574
rect 242992 7812 243044 7818
rect 242992 7754 243044 7760
rect 242900 3868 242952 3874
rect 242900 3810 242952 3816
rect 243004 3482 243032 7754
rect 244096 3868 244148 3874
rect 244096 3810 244148 3816
rect 242912 3454 243032 3482
rect 242912 480 242940 3454
rect 244108 480 244136 3810
rect 245212 480 245240 16546
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247604 480 247632 16546
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 20023
rect 249812 16574 249840 75958
rect 251180 33992 251232 33998
rect 251180 33934 251232 33940
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 3874 251220 33934
rect 251272 29980 251324 29986
rect 251272 29922 251324 29928
rect 251180 3868 251232 3874
rect 251180 3810 251232 3816
rect 251284 3482 251312 29922
rect 252572 16574 252600 77454
rect 267740 76900 267792 76906
rect 267740 76842 267792 76848
rect 260840 74112 260892 74118
rect 260840 74054 260892 74060
rect 256700 64456 256752 64462
rect 256700 64398 256752 64404
rect 253940 27192 253992 27198
rect 253940 27134 253992 27140
rect 253952 16574 253980 27134
rect 255320 20392 255372 20398
rect 255320 20334 255372 20340
rect 255332 16574 255360 20334
rect 252572 16546 253520 16574
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 252376 3868 252428 3874
rect 252376 3810 252428 3816
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3810
rect 253492 480 253520 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 64398
rect 259460 63096 259512 63102
rect 259460 63038 259512 63044
rect 258080 28416 258132 28422
rect 258080 28358 258132 28364
rect 258092 16574 258120 28358
rect 258092 16546 258304 16574
rect 258276 480 258304 16546
rect 259472 11694 259500 63038
rect 259552 33924 259604 33930
rect 259552 33866 259604 33872
rect 259460 11688 259512 11694
rect 259460 11630 259512 11636
rect 259564 6914 259592 33866
rect 260852 16574 260880 74054
rect 266358 71224 266414 71233
rect 266358 71159 266414 71168
rect 262220 35624 262272 35630
rect 262220 35566 262272 35572
rect 262232 16574 262260 35566
rect 266372 16574 266400 71159
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 266372 16546 266584 16574
rect 260656 11688 260708 11694
rect 260656 11630 260708 11636
rect 259472 6886 259592 6914
rect 259472 480 259500 6886
rect 260668 480 260696 11630
rect 261772 480 261800 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264150 8120 264206 8129
rect 264150 8055 264206 8064
rect 264164 480 264192 8055
rect 265346 7984 265402 7993
rect 265346 7919 265402 7928
rect 265360 480 265388 7919
rect 266556 480 266584 16546
rect 267752 480 267780 76842
rect 282918 73944 282974 73953
rect 282918 73879 282974 73888
rect 270500 64388 270552 64394
rect 270500 64330 270552 64336
rect 267832 29912 267884 29918
rect 267832 29854 267884 29860
rect 267844 16574 267872 29854
rect 269120 20324 269172 20330
rect 269120 20266 269172 20272
rect 269132 16574 269160 20266
rect 270512 16574 270540 64330
rect 274640 61736 274692 61742
rect 274640 61678 274692 61684
rect 273260 35556 273312 35562
rect 273260 35498 273312 35504
rect 271880 27124 271932 27130
rect 271880 27066 271932 27072
rect 271892 16574 271920 27066
rect 267844 16546 268424 16574
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 271892 16546 272472 16574
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 270052 480 270080 16546
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272444 480 272472 16546
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 35498
rect 274652 16574 274680 61678
rect 276020 35488 276072 35494
rect 276020 35430 276072 35436
rect 276032 16574 276060 35430
rect 280158 35320 280214 35329
rect 280158 35255 280214 35264
rect 278780 25764 278832 25770
rect 278780 25706 278832 25712
rect 278792 16574 278820 25706
rect 280172 16574 280200 35255
rect 282932 16574 282960 73879
rect 274652 16546 274864 16574
rect 276032 16546 276704 16574
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 282932 16546 283144 16574
rect 274836 480 274864 16546
rect 276020 6520 276072 6526
rect 276020 6462 276072 6468
rect 276032 480 276060 6462
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 16546
rect 278320 7744 278372 7750
rect 278320 7686 278372 7692
rect 278332 480 278360 7686
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 281906 9344 281962 9353
rect 281906 9279 281962 9288
rect 281920 480 281948 9279
rect 283116 480 283144 16546
rect 284312 3874 284340 77522
rect 284956 75818 284984 87586
rect 393976 78062 394004 231814
rect 395344 230444 395396 230450
rect 395344 230386 395396 230392
rect 394330 227760 394386 227769
rect 394330 227695 394386 227704
rect 394344 223106 394372 227695
rect 394332 223100 394384 223106
rect 394332 223042 394384 223048
rect 395356 210458 395384 230386
rect 395448 227798 395476 232358
rect 396460 230450 396488 675446
rect 396724 430636 396776 430642
rect 396724 430578 396776 430584
rect 396632 240032 396684 240038
rect 396632 239974 396684 239980
rect 396540 238740 396592 238746
rect 396540 238682 396592 238688
rect 396552 232422 396580 238682
rect 396540 232416 396592 232422
rect 396540 232358 396592 232364
rect 396644 231130 396672 239974
rect 396632 231124 396684 231130
rect 396632 231066 396684 231072
rect 396448 230444 396500 230450
rect 396448 230386 396500 230392
rect 395436 227792 395488 227798
rect 395436 227734 395488 227740
rect 395344 210452 395396 210458
rect 395344 210394 395396 210400
rect 393964 78056 394016 78062
rect 393964 77998 394016 78004
rect 302240 77444 302292 77450
rect 302240 77386 302292 77392
rect 288440 75948 288492 75954
rect 288440 75890 288492 75896
rect 284944 75812 284996 75818
rect 284944 75754 284996 75760
rect 284390 69864 284446 69873
rect 284390 69799 284446 69808
rect 284300 3868 284352 3874
rect 284300 3810 284352 3816
rect 284404 3482 284432 69799
rect 287060 35420 287112 35426
rect 287060 35362 287112 35368
rect 285680 29844 285732 29850
rect 285680 29786 285732 29792
rect 285692 16574 285720 29786
rect 287072 16574 287100 35362
rect 288452 16574 288480 75890
rect 296720 74044 296772 74050
rect 296720 73986 296772 73992
rect 292580 60240 292632 60246
rect 292580 60182 292632 60188
rect 289820 29776 289872 29782
rect 289820 29718 289872 29724
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 288452 16546 289032 16574
rect 285036 3868 285088 3874
rect 285036 3810 285088 3816
rect 284312 3454 284432 3482
rect 284312 480 284340 3454
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285048 354 285076 3810
rect 286612 480 286640 16546
rect 285374 354 285486 480
rect 285048 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 289004 480 289032 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 29718
rect 291384 13592 291436 13598
rect 291384 13534 291436 13540
rect 291396 480 291424 13534
rect 292592 480 292620 60182
rect 295340 54596 295392 54602
rect 295340 54538 295392 54544
rect 295352 16574 295380 54538
rect 296732 16574 296760 73986
rect 298098 69728 298154 69737
rect 298098 69663 298154 69672
rect 295352 16546 295656 16574
rect 296732 16546 297312 16574
rect 294880 16176 294932 16182
rect 294880 16118 294932 16124
rect 293684 7676 293736 7682
rect 293684 7618 293736 7624
rect 293696 480 293724 7618
rect 294892 480 294920 16118
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 297284 480 297312 16546
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 69663
rect 300858 19952 300914 19961
rect 300858 19887 300914 19896
rect 300872 16574 300900 19887
rect 302252 16574 302280 77386
rect 320180 77376 320232 77382
rect 320180 77318 320232 77324
rect 306380 76832 306432 76838
rect 306380 76774 306432 76780
rect 305000 70032 305052 70038
rect 305000 69974 305052 69980
rect 303620 31544 303672 31550
rect 303620 31486 303672 31492
rect 303632 16574 303660 31486
rect 305012 16574 305040 69974
rect 300872 16546 301544 16574
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 300766 9208 300822 9217
rect 300766 9143 300822 9152
rect 299662 9072 299718 9081
rect 299662 9007 299718 9016
rect 299676 480 299704 9007
rect 300780 480 300808 9143
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303172 480 303200 16546
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 76774
rect 311900 69964 311952 69970
rect 311900 69906 311952 69912
rect 309140 60172 309192 60178
rect 309140 60114 309192 60120
rect 307760 35352 307812 35358
rect 307760 35294 307812 35300
rect 307772 3398 307800 35294
rect 307852 31476 307904 31482
rect 307852 31418 307904 31424
rect 307864 16574 307892 31418
rect 309152 16574 309180 60114
rect 311912 16574 311940 69906
rect 318798 69592 318854 69601
rect 318798 69527 318854 69536
rect 316040 53100 316092 53106
rect 316040 53042 316092 53048
rect 307864 16546 307984 16574
rect 309152 16546 309824 16574
rect 311912 16546 312216 16574
rect 307760 3392 307812 3398
rect 307760 3334 307812 3340
rect 307956 480 307984 16546
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311440 9240 311492 9246
rect 311440 9182 311492 9188
rect 311452 480 311480 9182
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 314660 10736 314712 10742
rect 314660 10678 314712 10684
rect 313832 9172 313884 9178
rect 313832 9114 313884 9120
rect 313844 480 313872 9114
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 10678
rect 316052 3398 316080 53042
rect 316130 35184 316186 35193
rect 316130 35119 316186 35128
rect 316144 16574 316172 35119
rect 317418 25528 317474 25537
rect 317418 25463 317474 25472
rect 317432 16574 317460 25463
rect 318812 16574 318840 69527
rect 320192 16574 320220 77318
rect 396736 77081 396764 430578
rect 396816 378208 396868 378214
rect 396816 378150 396868 378156
rect 396828 77625 396856 378150
rect 397000 324352 397052 324358
rect 397000 324294 397052 324300
rect 396908 271924 396960 271930
rect 396908 271866 396960 271872
rect 396920 77858 396948 271866
rect 396908 77852 396960 77858
rect 396908 77794 396960 77800
rect 396814 77616 396870 77625
rect 396814 77551 396870 77560
rect 397012 77489 397040 324294
rect 396998 77480 397054 77489
rect 396998 77415 397054 77424
rect 397472 77217 397500 703520
rect 410524 700528 410576 700534
rect 410524 700470 410576 700476
rect 399484 700460 399536 700466
rect 399484 700402 399536 700408
rect 398104 364404 398156 364410
rect 398104 364346 398156 364352
rect 398116 142866 398144 364346
rect 398196 311908 398248 311914
rect 398196 311850 398248 311856
rect 398104 142860 398156 142866
rect 398104 142802 398156 142808
rect 398208 141506 398236 311850
rect 398288 258120 398340 258126
rect 398288 258062 398340 258068
rect 398300 141574 398328 258062
rect 399496 187678 399524 700402
rect 409144 700392 409196 700398
rect 409144 700334 409196 700340
rect 407764 700324 407816 700330
rect 407764 700266 407816 700272
rect 406384 616888 406436 616894
rect 406384 616830 406436 616836
rect 405004 563100 405056 563106
rect 405004 563042 405056 563048
rect 403624 510672 403676 510678
rect 403624 510614 403676 510620
rect 400864 456816 400916 456822
rect 400864 456758 400916 456764
rect 399484 187672 399536 187678
rect 399484 187614 399536 187620
rect 398288 141568 398340 141574
rect 398288 141510 398340 141516
rect 398196 141500 398248 141506
rect 398196 141442 398248 141448
rect 400876 95198 400904 456758
rect 403636 97986 403664 510614
rect 405016 99346 405044 563042
rect 406396 100706 406424 616830
rect 407776 103494 407804 700266
rect 409156 104854 409184 700334
rect 410536 106282 410564 700470
rect 412652 140214 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 700534 429884 703520
rect 429844 700528 429896 700534
rect 429844 700470 429896 700476
rect 446140 700466 446168 703520
rect 446128 700460 446180 700466
rect 446128 700402 446180 700408
rect 418804 404388 418856 404394
rect 418804 404330 418856 404336
rect 417424 351960 417476 351966
rect 417424 351902 417476 351908
rect 414664 298172 414716 298178
rect 414664 298114 414716 298120
rect 413284 244316 413336 244322
rect 413284 244258 413336 244264
rect 412640 140208 412692 140214
rect 412640 140150 412692 140156
rect 410524 106276 410576 106282
rect 410524 106218 410576 106224
rect 409144 104848 409196 104854
rect 409144 104790 409196 104796
rect 407764 103488 407816 103494
rect 407764 103430 407816 103436
rect 406384 100700 406436 100706
rect 406384 100642 406436 100648
rect 405004 99340 405056 99346
rect 405004 99282 405056 99288
rect 403624 97980 403676 97986
rect 403624 97922 403676 97928
rect 400864 95192 400916 95198
rect 400864 95134 400916 95140
rect 413296 89690 413324 244258
rect 414676 91050 414704 298114
rect 417436 92478 417464 351902
rect 418816 93838 418844 404330
rect 418804 93832 418856 93838
rect 418804 93774 418856 93780
rect 417424 92472 417476 92478
rect 417424 92414 417476 92420
rect 414664 91044 414716 91050
rect 414664 90986 414716 90992
rect 413284 89684 413336 89690
rect 413284 89626 413336 89632
rect 397458 77208 397514 77217
rect 397458 77143 397514 77152
rect 396722 77072 396778 77081
rect 396722 77007 396778 77016
rect 431960 76764 432012 76770
rect 431960 76706 432012 76712
rect 426440 76696 426492 76702
rect 426440 76638 426492 76644
rect 391204 75540 391256 75546
rect 391204 75482 391256 75488
rect 382280 73976 382332 73982
rect 382280 73918 382332 73924
rect 375380 71120 375432 71126
rect 375380 71062 375432 71068
rect 325700 69896 325752 69902
rect 325700 69838 325752 69844
rect 324320 64320 324372 64326
rect 324320 64262 324372 64268
rect 321560 31408 321612 31414
rect 321560 31350 321612 31356
rect 321572 16574 321600 31350
rect 322940 18964 322992 18970
rect 322940 18906 322992 18912
rect 316144 16546 316264 16574
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 316040 3392 316092 3398
rect 316040 3334 316092 3340
rect 316236 480 316264 16546
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317340 480 317368 3334
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 18906
rect 324332 3210 324360 64262
rect 324412 24472 324464 24478
rect 324412 24414 324464 24420
rect 324424 3398 324452 24414
rect 325712 16574 325740 69838
rect 332600 69828 332652 69834
rect 332600 69770 332652 69776
rect 331220 61668 331272 61674
rect 331220 61610 331272 61616
rect 329840 23180 329892 23186
rect 329840 23122 329892 23128
rect 329852 16574 329880 23122
rect 325712 16546 326384 16574
rect 329852 16546 330432 16574
rect 324412 3392 324464 3398
rect 324412 3334 324464 3340
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324332 3182 324452 3210
rect 324424 480 324452 3182
rect 325620 480 325648 3334
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328000 10668 328052 10674
rect 328000 10610 328052 10616
rect 328012 480 328040 10610
rect 329196 5228 329248 5234
rect 329196 5170 329248 5176
rect 329208 480 329236 5170
rect 330404 480 330432 16546
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 354 331260 61610
rect 332612 3398 332640 69770
rect 340880 69760 340932 69766
rect 340880 69702 340932 69708
rect 332692 65816 332744 65822
rect 332692 65758 332744 65764
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 65758
rect 338120 55888 338172 55894
rect 338120 55830 338172 55836
rect 338132 16574 338160 55830
rect 338132 16546 338712 16574
rect 334622 10432 334678 10441
rect 334622 10367 334678 10376
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 10367
rect 336278 10296 336334 10305
rect 336278 10231 336334 10240
rect 336292 480 336320 10231
rect 337474 7848 337530 7857
rect 337474 7783 337530 7792
rect 337488 480 337516 7783
rect 338684 480 338712 16546
rect 339500 13524 339552 13530
rect 339500 13466 339552 13472
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 354 339540 13466
rect 340892 3210 340920 69702
rect 367098 68232 367154 68241
rect 367098 68167 367154 68176
rect 353298 66872 353354 66881
rect 353298 66807 353354 66816
rect 347780 63028 347832 63034
rect 347780 62970 347832 62976
rect 340972 62960 341024 62966
rect 340972 62902 341024 62908
rect 340984 3398 341012 62902
rect 346400 25696 346452 25702
rect 346400 25638 346452 25644
rect 346412 16574 346440 25638
rect 347792 16574 347820 62970
rect 350538 17368 350594 17377
rect 350538 17303 350594 17312
rect 350552 16574 350580 17303
rect 353312 16574 353340 66807
rect 358820 61600 358872 61606
rect 358820 61542 358872 61548
rect 356060 60104 356112 60110
rect 356060 60046 356112 60052
rect 354680 58812 354732 58818
rect 354680 58754 354732 58760
rect 354692 16574 354720 58754
rect 356072 16574 356100 60046
rect 357440 27056 357492 27062
rect 357440 26998 357492 27004
rect 357452 16574 357480 26998
rect 358832 16574 358860 61542
rect 361580 21820 361632 21826
rect 361580 21762 361632 21768
rect 361592 16574 361620 21762
rect 367112 16574 367140 68167
rect 368480 64252 368532 64258
rect 368480 64194 368532 64200
rect 368492 16574 368520 64194
rect 374000 57384 374052 57390
rect 374000 57326 374052 57332
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 350552 16546 351224 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 356072 16546 356376 16574
rect 357452 16546 357572 16574
rect 358832 16546 359504 16574
rect 361592 16546 361896 16574
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 342904 14680 342956 14686
rect 342904 14622 342956 14628
rect 340972 3392 341024 3398
rect 340972 3334 341024 3340
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 340892 3182 341012 3210
rect 340984 480 341012 3182
rect 342180 480 342208 3334
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 14622
rect 345296 10600 345348 10606
rect 345296 10542 345348 10548
rect 344560 3800 344612 3806
rect 344560 3742 344612 3748
rect 344572 480 344600 3742
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 10542
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349158 14920 349214 14929
rect 349158 14855 349214 14864
rect 349172 1426 349200 14855
rect 349252 11960 349304 11966
rect 349252 11902 349304 11908
rect 349160 1420 349212 1426
rect 349160 1362 349212 1368
rect 349264 480 349292 11902
rect 350448 1420 350500 1426
rect 350448 1362 350500 1368
rect 350460 480 350488 1362
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352838 12064 352894 12073
rect 352838 11999 352894 12008
rect 352852 480 352880 11999
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356348 480 356376 16546
rect 357544 480 357572 16546
rect 358728 5160 358780 5166
rect 358728 5102 358780 5108
rect 358740 480 358768 5102
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 361120 11892 361172 11898
rect 361120 11834 361172 11840
rect 361132 480 361160 11834
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 365720 13456 365772 13462
rect 365720 13398 365772 13404
rect 363512 11824 363564 11830
rect 363512 11766 363564 11772
rect 363524 480 363552 11766
rect 364616 11756 364668 11762
rect 364616 11698 364668 11704
rect 364628 480 364656 11698
rect 365732 3398 365760 13398
rect 365812 9104 365864 9110
rect 365812 9046 365864 9052
rect 365720 3392 365772 3398
rect 365720 3334 365772 3340
rect 365824 480 365852 9046
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367020 480 367048 3334
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 371238 16280 371294 16289
rect 371238 16215 371294 16224
rect 370134 13016 370190 13025
rect 370134 12951 370190 12960
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 12951
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 371252 354 371280 16215
rect 372894 11928 372950 11937
rect 372894 11863 372950 11872
rect 372908 480 372936 11863
rect 374012 1170 374040 57326
rect 374092 29708 374144 29714
rect 374092 29650 374144 29656
rect 374104 3398 374132 29650
rect 375392 16574 375420 71062
rect 376760 62892 376812 62898
rect 376760 62834 376812 62840
rect 376772 16574 376800 62834
rect 379520 35284 379572 35290
rect 379520 35226 379572 35232
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374012 1142 374132 1170
rect 374104 480 374132 1142
rect 375300 480 375328 3334
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 378416 16108 378468 16114
rect 378416 16050 378468 16056
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16050
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 35226
rect 381176 13388 381228 13394
rect 381176 13330 381228 13336
rect 381188 480 381216 13330
rect 382292 3210 382320 73918
rect 390560 73908 390612 73914
rect 390560 73850 390612 73856
rect 389178 72856 389234 72865
rect 389178 72791 389234 72800
rect 382372 69692 382424 69698
rect 382372 69634 382424 69640
rect 382384 3398 382412 69634
rect 386420 35216 386472 35222
rect 386420 35158 386472 35164
rect 385040 31340 385092 31346
rect 385040 31282 385092 31288
rect 385052 16574 385080 31282
rect 386432 16574 386460 35158
rect 389192 16574 389220 72791
rect 385052 16546 386000 16574
rect 386432 16546 386736 16574
rect 389192 16546 389496 16574
rect 384304 14612 384356 14618
rect 384304 14554 384356 14560
rect 382372 3392 382424 3398
rect 382372 3334 382424 3340
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 382292 3182 382412 3210
rect 382384 480 382412 3182
rect 383580 480 383608 3334
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 14554
rect 385972 480 386000 16546
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387798 14784 387854 14793
rect 387798 14719 387854 14728
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 14719
rect 389468 480 389496 16546
rect 390572 3210 390600 73850
rect 390652 14476 390704 14482
rect 390652 14418 390704 14424
rect 390664 3398 390692 14418
rect 391216 6526 391244 75482
rect 402978 72720 403034 72729
rect 402978 72655 403034 72664
rect 396080 67108 396132 67114
rect 396080 67050 396132 67056
rect 395344 16040 395396 16046
rect 395344 15982 395396 15988
rect 392584 13320 392636 13326
rect 392584 13262 392636 13268
rect 391204 6520 391256 6526
rect 391204 6462 391256 6468
rect 390652 3392 390704 3398
rect 390652 3334 390704 3340
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 390572 3182 390692 3210
rect 390664 480 390692 3182
rect 391860 480 391888 3334
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 13262
rect 394240 6452 394292 6458
rect 394240 6394 394292 6400
rect 394252 480 394280 6394
rect 395356 480 395384 15982
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 67050
rect 401600 54528 401652 54534
rect 401600 54470 401652 54476
rect 398840 50516 398892 50522
rect 398840 50458 398892 50464
rect 398852 16574 398880 50458
rect 401612 16574 401640 54470
rect 402992 16574 403020 72655
rect 408500 65748 408552 65754
rect 408500 65690 408552 65696
rect 405738 54496 405794 54505
rect 405738 54431 405794 54440
rect 405752 16574 405780 54431
rect 408512 16574 408540 65690
rect 412640 62824 412692 62830
rect 412640 62766 412692 62772
rect 411260 18896 411312 18902
rect 411260 18838 411312 18844
rect 411272 16574 411300 18838
rect 398852 16546 398972 16574
rect 401612 16546 402560 16574
rect 402992 16546 403664 16574
rect 405752 16546 406056 16574
rect 408512 16546 409184 16574
rect 411272 16546 411944 16574
rect 397736 10532 397788 10538
rect 397736 10474 397788 10480
rect 397748 480 397776 10474
rect 398944 480 398972 16546
rect 400864 13252 400916 13258
rect 400864 13194 400916 13200
rect 400128 6384 400180 6390
rect 400128 6326 400180 6332
rect 400140 480 400168 6326
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 13194
rect 402532 480 402560 16546
rect 403636 480 403664 16546
rect 404360 14544 404412 14550
rect 404360 14486 404412 14492
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 14486
rect 406028 480 406056 16546
rect 407118 16144 407174 16153
rect 407118 16079 407174 16088
rect 407132 3398 407160 16079
rect 407210 14648 407266 14657
rect 407210 14583 407266 14592
rect 407120 3392 407172 3398
rect 407120 3334 407172 3340
rect 407224 480 407252 14583
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 408420 480 408448 3334
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410800 13184 410852 13190
rect 410800 13126 410852 13132
rect 410812 480 410840 13126
rect 411916 480 411944 16546
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 62766
rect 415400 60036 415452 60042
rect 415400 59978 415452 59984
rect 414296 5092 414348 5098
rect 414296 5034 414348 5040
rect 414308 480 414336 5034
rect 415412 3398 415440 59978
rect 422298 36544 422354 36553
rect 422298 36479 422354 36488
rect 415492 23112 415544 23118
rect 415492 23054 415544 23060
rect 415400 3392 415452 3398
rect 415400 3334 415452 3340
rect 415504 480 415532 23054
rect 418160 20188 418212 20194
rect 418160 20130 418212 20136
rect 418172 16574 418200 20130
rect 422312 16574 422340 36479
rect 425060 32632 425112 32638
rect 425060 32574 425112 32580
rect 425072 16574 425100 32574
rect 426452 16574 426480 76638
rect 431972 73166 432000 76706
rect 462332 76634 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 477512 145586 477540 702406
rect 494808 700398 494836 703520
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 504364 696992 504416 696998
rect 504364 696934 504416 696940
rect 477500 145580 477552 145586
rect 477500 145522 477552 145528
rect 462412 77308 462464 77314
rect 462412 77250 462464 77256
rect 462320 76628 462372 76634
rect 462320 76570 462372 76576
rect 431960 73160 432012 73166
rect 431960 73102 432012 73108
rect 431960 72752 432012 72758
rect 431960 72694 432012 72700
rect 430580 61532 430632 61538
rect 430580 61474 430632 61480
rect 429200 21684 429252 21690
rect 429200 21626 429252 21632
rect 418172 16546 418568 16574
rect 422312 16546 422616 16574
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 417884 9036 417936 9042
rect 417884 8978 417936 8984
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416700 480 416728 3334
rect 417896 480 417924 8978
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418540 354 418568 16546
rect 420918 16008 420974 16017
rect 420184 15972 420236 15978
rect 420918 15943 420974 15952
rect 420184 15914 420236 15920
rect 420196 480 420224 15914
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 15943
rect 422588 480 422616 16546
rect 423770 15872 423826 15881
rect 423770 15807 423826 15816
rect 423784 480 423812 15807
rect 424966 7712 425022 7721
rect 424966 7647 425022 7656
rect 424980 480 425008 7647
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428464 10464 428516 10470
rect 428464 10406 428516 10412
rect 428476 480 428504 10406
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 21626
rect 430592 16574 430620 61474
rect 430592 16546 430896 16574
rect 430868 480 430896 16546
rect 431972 1170 432000 72694
rect 438860 72684 438912 72690
rect 438860 72626 438912 72632
rect 437480 64184 437532 64190
rect 437480 64126 437532 64132
rect 434720 31272 434772 31278
rect 434720 31214 434772 31220
rect 432052 21752 432104 21758
rect 432052 21694 432104 21700
rect 432064 3398 432092 21694
rect 433340 17604 433392 17610
rect 433340 17546 433392 17552
rect 433352 16574 433380 17546
rect 434732 16574 434760 31214
rect 436100 21616 436152 21622
rect 436100 21558 436152 21564
rect 436112 16574 436140 21558
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 436112 16546 436784 16574
rect 432052 3392 432104 3398
rect 432052 3334 432104 3340
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 431972 1142 432092 1170
rect 432064 480 432092 1142
rect 433260 480 433288 3334
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 64126
rect 438872 16574 438900 72626
rect 454040 72616 454092 72622
rect 454040 72558 454092 72564
rect 441618 59936 441674 59945
rect 441618 59871 441674 59880
rect 440240 24404 440292 24410
rect 440240 24346 440292 24352
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 3210 440280 24346
rect 440332 17536 440384 17542
rect 440332 17478 440384 17484
rect 440344 3398 440372 17478
rect 441632 16574 441660 59871
rect 448520 58744 448572 58750
rect 448520 58686 448572 58692
rect 447140 26988 447192 26994
rect 447140 26930 447192 26936
rect 442998 21448 443054 21457
rect 442998 21383 443054 21392
rect 443012 16574 443040 21383
rect 447152 16574 447180 26930
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 447152 16546 447456 16574
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 440252 3182 440372 3210
rect 440344 480 440372 3182
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 446220 6316 446272 6322
rect 446220 6258 446272 6264
rect 445024 3732 445076 3738
rect 445024 3674 445076 3680
rect 445036 480 445064 3674
rect 446232 480 446260 6258
rect 447428 480 447456 16546
rect 448532 3210 448560 58686
rect 449900 20256 449952 20262
rect 449900 20198 449952 20204
rect 448612 17468 448664 17474
rect 448612 17410 448664 17416
rect 448624 3398 448652 17410
rect 449912 16574 449940 20198
rect 451280 17400 451332 17406
rect 451280 17342 451332 17348
rect 451292 16574 451320 17342
rect 452660 17332 452712 17338
rect 452660 17274 452712 17280
rect 452672 16574 452700 17274
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 450924 480 450952 16546
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 72558
rect 456800 33856 456852 33862
rect 456800 33798 456852 33804
rect 455420 17264 455472 17270
rect 455420 17206 455472 17212
rect 455432 16574 455460 17206
rect 455432 16546 455736 16574
rect 455708 480 455736 16546
rect 456812 3398 456840 33798
rect 460938 30968 460994 30977
rect 460938 30903 460994 30912
rect 458178 18592 458234 18601
rect 458178 18527 458234 18536
rect 458192 16574 458220 18527
rect 459558 17232 459614 17241
rect 459558 17167 459614 17176
rect 459572 16574 459600 17167
rect 460952 16574 460980 30903
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 456890 11792 456946 11801
rect 456890 11727 456946 11736
rect 456800 3392 456852 3398
rect 456800 3334 456852 3340
rect 456904 480 456932 11727
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462424 354 462452 77250
rect 471244 75472 471296 75478
rect 471244 75414 471296 75420
rect 469220 50448 469272 50454
rect 469220 50390 469272 50396
rect 466460 29640 466512 29646
rect 466460 29582 466512 29588
rect 463700 28348 463752 28354
rect 463700 28290 463752 28296
rect 463712 16574 463740 28290
rect 465172 18828 465224 18834
rect 465172 18770 465224 18776
rect 465184 16574 465212 18770
rect 466472 16574 466500 29582
rect 469232 16574 469260 50390
rect 470600 26920 470652 26926
rect 470600 26862 470652 26868
rect 463712 16546 464016 16574
rect 465184 16546 465856 16574
rect 466472 16546 467512 16574
rect 469232 16546 469904 16574
rect 463988 480 464016 16546
rect 465172 3664 465224 3670
rect 465172 3606 465224 3612
rect 465184 480 465212 3606
rect 462750 354 462862 480
rect 462424 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 16546
rect 467484 480 467512 16546
rect 468668 3596 468720 3602
rect 468668 3538 468720 3544
rect 468680 480 468708 3538
rect 469876 480 469904 16546
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 26862
rect 471256 3534 471284 75414
rect 478144 75404 478196 75410
rect 478144 75346 478196 75352
rect 476118 39264 476174 39273
rect 476118 39199 476174 39208
rect 473358 29608 473414 29617
rect 473358 29543 473414 29552
rect 473372 16574 473400 29543
rect 476132 16574 476160 39199
rect 473372 16546 474136 16574
rect 476132 16546 476528 16574
rect 473452 7608 473504 7614
rect 473452 7550 473504 7556
rect 471244 3528 471296 3534
rect 471244 3470 471296 3476
rect 472256 3528 472308 3534
rect 472256 3470 472308 3476
rect 472268 480 472296 3470
rect 473464 480 473492 7550
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475752 3596 475804 3602
rect 475752 3538 475804 3544
rect 475764 480 475792 3538
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478156 3194 478184 75346
rect 483020 75336 483072 75342
rect 483020 75278 483072 75284
rect 481640 58676 481692 58682
rect 481640 58618 481692 58624
rect 478234 7576 478290 7585
rect 478234 7511 478290 7520
rect 478144 3188 478196 3194
rect 478144 3130 478196 3136
rect 478248 3074 478276 7511
rect 481652 6914 481680 58618
rect 481732 50380 481784 50386
rect 481732 50322 481784 50328
rect 481744 16574 481772 50322
rect 483032 16574 483060 75278
rect 498200 75268 498252 75274
rect 498200 75210 498252 75216
rect 496818 72584 496874 72593
rect 489920 72548 489972 72554
rect 496818 72519 496874 72528
rect 489920 72490 489972 72496
rect 487160 68536 487212 68542
rect 487160 68478 487212 68484
rect 485780 32564 485832 32570
rect 485780 32506 485832 32512
rect 484400 20120 484452 20126
rect 484400 20062 484452 20068
rect 484412 16574 484440 20062
rect 485792 16574 485820 32506
rect 481744 16546 482416 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 485792 16546 486464 16574
rect 481652 6886 481772 6914
rect 480536 5024 480588 5030
rect 480536 4966 480588 4972
rect 479340 3188 479392 3194
rect 479340 3130 479392 3136
rect 478156 3046 478276 3074
rect 478156 480 478184 3046
rect 479352 480 479380 3130
rect 480548 480 480576 4966
rect 481744 480 481772 6886
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 16546
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486436 480 486464 16546
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 68478
rect 488540 20052 488592 20058
rect 488540 19994 488592 20000
rect 488552 16574 488580 19994
rect 488552 16546 488856 16574
rect 488828 480 488856 16546
rect 489932 480 489960 72490
rect 496832 16574 496860 72519
rect 496832 16546 497136 16574
rect 495438 14512 495494 14521
rect 495438 14447 495494 14456
rect 492312 8968 492364 8974
rect 492312 8910 492364 8916
rect 491116 4956 491168 4962
rect 491116 4898 491168 4904
rect 491128 480 491156 4898
rect 492324 480 492352 8910
rect 493508 6248 493560 6254
rect 493508 6190 493560 6196
rect 493520 480 493548 6190
rect 494702 3496 494758 3505
rect 494702 3431 494758 3440
rect 494716 480 494744 3431
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495452 354 495480 14447
rect 497108 480 497136 16546
rect 498212 480 498240 75210
rect 504376 74769 504404 696934
rect 527192 77353 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 542372 140146 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 544384 670744 544436 670750
rect 580172 670744 580224 670750
rect 544384 670686 544436 670692
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 542360 140140 542412 140146
rect 542360 140082 542412 140088
rect 544396 102134 544424 670686
rect 580170 670647 580226 670656
rect 579710 617536 579766 617545
rect 579710 617471 579766 617480
rect 579724 616894 579752 617471
rect 579712 616888 579764 616894
rect 579712 616830 579764 616836
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 579986 431624 580042 431633
rect 579986 431559 580042 431568
rect 580000 430642 580028 431559
rect 579988 430636 580040 430642
rect 579988 430578 580040 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580078 404968 580134 404977
rect 580078 404903 580134 404912
rect 580092 404394 580120 404903
rect 580080 404388 580132 404394
rect 580080 404330 580132 404336
rect 580078 378448 580134 378457
rect 580078 378383 580134 378392
rect 580092 378214 580120 378383
rect 580080 378208 580132 378214
rect 580080 378150 580132 378156
rect 579802 365120 579858 365129
rect 579802 365055 579858 365064
rect 579816 364410 579844 365055
rect 579804 364404 579856 364410
rect 579804 364346 579856 364352
rect 580080 351960 580132 351966
rect 580078 351928 580080 351937
rect 580132 351928 580134 351937
rect 580078 351863 580134 351872
rect 580078 325272 580134 325281
rect 580078 325207 580134 325216
rect 580092 324358 580120 325207
rect 580080 324352 580132 324358
rect 580080 324294 580132 324300
rect 580078 312080 580134 312089
rect 580078 312015 580134 312024
rect 580092 311914 580120 312015
rect 580080 311908 580132 311914
rect 580080 311850 580132 311856
rect 580078 298752 580134 298761
rect 580078 298687 580134 298696
rect 580092 298178 580120 298687
rect 580080 298172 580132 298178
rect 580080 298114 580132 298120
rect 579802 272232 579858 272241
rect 579802 272167 579858 272176
rect 579816 271930 579844 272167
rect 579804 271924 579856 271930
rect 579804 271866 579856 271872
rect 579986 258904 580042 258913
rect 579986 258839 580042 258848
rect 580000 258126 580028 258839
rect 579988 258120 580040 258126
rect 579988 258062 580040 258068
rect 579986 245576 580042 245585
rect 579986 245511 580042 245520
rect 580000 244322 580028 245511
rect 579988 244316 580040 244322
rect 579988 244258 580040 244264
rect 580078 232384 580134 232393
rect 580078 232319 580134 232328
rect 580092 231878 580120 232319
rect 580080 231872 580132 231878
rect 580080 231814 580132 231820
rect 580078 219056 580134 219065
rect 580078 218991 580134 219000
rect 580092 218074 580120 218991
rect 580080 218068 580132 218074
rect 580080 218010 580132 218016
rect 580078 205728 580134 205737
rect 580078 205663 580080 205672
rect 580132 205663 580134 205672
rect 580080 205634 580132 205640
rect 580078 192536 580134 192545
rect 580078 192471 580134 192480
rect 580092 191894 580120 192471
rect 580080 191888 580132 191894
rect 580080 191830 580132 191836
rect 580078 179208 580134 179217
rect 580078 179143 580134 179152
rect 580092 146946 580120 179143
rect 580184 171834 580212 418231
rect 580172 171828 580224 171834
rect 580172 171770 580224 171776
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580184 151842 580212 152623
rect 580172 151836 580224 151842
rect 580172 151778 580224 151784
rect 580080 146940 580132 146946
rect 580080 146882 580132 146888
rect 580276 144226 580304 683839
rect 580446 630864 580502 630873
rect 580446 630799 580502 630808
rect 580354 591016 580410 591025
rect 580354 590951 580410 590960
rect 580264 144220 580316 144226
rect 580264 144162 580316 144168
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 580184 138038 580212 139295
rect 580172 138032 580224 138038
rect 580172 137974 580224 137980
rect 580078 126032 580134 126041
rect 580078 125967 580134 125976
rect 580092 125662 580120 125967
rect 580080 125656 580132 125662
rect 580080 125598 580132 125604
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580184 111858 580212 112775
rect 580172 111852 580224 111858
rect 580172 111794 580224 111800
rect 544384 102128 544436 102134
rect 544384 102070 544436 102076
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580184 99414 580212 99447
rect 580172 99408 580224 99414
rect 580172 99350 580224 99356
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580184 85610 580212 86119
rect 580172 85604 580224 85610
rect 580172 85546 580224 85552
rect 555424 80096 555476 80102
rect 555424 80038 555476 80044
rect 527178 77344 527234 77353
rect 527178 77279 527234 77288
rect 532700 75200 532752 75206
rect 518898 75168 518954 75177
rect 532700 75142 532752 75148
rect 518898 75103 518954 75112
rect 504362 74760 504418 74769
rect 504362 74695 504418 74704
rect 514758 72448 514814 72457
rect 514758 72383 514814 72392
rect 500960 68468 501012 68474
rect 500960 68410 501012 68416
rect 499580 25628 499632 25634
rect 499580 25570 499632 25576
rect 498292 19984 498344 19990
rect 498292 19926 498344 19932
rect 498304 16574 498332 19926
rect 499592 16574 499620 25570
rect 500972 16574 501000 68410
rect 505100 68400 505152 68406
rect 505100 68342 505152 68348
rect 503720 25560 503772 25566
rect 503720 25502 503772 25508
rect 498304 16546 498976 16574
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500604 480 500632 16546
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502984 10396 503036 10402
rect 502984 10338 503036 10344
rect 502996 480 503024 10338
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 25502
rect 505112 16574 505140 68342
rect 507860 57316 507912 57322
rect 507860 57258 507912 57264
rect 506480 31204 506532 31210
rect 506480 31146 506532 31152
rect 505112 16546 505416 16574
rect 505388 480 505416 16546
rect 506492 3534 506520 31146
rect 507872 16574 507900 57258
rect 513378 21312 513434 21321
rect 513378 21247 513434 21256
rect 507872 16546 508912 16574
rect 506572 13116 506624 13122
rect 506572 13058 506624 13064
rect 506480 3528 506532 3534
rect 506480 3470 506532 3476
rect 506584 3346 506612 13058
rect 507308 3528 507360 3534
rect 507308 3470 507360 3476
rect 506492 3318 506612 3346
rect 506492 480 506520 3318
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 3470
rect 508884 480 508912 16546
rect 509608 15904 509660 15910
rect 509608 15846 509660 15852
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 15846
rect 511262 8936 511318 8945
rect 511262 8871 511318 8880
rect 511276 480 511304 8871
rect 512460 3460 512512 3466
rect 512460 3402 512512 3408
rect 512472 480 512500 3402
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513392 354 513420 21247
rect 514772 480 514800 72383
rect 516140 61464 516192 61470
rect 516140 61406 516192 61412
rect 514852 42084 514904 42090
rect 514852 42026 514904 42032
rect 514864 16574 514892 42026
rect 516152 16574 516180 61406
rect 517520 31136 517572 31142
rect 517520 31078 517572 31084
rect 517532 16574 517560 31078
rect 518912 16574 518940 75103
rect 523040 67040 523092 67046
rect 523040 66982 523092 66988
rect 521660 31068 521712 31074
rect 521660 31010 521712 31016
rect 520280 21548 520332 21554
rect 520280 21490 520332 21496
rect 514864 16546 515536 16574
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515508 354 515536 16546
rect 517164 480 517192 16546
rect 515926 354 516038 480
rect 515508 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 21490
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 31010
rect 523052 480 523080 66982
rect 529938 62792 529994 62801
rect 529938 62727 529994 62736
rect 525800 57248 525852 57254
rect 525800 57190 525852 57196
rect 524420 28280 524472 28286
rect 524420 28222 524472 28228
rect 523132 21480 523184 21486
rect 523132 21422 523184 21428
rect 523144 16574 523172 21422
rect 524432 16574 524460 28222
rect 525812 16574 525840 57190
rect 528558 32736 528614 32745
rect 528558 32671 528614 32680
rect 527180 21412 527232 21418
rect 527180 21354 527232 21360
rect 527192 16574 527220 21354
rect 523144 16546 523816 16574
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 527192 16546 527864 16574
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527836 480 527864 16546
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 32671
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 62727
rect 531318 22672 531374 22681
rect 531318 22607 531374 22616
rect 531332 480 531360 22607
rect 532712 16574 532740 75142
rect 535460 72480 535512 72486
rect 535460 72422 535512 72428
rect 534080 23044 534132 23050
rect 534080 22986 534132 22992
rect 534092 16574 534120 22986
rect 535472 16574 535500 72422
rect 536840 66972 536892 66978
rect 536840 66914 536892 66920
rect 536852 16574 536880 66914
rect 550640 66904 550692 66910
rect 550640 66846 550692 66852
rect 539600 65680 539652 65686
rect 539600 65622 539652 65628
rect 538220 22976 538272 22982
rect 538220 22918 538272 22924
rect 532712 16546 533752 16574
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 532514 4992 532570 5001
rect 532514 4927 532570 4936
rect 532528 480 532556 4927
rect 533724 480 533752 16546
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 22918
rect 539612 3534 539640 65622
rect 543740 65612 543792 65618
rect 543740 65554 543792 65560
rect 542360 32496 542412 32502
rect 542360 32438 542412 32444
rect 540980 22908 541032 22914
rect 540980 22850 541032 22856
rect 540992 16574 541020 22850
rect 542372 16574 542400 32438
rect 543752 16574 543780 65554
rect 546498 32600 546554 32609
rect 546498 32535 546554 32544
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 539692 10328 539744 10334
rect 539692 10270 539744 10276
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539704 3346 539732 10270
rect 540428 3528 540480 3534
rect 540428 3470 540480 3476
rect 539612 3318 539732 3346
rect 539612 480 539640 3318
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540440 354 540468 3470
rect 542004 480 542032 16546
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545488 4888 545540 4894
rect 545488 4830 545540 4836
rect 545500 480 545528 4830
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 32535
rect 549258 32464 549314 32473
rect 549258 32399 549314 32408
rect 547878 24304 547934 24313
rect 547878 24239 547934 24248
rect 547892 16574 547920 24239
rect 549272 16574 549300 32399
rect 550652 16574 550680 66846
rect 552020 24336 552072 24342
rect 552020 24278 552072 24284
rect 552032 16574 552060 24278
rect 553400 18760 553452 18766
rect 553400 18702 553452 18708
rect 553412 16574 553440 18702
rect 547892 16546 548656 16574
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 547878 4856 547934 4865
rect 547878 4791 547934 4800
rect 547892 480 547920 4791
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 550284 480 550312 16546
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 555436 6866 555464 80038
rect 580368 77994 580396 590951
rect 580460 141438 580488 630799
rect 580630 577688 580686 577697
rect 580630 577623 580686 577632
rect 580538 537840 580594 537849
rect 580538 537775 580594 537784
rect 580448 141432 580500 141438
rect 580448 141374 580500 141380
rect 580552 79354 580580 537775
rect 580644 138718 580672 577623
rect 580814 524512 580870 524521
rect 580814 524447 580870 524456
rect 580722 484664 580778 484673
rect 580722 484599 580778 484608
rect 580632 138712 580684 138718
rect 580632 138654 580684 138660
rect 580540 79348 580592 79354
rect 580540 79290 580592 79296
rect 580356 77988 580408 77994
rect 580356 77930 580408 77936
rect 557540 76560 557592 76566
rect 557540 76502 557592 76508
rect 556160 24268 556212 24274
rect 556160 24210 556212 24216
rect 555424 6860 555476 6866
rect 555424 6802 555476 6808
rect 554962 3360 555018 3369
rect 554962 3295 555018 3304
rect 554976 480 555004 3295
rect 556172 480 556200 24210
rect 556252 18692 556304 18698
rect 556252 18634 556304 18640
rect 556264 16574 556292 18634
rect 557552 16574 557580 76502
rect 580736 74798 580764 484599
rect 580828 179382 580856 524447
rect 580906 471472 580962 471481
rect 580906 471407 580962 471416
rect 580816 179376 580868 179382
rect 580816 179318 580868 179324
rect 580920 140078 580948 471407
rect 580908 140072 580960 140078
rect 580908 140014 580960 140020
rect 580724 74792 580776 74798
rect 580724 74734 580776 74740
rect 558920 73840 558972 73846
rect 558920 73782 558972 73788
rect 565818 73808 565874 73817
rect 558932 16574 558960 73782
rect 565818 73743 565874 73752
rect 564440 71052 564492 71058
rect 564440 70994 564492 71000
rect 563060 24200 563112 24206
rect 563060 24142 563112 24148
rect 560300 18624 560352 18630
rect 560300 18566 560352 18572
rect 560312 16574 560340 18566
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562048 6180 562100 6186
rect 562048 6122 562100 6128
rect 562060 480 562088 6122
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 24142
rect 564452 480 564480 70994
rect 564532 68332 564584 68338
rect 564532 68274 564584 68280
rect 564544 16574 564572 68274
rect 565832 16574 565860 73743
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 578238 71088 578294 71097
rect 578238 71023 578294 71032
rect 568580 65544 568632 65550
rect 568580 65486 568632 65492
rect 567198 26888 567254 26897
rect 567198 26823 567254 26832
rect 567212 16574 567240 26823
rect 568592 16574 568620 65486
rect 572720 61396 572772 61402
rect 572720 61338 572772 61344
rect 571340 32428 571392 32434
rect 571340 32370 571392 32376
rect 569960 22840 570012 22846
rect 569960 22782 570012 22788
rect 569972 16574 570000 22782
rect 564544 16546 565216 16574
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 566844 480 566872 16546
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 570340 480 570368 16546
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571352 354 571380 32370
rect 572732 480 572760 61338
rect 574100 33788 574152 33794
rect 574100 33730 574152 33736
rect 572812 24132 572864 24138
rect 572812 24074 572864 24080
rect 572824 16574 572852 24074
rect 574112 16574 574140 33730
rect 576858 24168 576914 24177
rect 576858 24103 576914 24112
rect 576872 16574 576900 24103
rect 578252 16574 578280 71023
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 582378 50280 582434 50289
rect 582378 50215 582434 50224
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 580172 22772 580224 22778
rect 580172 22714 580224 22720
rect 580184 19825 580212 22714
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 582392 16574 582420 50215
rect 572824 16546 573496 16574
rect 574112 16546 575152 16574
rect 576872 16546 576992 16574
rect 578252 16546 578648 16574
rect 582392 16546 583432 16574
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573468 354 573496 16546
rect 575124 480 575152 16546
rect 576308 4820 576360 4826
rect 576308 4762 576360 4768
rect 576320 480 576348 4762
rect 573886 354 573998 480
rect 573468 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576964 354 576992 16546
rect 578620 480 578648 16546
rect 580998 11656 581054 11665
rect 580998 11591 581054 11600
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 581012 480 581040 11591
rect 582196 6520 582248 6526
rect 582196 6462 582248 6468
rect 582208 480 582236 6462
rect 583404 480 583432 16546
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 2778 671200 2834 671256
rect 3330 579944 3386 580000
rect 3054 566888 3110 566944
rect 2962 527856 3018 527912
rect 2778 514820 2834 514856
rect 2778 514800 2780 514820
rect 2780 514800 2832 514820
rect 2832 514800 2834 514820
rect 3330 475632 3386 475688
rect 3238 462596 3294 462632
rect 3238 462576 3240 462596
rect 3240 462576 3292 462596
rect 3292 462576 3294 462596
rect 3146 423544 3202 423600
rect 3146 410488 3202 410544
rect 3238 371320 3294 371376
rect 3238 358400 3294 358456
rect 3238 319232 3294 319288
rect 3238 306176 3294 306232
rect 2778 293120 2834 293176
rect 3054 267144 3110 267200
rect 3146 254088 3202 254144
rect 2778 241032 2834 241088
rect 2962 201864 3018 201920
rect 3330 214920 3386 214976
rect 3330 188808 3386 188864
rect 3330 162868 3332 162888
rect 3332 162868 3384 162888
rect 3384 162868 3386 162888
rect 3330 162832 3386 162868
rect 3330 149776 3386 149832
rect 3606 632032 3662 632088
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3422 136740 3478 136776
rect 3422 136720 3424 136740
rect 3424 136720 3476 136740
rect 3476 136720 3478 136740
rect 3238 110608 3294 110664
rect 3330 97552 3386 97608
rect 3146 84632 3202 84688
rect 1398 73752 1454 73808
rect 2778 72392 2834 72448
rect 3698 553832 3754 553888
rect 3514 76472 3570 76528
rect 3514 71576 3570 71632
rect 3790 501744 3846 501800
rect 3698 77968 3754 78024
rect 3882 449520 3938 449576
rect 3974 397432 4030 397488
rect 4066 345344 4122 345400
rect 3974 76880 4030 76936
rect 3790 76608 3846 76664
rect 387062 643728 387118 643784
rect 6918 78104 6974 78160
rect 117318 137128 117374 137184
rect 117318 134000 117374 134056
rect 117318 132524 117374 132560
rect 117318 132504 117320 132524
rect 117320 132504 117372 132524
rect 117372 132504 117374 132524
rect 117318 131164 117374 131200
rect 117318 131144 117320 131164
rect 117320 131144 117372 131164
rect 117372 131144 117374 131164
rect 117318 129684 117320 129704
rect 117320 129684 117372 129704
rect 117372 129684 117374 129704
rect 117318 129648 117374 129684
rect 117318 128152 117374 128208
rect 117318 126792 117374 126848
rect 117318 123800 117374 123856
rect 117318 122748 117320 122768
rect 117320 122748 117372 122768
rect 117372 122748 117374 122768
rect 117318 122712 117374 122748
rect 117318 121216 117374 121272
rect 117318 119720 117374 119776
rect 117318 118224 117374 118280
rect 117318 116728 117374 116784
rect 117318 115232 117374 115288
rect 117318 113092 117320 113112
rect 117320 113092 117372 113112
rect 117372 113092 117374 113112
rect 117318 113056 117374 113092
rect 117318 111732 117320 111752
rect 117320 111732 117372 111752
rect 117372 111732 117374 111752
rect 117318 111696 117374 111732
rect 117318 110200 117374 110256
rect 117318 108840 117374 108896
rect 117318 107480 117374 107536
rect 118146 137128 118202 137184
rect 118238 135496 118294 135552
rect 118146 125432 118202 125488
rect 117870 83680 117926 83736
rect 118238 95104 118294 95160
rect 118330 91024 118386 91080
rect 118422 89664 118478 89720
rect 118606 106120 118662 106176
rect 118698 92384 118754 92440
rect 118514 88168 118570 88224
rect 118146 86808 118202 86864
rect 119066 103128 119122 103184
rect 118974 100272 119030 100328
rect 119158 98776 119214 98832
rect 138110 195916 138112 195936
rect 138112 195916 138164 195936
rect 138164 195916 138166 195936
rect 138110 195880 138166 195916
rect 140410 195880 140466 195936
rect 158902 195872 158958 195928
rect 160834 195880 160890 195936
rect 140778 195608 140834 195664
rect 157154 195608 157210 195664
rect 139398 195472 139454 195528
rect 140962 191800 141018 191856
rect 140870 191664 140926 191720
rect 140778 191528 140834 191584
rect 144550 190984 144606 191040
rect 140962 190848 141018 190904
rect 140870 190304 140926 190360
rect 140778 184184 140834 184240
rect 140962 184320 141018 184376
rect 140870 184048 140926 184104
rect 120630 136176 120686 136232
rect 119342 104760 119398 104816
rect 145838 188944 145894 189000
rect 144918 182144 144974 182200
rect 144918 181192 144974 181248
rect 145194 181192 145250 181248
rect 144642 180920 144698 180976
rect 144090 178880 144146 178936
rect 141606 178744 141662 178800
rect 141790 178744 141846 178800
rect 142066 178608 142122 178664
rect 145470 177384 145526 177440
rect 142526 172896 142582 172952
rect 158810 176432 158866 176488
rect 149242 175752 149298 175808
rect 159178 175752 159234 175808
rect 149334 175344 149390 175400
rect 159086 175344 159142 175400
rect 148690 175208 148746 175264
rect 154578 175208 154634 175264
rect 158442 172896 158498 172952
rect 154486 169496 154542 169552
rect 164238 175752 164294 175808
rect 166998 175752 167054 175808
rect 171138 157936 171194 157992
rect 179510 131688 179566 131744
rect 179602 118224 179658 118280
rect 179418 111832 179474 111888
rect 120630 101768 120686 101824
rect 119250 97280 119306 97336
rect 118882 93744 118938 93800
rect 118790 85312 118846 85368
rect 120630 81504 120686 81560
rect 118514 80144 118570 80200
rect 118422 78648 118478 78704
rect 20718 73888 20774 73944
rect 3606 58520 3662 58576
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3514 6432 3570 6488
rect 4066 3304 4122 3360
rect 20626 6160 20682 6216
rect 35898 71032 35954 71088
rect 38382 8880 38438 8936
rect 41878 9016 41934 9072
rect 40682 6296 40738 6352
rect 53838 72528 53894 72584
rect 57978 72664 58034 72720
rect 57242 9152 57298 9208
rect 56046 7520 56102 7576
rect 74998 11600 75054 11656
rect 73802 6432 73858 6488
rect 89718 71168 89774 71224
rect 88154 6568 88210 6624
rect 92478 10240 92534 10296
rect 91558 7656 91614 7712
rect 109314 9288 109370 9344
rect 111798 74024 111854 74080
rect 121366 73888 121422 73944
rect 110510 10376 110566 10432
rect 114006 10512 114062 10568
rect 123758 77832 123814 77888
rect 124770 77152 124826 77208
rect 125322 75112 125378 75168
rect 125506 73752 125562 73808
rect 126012 77832 126068 77888
rect 126288 77832 126344 77888
rect 126242 77696 126298 77752
rect 125690 72392 125746 72448
rect 126242 71848 126298 71904
rect 127576 77832 127632 77888
rect 128036 77832 128092 77888
rect 126610 75384 126666 75440
rect 126610 71304 126666 71360
rect 127530 77696 127586 77752
rect 127254 76744 127310 76800
rect 127070 76336 127126 76392
rect 128450 76744 128506 76800
rect 128450 76336 128506 76392
rect 128542 75792 128598 75848
rect 128174 3304 128230 3360
rect 129048 77832 129104 77888
rect 128818 76064 128874 76120
rect 128726 75520 128782 75576
rect 128634 74160 128690 74216
rect 129278 77152 129334 77208
rect 129876 77832 129932 77888
rect 129738 76336 129794 76392
rect 129830 72664 129886 72720
rect 130014 76336 130070 76392
rect 130520 77832 130576 77888
rect 130566 75656 130622 75712
rect 130382 71712 130438 71768
rect 130842 77696 130898 77752
rect 131716 77832 131772 77888
rect 131992 77832 132048 77888
rect 131118 74840 131174 74896
rect 131210 74704 131266 74760
rect 131394 77424 131450 77480
rect 131302 74568 131358 74624
rect 131946 77696 132002 77752
rect 132360 77832 132416 77888
rect 132544 77832 132600 77888
rect 132912 77832 132968 77888
rect 133188 77832 133244 77888
rect 133648 77832 133704 77888
rect 133832 77832 133888 77888
rect 132038 77424 132094 77480
rect 132498 77152 132554 77208
rect 132590 76336 132646 76392
rect 132682 74976 132738 75032
rect 132866 76200 132922 76256
rect 132774 74432 132830 74488
rect 132590 74160 132646 74216
rect 132498 71168 132554 71224
rect 133510 77696 133566 77752
rect 133786 77696 133842 77752
rect 134384 77832 134440 77888
rect 134154 77308 134210 77344
rect 134154 77288 134156 77308
rect 134156 77288 134208 77308
rect 134208 77288 134210 77308
rect 134752 77832 134808 77888
rect 134338 76336 134394 76392
rect 134062 74976 134118 75032
rect 134154 74296 134210 74352
rect 134522 77696 134578 77752
rect 135396 77730 135452 77786
rect 136040 77832 136096 77888
rect 136224 77832 136280 77888
rect 136408 77832 136464 77888
rect 136684 77832 136740 77888
rect 136868 77832 136924 77888
rect 135442 74976 135498 75032
rect 136178 77696 136234 77752
rect 136086 74976 136142 75032
rect 136822 77696 136878 77752
rect 136546 77424 136602 77480
rect 137420 77832 137476 77888
rect 137374 77696 137430 77752
rect 137282 73344 137338 73400
rect 137926 74976 137982 75032
rect 138110 77424 138166 77480
rect 138018 73752 138074 73808
rect 138386 77424 138442 77480
rect 138294 73888 138350 73944
rect 138846 77696 138902 77752
rect 138570 77424 138626 77480
rect 138570 77324 138572 77344
rect 138572 77324 138624 77344
rect 138624 77324 138626 77344
rect 138570 77288 138626 77324
rect 139030 76336 139086 76392
rect 138938 74976 138994 75032
rect 139306 76336 139362 76392
rect 139122 72936 139178 72992
rect 139904 77696 139960 77752
rect 139582 77152 139638 77208
rect 139858 74976 139914 75032
rect 140502 77560 140558 77616
rect 140502 77424 140558 77480
rect 140594 74976 140650 75032
rect 140686 74840 140742 74896
rect 142066 74568 142122 74624
rect 141974 74160 142030 74216
rect 143124 77696 143180 77752
rect 143078 77560 143134 77616
rect 143584 77696 143640 77752
rect 143262 74840 143318 74896
rect 143170 74704 143226 74760
rect 143446 74704 143502 74760
rect 143354 74568 143410 74624
rect 143630 77016 143686 77072
rect 144550 77696 144606 77752
rect 144872 77832 144928 77888
rect 144550 77288 144606 77344
rect 145608 77732 145610 77752
rect 145610 77732 145662 77752
rect 145662 77732 145664 77752
rect 145608 77696 145664 77732
rect 144642 74976 144698 75032
rect 144918 75112 144974 75168
rect 144734 74024 144790 74080
rect 145102 74976 145158 75032
rect 145470 77444 145526 77480
rect 145470 77424 145472 77444
rect 145472 77424 145524 77444
rect 145524 77424 145526 77444
rect 145838 77696 145894 77752
rect 145838 77580 145894 77616
rect 145838 77560 145840 77580
rect 145840 77560 145892 77580
rect 145892 77560 145894 77580
rect 145930 77424 145986 77480
rect 145838 76200 145894 76256
rect 146252 77696 146308 77752
rect 146114 76336 146170 76392
rect 146298 77560 146354 77616
rect 146666 77560 146722 77616
rect 146206 71168 146262 71224
rect 146574 77424 146630 77480
rect 146896 77696 146952 77752
rect 147034 77560 147090 77616
rect 147310 76744 147366 76800
rect 147586 73888 147642 73944
rect 147402 73480 147458 73536
rect 148690 77696 148746 77752
rect 148598 77560 148654 77616
rect 148874 75656 148930 75712
rect 148782 74976 148838 75032
rect 149058 77308 149114 77344
rect 149058 77288 149060 77308
rect 149060 77288 149112 77308
rect 149112 77288 149114 77308
rect 148966 74568 149022 74624
rect 149058 69672 149114 69728
rect 149334 77424 149390 77480
rect 149978 75656 150034 75712
rect 150162 76200 150218 76256
rect 150162 69808 150218 69864
rect 150438 77288 150494 77344
rect 150346 69536 150402 69592
rect 150944 77832 151000 77888
rect 151680 77832 151736 77888
rect 151082 77696 151138 77752
rect 151174 75792 151230 75848
rect 152048 77832 152104 77888
rect 152324 77832 152380 77888
rect 152600 77832 152656 77888
rect 152784 77832 152840 77888
rect 151542 75656 151598 75712
rect 151542 75520 151598 75576
rect 151726 72800 151782 72856
rect 152738 77696 152794 77752
rect 152278 75792 152334 75848
rect 152278 75520 152334 75576
rect 153428 77832 153484 77888
rect 152830 76064 152886 76120
rect 152830 75948 152886 75984
rect 152830 75928 152832 75948
rect 152832 75928 152884 75948
rect 152884 75928 152886 75948
rect 153198 77580 153254 77616
rect 153198 77560 153200 77580
rect 153200 77560 153252 77580
rect 153252 77560 153254 77580
rect 153198 76744 153254 76800
rect 152922 75656 152978 75712
rect 153290 75248 153346 75304
rect 153704 77832 153760 77888
rect 154072 77832 154128 77888
rect 153658 76200 153714 76256
rect 153842 77152 153898 77208
rect 154210 77560 154266 77616
rect 154118 76744 154174 76800
rect 154026 76336 154082 76392
rect 154026 74976 154082 75032
rect 154210 75792 154266 75848
rect 154532 77832 154588 77888
rect 154302 75656 154358 75712
rect 154486 75520 154542 75576
rect 154992 77832 155048 77888
rect 154854 77016 154910 77072
rect 154854 75792 154910 75848
rect 154762 75520 154818 75576
rect 155912 77866 155968 77922
rect 155314 77424 155370 77480
rect 155682 76744 155738 76800
rect 156188 77866 156244 77922
rect 155958 77560 156014 77616
rect 155774 72800 155830 72856
rect 156050 75792 156106 75848
rect 156050 75656 156106 75712
rect 156326 77016 156382 77072
rect 156694 77560 156750 77616
rect 157108 77866 157164 77922
rect 157384 77832 157440 77888
rect 157752 77866 157808 77922
rect 157246 77696 157302 77752
rect 157430 77696 157486 77752
rect 157062 75384 157118 75440
rect 157430 75656 157486 75712
rect 157154 72664 157210 72720
rect 157890 77696 157946 77752
rect 158488 77832 158544 77888
rect 158672 77832 158728 77888
rect 158258 77560 158314 77616
rect 158534 77696 158590 77752
rect 159224 77696 159280 77752
rect 159730 77696 159786 77752
rect 158350 76064 158406 76120
rect 158534 77016 158590 77072
rect 158902 75112 158958 75168
rect 159546 77424 159602 77480
rect 159546 77016 159602 77072
rect 159638 74568 159694 74624
rect 160006 74976 160062 75032
rect 160696 77696 160752 77752
rect 158902 16360 158958 16416
rect 160466 77560 160522 77616
rect 160742 75520 160798 75576
rect 160466 74432 160522 74488
rect 161018 77662 161074 77718
rect 161478 77560 161534 77616
rect 161386 75928 161442 75984
rect 161294 75520 161350 75576
rect 162352 77832 162408 77888
rect 162720 77866 162776 77922
rect 163088 77832 163144 77888
rect 161754 76064 161810 76120
rect 162582 77696 162638 77752
rect 163456 77832 163512 77888
rect 164008 77866 164064 77922
rect 162674 76780 162676 76800
rect 162676 76780 162728 76800
rect 162728 76780 162730 76800
rect 162674 76744 162730 76780
rect 162582 76336 162638 76392
rect 162490 76200 162546 76256
rect 162950 77460 162952 77480
rect 162952 77460 163004 77480
rect 163004 77460 163006 77480
rect 162950 77424 163006 77460
rect 163042 77152 163098 77208
rect 164192 77832 164248 77888
rect 163410 75928 163466 75984
rect 163594 75520 163650 75576
rect 164054 76200 164110 76256
rect 163870 73072 163926 73128
rect 160098 4800 160154 4856
rect 161294 3304 161350 3360
rect 164238 77424 164294 77480
rect 164422 77560 164478 77616
rect 164836 77866 164892 77922
rect 165296 77832 165352 77888
rect 164514 75248 164570 75304
rect 164882 77424 164938 77480
rect 164974 75112 165030 75168
rect 165480 77866 165536 77922
rect 165342 77016 165398 77072
rect 165526 76780 165528 76800
rect 165528 76780 165580 76800
rect 165580 76780 165582 76800
rect 165526 76744 165582 76780
rect 165342 72528 165398 72584
rect 165848 77832 165904 77888
rect 165894 77424 165950 77480
rect 165710 73480 165766 73536
rect 166170 77560 166226 77616
rect 166078 75112 166134 75168
rect 166952 77832 167008 77888
rect 166078 70896 166134 70952
rect 166446 77424 166502 77480
rect 166630 77016 166686 77072
rect 167228 77832 167284 77888
rect 166722 76200 166778 76256
rect 166722 76064 166778 76120
rect 166906 77560 166962 77616
rect 166998 77424 167054 77480
rect 166906 77016 166962 77072
rect 166906 76744 166962 76800
rect 167090 77152 167146 77208
rect 167090 77016 167146 77072
rect 166906 75792 166962 75848
rect 167504 77866 167560 77922
rect 168056 77832 168112 77888
rect 167550 77288 167606 77344
rect 167274 76200 167330 76256
rect 166998 74296 167054 74352
rect 166998 74160 167054 74216
rect 166998 73752 167054 73808
rect 167550 76200 167606 76256
rect 168608 77832 168664 77888
rect 168010 77152 168066 77208
rect 168102 76744 168158 76800
rect 167826 74704 167882 74760
rect 169160 77832 169216 77888
rect 168378 77560 168434 77616
rect 168562 77560 168618 77616
rect 168286 76336 168342 76392
rect 168194 75792 168250 75848
rect 168470 76336 168526 76392
rect 169344 77832 169400 77888
rect 169528 77832 169584 77888
rect 169114 77560 169170 77616
rect 169298 77560 169354 77616
rect 169482 77560 169538 77616
rect 169390 74296 169446 74352
rect 169666 76336 169722 76392
rect 170080 77832 170136 77888
rect 170264 77866 170320 77922
rect 169574 73616 169630 73672
rect 170448 77696 170504 77752
rect 170632 77832 170688 77888
rect 170310 75656 170366 75712
rect 170586 75656 170642 75712
rect 170218 74976 170274 75032
rect 171000 77832 171056 77888
rect 171644 77832 171700 77888
rect 170770 74704 170826 74760
rect 170494 72392 170550 72448
rect 171138 77288 171194 77344
rect 171506 77288 171562 77344
rect 172196 77832 172252 77888
rect 172380 77866 172436 77922
rect 171598 77016 171654 77072
rect 171782 76744 171838 76800
rect 170862 73208 170918 73264
rect 171690 74568 171746 74624
rect 171966 77424 172022 77480
rect 172150 77424 172206 77480
rect 172058 77288 172114 77344
rect 172748 77832 172804 77888
rect 172426 77424 172482 77480
rect 172334 75384 172390 75440
rect 171966 73752 172022 73808
rect 172150 69944 172206 70000
rect 172978 77288 173034 77344
rect 173484 77832 173540 77888
rect 173852 77832 173908 77888
rect 173346 77560 173402 77616
rect 173622 77596 173624 77616
rect 173624 77596 173676 77616
rect 173676 77596 173678 77616
rect 173622 77560 173678 77596
rect 173530 76880 173586 76936
rect 173438 76608 173494 76664
rect 173162 76472 173218 76528
rect 173070 76336 173126 76392
rect 172978 76200 173034 76256
rect 172518 65456 172574 65512
rect 173254 70352 173310 70408
rect 173898 72936 173954 72992
rect 174358 77832 174414 77888
rect 178958 78512 179014 78568
rect 174818 78376 174874 78432
rect 174542 75520 174598 75576
rect 175646 77696 175702 77752
rect 175830 77716 175886 77752
rect 180890 135360 180946 135416
rect 180798 122712 180854 122768
rect 180154 78376 180210 78432
rect 176290 77832 176346 77888
rect 175830 77696 175832 77716
rect 175832 77696 175884 77716
rect 175884 77696 175886 77716
rect 175830 77580 175886 77616
rect 175830 77560 175832 77580
rect 175832 77560 175884 77580
rect 175884 77560 175886 77580
rect 175830 77424 175886 77480
rect 178406 77152 178462 77208
rect 176290 77016 176346 77072
rect 176198 76064 176254 76120
rect 175646 74704 175702 74760
rect 175278 63008 175334 63064
rect 176658 33904 176714 33960
rect 180982 129648 181038 129704
rect 181074 115232 181130 115288
rect 182178 133184 182234 133240
rect 182362 128288 182418 128344
rect 182270 124072 182326 124128
rect 181166 113056 181222 113112
rect 182730 125296 182786 125352
rect 183006 133864 183062 133920
rect 182914 126928 182970 126984
rect 182822 121216 182878 121272
rect 182638 119720 182694 119776
rect 182546 116728 182602 116784
rect 182454 110336 182510 110392
rect 182822 100136 182878 100192
rect 182822 98776 182878 98832
rect 182270 89392 182326 89448
rect 182178 85040 182234 85096
rect 182270 83816 182326 83872
rect 182822 81504 182878 81560
rect 181442 77832 181498 77888
rect 181442 77424 181498 77480
rect 183466 108840 183522 108896
rect 183466 107344 183522 107400
rect 183466 105984 183522 106040
rect 183466 104488 183522 104544
rect 183466 102992 183522 103048
rect 183466 101632 183522 101688
rect 183466 97280 183522 97336
rect 183466 95140 183468 95160
rect 183468 95140 183520 95160
rect 183520 95140 183522 95160
rect 183466 95104 183522 95140
rect 183466 93780 183468 93800
rect 183468 93780 183520 93800
rect 183520 93780 183522 93800
rect 183466 93744 183522 93780
rect 183466 92248 183522 92304
rect 183466 90888 183522 90944
rect 183466 88032 183522 88088
rect 183466 86536 183522 86592
rect 183466 80144 183522 80200
rect 193218 62872 193274 62928
rect 191838 18672 191894 18728
rect 194598 57296 194654 57352
rect 193310 26968 193366 27024
rect 213366 12144 213422 12200
rect 230478 71440 230534 71496
rect 226430 33768 226486 33824
rect 229098 28192 229154 28248
rect 228730 6160 228786 6216
rect 247038 74024 247094 74080
rect 244278 71304 244334 71360
rect 245658 57160 245714 57216
rect 248418 20032 248474 20088
rect 266358 71168 266414 71224
rect 264150 8064 264206 8120
rect 265346 7928 265402 7984
rect 282918 73888 282974 73944
rect 280158 35264 280214 35320
rect 281906 9288 281962 9344
rect 394330 227704 394386 227760
rect 284390 69808 284446 69864
rect 298098 69672 298154 69728
rect 300858 19896 300914 19952
rect 300766 9152 300822 9208
rect 299662 9016 299718 9072
rect 318798 69536 318854 69592
rect 316130 35128 316186 35184
rect 317418 25472 317474 25528
rect 396814 77560 396870 77616
rect 396998 77424 397054 77480
rect 397458 77152 397514 77208
rect 396722 77016 396778 77072
rect 334622 10376 334678 10432
rect 336278 10240 336334 10296
rect 337474 7792 337530 7848
rect 367098 68176 367154 68232
rect 353298 66816 353354 66872
rect 350538 17312 350594 17368
rect 349158 14864 349214 14920
rect 352838 12008 352894 12064
rect 371238 16224 371294 16280
rect 370134 12960 370190 13016
rect 372894 11872 372950 11928
rect 389178 72800 389234 72856
rect 387798 14728 387854 14784
rect 402978 72664 403034 72720
rect 405738 54440 405794 54496
rect 407118 16088 407174 16144
rect 407210 14592 407266 14648
rect 422298 36488 422354 36544
rect 420918 15952 420974 16008
rect 423770 15816 423826 15872
rect 424966 7656 425022 7712
rect 441618 59880 441674 59936
rect 442998 21392 443054 21448
rect 460938 30912 460994 30968
rect 458178 18536 458234 18592
rect 459558 17176 459614 17232
rect 456890 11736 456946 11792
rect 476118 39208 476174 39264
rect 473358 29552 473414 29608
rect 478234 7520 478290 7576
rect 496818 72528 496874 72584
rect 495438 14456 495494 14512
rect 494702 3440 494758 3496
rect 580170 697176 580226 697232
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 579710 617480 579766 617536
rect 580170 564304 580226 564360
rect 580170 511264 580226 511320
rect 580170 458088 580226 458144
rect 579986 431568 580042 431624
rect 580170 418240 580226 418296
rect 580078 404912 580134 404968
rect 580078 378392 580134 378448
rect 579802 365064 579858 365120
rect 580078 351908 580080 351928
rect 580080 351908 580132 351928
rect 580132 351908 580134 351928
rect 580078 351872 580134 351908
rect 580078 325216 580134 325272
rect 580078 312024 580134 312080
rect 580078 298696 580134 298752
rect 579802 272176 579858 272232
rect 579986 258848 580042 258904
rect 579986 245520 580042 245576
rect 580078 232328 580134 232384
rect 580078 219000 580134 219056
rect 580078 205692 580134 205728
rect 580078 205672 580080 205692
rect 580080 205672 580132 205692
rect 580132 205672 580134 205692
rect 580078 192480 580134 192536
rect 580078 179152 580134 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580446 630808 580502 630864
rect 580354 590960 580410 591016
rect 580170 139304 580226 139360
rect 580078 125976 580134 126032
rect 580170 112784 580226 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 527178 77288 527234 77344
rect 518898 75112 518954 75168
rect 504362 74704 504418 74760
rect 514758 72392 514814 72448
rect 513378 21256 513434 21312
rect 511262 8880 511318 8936
rect 529938 62736 529994 62792
rect 528558 32680 528614 32736
rect 531318 22616 531374 22672
rect 532514 4936 532570 4992
rect 546498 32544 546554 32600
rect 549258 32408 549314 32464
rect 547878 24248 547934 24304
rect 547878 4800 547934 4856
rect 580630 577632 580686 577688
rect 580538 537784 580594 537840
rect 580814 524456 580870 524512
rect 580722 484608 580778 484664
rect 554962 3304 555018 3360
rect 580906 471416 580962 471472
rect 565818 73752 565874 73808
rect 580170 72936 580226 72992
rect 578238 71032 578294 71088
rect 567198 26832 567254 26888
rect 576858 24112 576914 24168
rect 580170 59608 580226 59664
rect 582378 50224 582434 50280
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 19760 580226 19816
rect 580998 11600 581054 11656
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 2773 671258 2839 671261
rect -960 671256 2839 671258
rect -960 671200 2778 671256
rect 2834 671200 2839 671256
rect -960 671198 2839 671200
rect -960 671108 480 671198
rect 2773 671195 2839 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3366 658202 3372 658204
rect -960 658142 3372 658202
rect -960 658052 480 658142
rect 3366 658140 3372 658142
rect 3436 658140 3442 658204
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 644058 584960 644148
rect 583342 643998 584960 644058
rect 583342 643922 583402 643998
rect 583520 643922 584960 643998
rect 583342 643908 584960 643922
rect 583342 643862 583586 643908
rect 387057 643786 387123 643789
rect 396758 643786 396764 643788
rect 387057 643784 396764 643786
rect 387057 643728 387062 643784
rect 387118 643728 396764 643784
rect 387057 643726 396764 643728
rect 387057 643723 387123 643726
rect 396758 643724 396764 643726
rect 396828 643724 396834 643788
rect 396574 643180 396580 643244
rect 396644 643242 396650 643244
rect 583526 643242 583586 643862
rect 396644 643182 583586 643242
rect 396644 643180 396650 643182
rect -960 632090 480 632180
rect 3601 632090 3667 632093
rect -960 632088 3667 632090
rect -960 632032 3606 632088
rect 3662 632032 3667 632088
rect -960 632030 3667 632032
rect -960 631940 480 632030
rect 3601 632027 3667 632030
rect 580441 630866 580507 630869
rect 583520 630866 584960 630956
rect 580441 630864 584960 630866
rect 580441 630808 580446 630864
rect 580502 630808 584960 630864
rect 580441 630806 584960 630808
rect 580441 630803 580507 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 579705 617538 579771 617541
rect 583520 617538 584960 617628
rect 579705 617536 584960 617538
rect 579705 617480 579710 617536
rect 579766 617480 584960 617536
rect 579705 617478 584960 617480
rect 579705 617475 579771 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580349 591018 580415 591021
rect 583520 591018 584960 591108
rect 580349 591016 584960 591018
rect 580349 590960 580354 591016
rect 580410 590960 584960 591016
rect 580349 590958 584960 590960
rect 580349 590955 580415 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580625 577690 580691 577693
rect 583520 577690 584960 577780
rect 580625 577688 584960 577690
rect 580625 577632 580630 577688
rect 580686 577632 584960 577688
rect 580625 577630 584960 577632
rect 580625 577627 580691 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3049 566946 3115 566949
rect -960 566944 3115 566946
rect -960 566888 3054 566944
rect 3110 566888 3115 566944
rect -960 566886 3115 566888
rect -960 566796 480 566886
rect 3049 566883 3115 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3693 553890 3759 553893
rect -960 553888 3759 553890
rect -960 553832 3698 553888
rect 3754 553832 3759 553888
rect -960 553830 3759 553832
rect -960 553740 480 553830
rect 3693 553827 3759 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580533 537842 580599 537845
rect 583520 537842 584960 537932
rect 580533 537840 584960 537842
rect 580533 537784 580538 537840
rect 580594 537784 584960 537840
rect 580533 537782 584960 537784
rect 580533 537779 580599 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580809 524514 580875 524517
rect 583520 524514 584960 524604
rect 580809 524512 584960 524514
rect 580809 524456 580814 524512
rect 580870 524456 584960 524512
rect 580809 524454 584960 524456
rect 580809 524451 580875 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 2773 514858 2839 514861
rect -960 514856 2839 514858
rect -960 514800 2778 514856
rect 2834 514800 2839 514856
rect -960 514798 2839 514800
rect -960 514708 480 514798
rect 2773 514795 2839 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3785 501802 3851 501805
rect -960 501800 3851 501802
rect -960 501744 3790 501800
rect 3846 501744 3851 501800
rect -960 501742 3851 501744
rect -960 501652 480 501742
rect 3785 501739 3851 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580717 484666 580783 484669
rect 583520 484666 584960 484756
rect 580717 484664 584960 484666
rect 580717 484608 580722 484664
rect 580778 484608 584960 484664
rect 580717 484606 584960 484608
rect 580717 484603 580783 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 580901 471474 580967 471477
rect 583520 471474 584960 471564
rect 580901 471472 584960 471474
rect 580901 471416 580906 471472
rect 580962 471416 584960 471472
rect 580901 471414 584960 471416
rect 580901 471411 580967 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3877 449578 3943 449581
rect -960 449576 3943 449578
rect -960 449520 3882 449576
rect 3938 449520 3943 449576
rect -960 449518 3943 449520
rect -960 449428 480 449518
rect 3877 449515 3943 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 579981 431626 580047 431629
rect 583520 431626 584960 431716
rect 579981 431624 584960 431626
rect 579981 431568 579986 431624
rect 580042 431568 584960 431624
rect 579981 431566 584960 431568
rect 579981 431563 580047 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3141 423602 3207 423605
rect -960 423600 3207 423602
rect -960 423544 3146 423600
rect 3202 423544 3207 423600
rect -960 423542 3207 423544
rect -960 423452 480 423542
rect 3141 423539 3207 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 580073 404970 580139 404973
rect 583520 404970 584960 405060
rect 580073 404968 584960 404970
rect 580073 404912 580078 404968
rect 580134 404912 584960 404968
rect 580073 404910 584960 404912
rect 580073 404907 580139 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3969 397490 4035 397493
rect -960 397488 4035 397490
rect -960 397432 3974 397488
rect 4030 397432 4035 397488
rect -960 397430 4035 397432
rect -960 397340 480 397430
rect 3969 397427 4035 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580073 378450 580139 378453
rect 583520 378450 584960 378540
rect 580073 378448 584960 378450
rect 580073 378392 580078 378448
rect 580134 378392 584960 378448
rect 580073 378390 584960 378392
rect 580073 378387 580139 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3233 371378 3299 371381
rect -960 371376 3299 371378
rect -960 371320 3238 371376
rect 3294 371320 3299 371376
rect -960 371318 3299 371320
rect -960 371228 480 371318
rect 3233 371315 3299 371318
rect 579797 365122 579863 365125
rect 583520 365122 584960 365212
rect 579797 365120 584960 365122
rect 579797 365064 579802 365120
rect 579858 365064 584960 365120
rect 579797 365062 584960 365064
rect 579797 365059 579863 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3233 358458 3299 358461
rect -960 358456 3299 358458
rect -960 358400 3238 358456
rect 3294 358400 3299 358456
rect -960 358398 3299 358400
rect -960 358308 480 358398
rect 3233 358395 3299 358398
rect 580073 351930 580139 351933
rect 583520 351930 584960 352020
rect 580073 351928 584960 351930
rect 580073 351872 580078 351928
rect 580134 351872 584960 351928
rect 580073 351870 584960 351872
rect 580073 351867 580139 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 4061 345402 4127 345405
rect -960 345400 4127 345402
rect -960 345344 4066 345400
rect 4122 345344 4127 345400
rect -960 345342 4127 345344
rect -960 345252 480 345342
rect 4061 345339 4127 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580073 325274 580139 325277
rect 583520 325274 584960 325364
rect 580073 325272 584960 325274
rect 580073 325216 580078 325272
rect 580134 325216 584960 325272
rect 580073 325214 584960 325216
rect 580073 325211 580139 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3233 319290 3299 319293
rect -960 319288 3299 319290
rect -960 319232 3238 319288
rect 3294 319232 3299 319288
rect -960 319230 3299 319232
rect -960 319140 480 319230
rect 3233 319227 3299 319230
rect 580073 312082 580139 312085
rect 583520 312082 584960 312172
rect 580073 312080 584960 312082
rect 580073 312024 580078 312080
rect 580134 312024 584960 312080
rect 580073 312022 584960 312024
rect 580073 312019 580139 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 580073 298754 580139 298757
rect 583520 298754 584960 298844
rect 580073 298752 584960 298754
rect 580073 298696 580078 298752
rect 580134 298696 584960 298752
rect 580073 298694 584960 298696
rect 580073 298691 580139 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 2773 293178 2839 293181
rect -960 293176 2839 293178
rect -960 293120 2778 293176
rect 2834 293120 2839 293176
rect -960 293118 2839 293120
rect -960 293028 480 293118
rect 2773 293115 2839 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579797 272234 579863 272237
rect 583520 272234 584960 272324
rect 579797 272232 584960 272234
rect 579797 272176 579802 272232
rect 579858 272176 584960 272232
rect 579797 272174 584960 272176
rect 579797 272171 579863 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 579981 258906 580047 258909
rect 583520 258906 584960 258996
rect 579981 258904 584960 258906
rect 579981 258848 579986 258904
rect 580042 258848 584960 258904
rect 579981 258846 584960 258848
rect 579981 258843 580047 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 579981 245578 580047 245581
rect 583520 245578 584960 245668
rect 579981 245576 584960 245578
rect 579981 245520 579986 245576
rect 580042 245520 584960 245576
rect 579981 245518 584960 245520
rect 579981 245515 580047 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 580073 232386 580139 232389
rect 583520 232386 584960 232476
rect 580073 232384 584960 232386
rect 580073 232328 580078 232384
rect 580134 232328 584960 232384
rect 580073 232326 584960 232328
rect 580073 232323 580139 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 394325 227762 394391 227765
rect 396758 227762 396764 227764
rect 394325 227760 396764 227762
rect 394325 227704 394330 227760
rect 394386 227704 396764 227760
rect 394325 227702 396764 227704
rect 394325 227699 394391 227702
rect 396758 227700 396764 227702
rect 396828 227700 396834 227764
rect 580073 219058 580139 219061
rect 583520 219058 584960 219148
rect 580073 219056 584960 219058
rect 580073 219000 580078 219056
rect 580134 219000 584960 219056
rect 580073 218998 584960 219000
rect 580073 218995 580139 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 580073 205730 580139 205733
rect 583520 205730 584960 205820
rect 580073 205728 584960 205730
rect 580073 205672 580078 205728
rect 580134 205672 584960 205728
rect 580073 205670 584960 205672
rect 580073 205667 580139 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 2957 201922 3023 201925
rect -960 201920 3023 201922
rect -960 201864 2962 201920
rect 3018 201864 3023 201920
rect -960 201862 3023 201864
rect -960 201772 480 201862
rect 2957 201859 3023 201862
rect 138105 195938 138171 195941
rect 140405 195938 140471 195941
rect 160829 195938 160895 195941
rect 138105 195936 140471 195938
rect 138105 195880 138110 195936
rect 138166 195880 140410 195936
rect 140466 195880 140471 195936
rect 138105 195878 140471 195880
rect 138105 195875 138171 195878
rect 140405 195875 140471 195878
rect 158854 195936 160895 195938
rect 158854 195928 160834 195936
rect 158854 195872 158902 195928
rect 158958 195880 160834 195928
rect 160890 195880 160895 195936
rect 158958 195878 160895 195880
rect 158958 195872 158963 195878
rect 160829 195875 160895 195878
rect 158854 195870 158963 195872
rect 158897 195867 158963 195870
rect 140773 195666 140839 195669
rect 143582 195666 144164 195674
rect 157149 195666 157215 195669
rect 140773 195664 144164 195666
rect 140773 195608 140778 195664
rect 140834 195614 144164 195664
rect 155910 195664 157215 195666
rect 140834 195608 143642 195614
rect 140773 195606 143642 195608
rect 155910 195608 157154 195664
rect 157210 195608 157215 195664
rect 155910 195606 157215 195608
rect 140773 195603 140839 195606
rect 139393 195530 139459 195533
rect 139393 195528 142170 195530
rect 139393 195472 139398 195528
rect 139454 195498 142170 195528
rect 139454 195472 142692 195498
rect 139393 195470 142692 195472
rect 139393 195467 139459 195470
rect 142110 195438 142692 195470
rect 155910 195340 155970 195606
rect 157149 195603 157215 195606
rect 580073 192538 580139 192541
rect 583520 192538 584960 192628
rect 580073 192536 584960 192538
rect 580073 192480 580078 192536
rect 580134 192480 584960 192536
rect 580073 192478 584960 192480
rect 580073 192475 580139 192478
rect 583520 192388 584960 192478
rect 140957 191858 141023 191861
rect 143214 191858 143980 191900
rect 140957 191856 143980 191858
rect 140957 191800 140962 191856
rect 141018 191840 143980 191856
rect 141018 191800 143274 191840
rect 140957 191798 143274 191800
rect 140957 191795 141023 191798
rect 140865 191722 140931 191725
rect 143398 191722 143980 191760
rect 140865 191720 143980 191722
rect 140865 191664 140870 191720
rect 140926 191700 143980 191720
rect 140926 191664 143458 191700
rect 140865 191662 143458 191664
rect 140865 191659 140931 191662
rect 140773 191586 140839 191589
rect 143582 191586 144164 191630
rect 140773 191584 144164 191586
rect 140773 191528 140778 191584
rect 140834 191570 144164 191584
rect 140834 191528 143642 191570
rect 140773 191526 143642 191528
rect 140773 191523 140839 191526
rect 140957 190906 141023 190909
rect 144134 190906 144194 191460
rect 144545 191042 144611 191045
rect 144862 191042 144868 191044
rect 144545 191040 144868 191042
rect 144545 190984 144550 191040
rect 144606 190984 144868 191040
rect 144545 190982 144868 190984
rect 144545 190979 144611 190982
rect 144862 190980 144868 190982
rect 144932 190980 144938 191044
rect 140957 190904 144194 190906
rect 140957 190848 140962 190904
rect 141018 190848 144194 190904
rect 140957 190846 144194 190848
rect 140957 190843 141023 190846
rect 140865 190362 140931 190365
rect 140998 190362 141004 190364
rect 140865 190360 141004 190362
rect 140865 190304 140870 190360
rect 140926 190304 141004 190360
rect 140865 190302 141004 190304
rect 140865 190299 140931 190302
rect 140998 190300 141004 190302
rect 141068 190300 141074 190364
rect 145833 189000 145899 189005
rect -960 188866 480 188956
rect 145833 188944 145838 189000
rect 145894 188944 145899 189000
rect 145833 188939 145899 188944
rect 3325 188866 3391 188869
rect -960 188864 3391 188866
rect -960 188808 3330 188864
rect 3386 188808 3391 188864
rect -960 188806 3391 188808
rect -960 188716 480 188806
rect 3325 188803 3391 188806
rect 145836 188594 145896 188939
rect 146150 188594 146156 188596
rect 145836 188534 146156 188594
rect 146150 188532 146156 188534
rect 146220 188532 146226 188596
rect 140957 184378 141023 184381
rect 141734 184378 141740 184380
rect 140957 184376 141740 184378
rect 140957 184320 140962 184376
rect 141018 184320 141740 184376
rect 140957 184318 141740 184320
rect 140957 184315 141023 184318
rect 141734 184316 141740 184318
rect 141804 184316 141810 184380
rect 140773 184244 140839 184245
rect 140773 184240 140820 184244
rect 140884 184242 140890 184244
rect 140773 184184 140778 184240
rect 140773 184180 140820 184184
rect 140884 184182 140930 184242
rect 140884 184180 140890 184182
rect 140773 184179 140839 184180
rect 140865 184106 140931 184109
rect 142838 184106 142844 184108
rect 140865 184104 142844 184106
rect 140865 184048 140870 184104
rect 140926 184048 142844 184104
rect 140865 184046 142844 184048
rect 140865 184043 140931 184046
rect 142838 184044 142844 184046
rect 142908 184044 142914 184108
rect 144913 182204 144979 182205
rect 144862 182140 144868 182204
rect 144932 182202 144979 182204
rect 144932 182200 145024 182202
rect 144974 182144 145024 182200
rect 144932 182142 145024 182144
rect 144932 182140 144979 182142
rect 144913 182139 144979 182140
rect 144913 181250 144979 181253
rect 145046 181250 145052 181252
rect 144913 181248 145052 181250
rect 144913 181192 144918 181248
rect 144974 181192 145052 181248
rect 144913 181190 145052 181192
rect 144913 181187 144979 181190
rect 145046 181188 145052 181190
rect 145116 181188 145122 181252
rect 145189 181250 145255 181253
rect 152590 181250 152596 181252
rect 145189 181248 152596 181250
rect 145189 181192 145194 181248
rect 145250 181192 152596 181248
rect 145189 181190 152596 181192
rect 145189 181187 145255 181190
rect 152590 181188 152596 181190
rect 152660 181188 152666 181252
rect 142470 180916 142476 180980
rect 142540 180978 142546 180980
rect 144637 180978 144703 180981
rect 142540 180976 144703 180978
rect 142540 180920 144642 180976
rect 144698 180920 144703 180976
rect 142540 180918 144703 180920
rect 142540 180916 142546 180918
rect 144637 180915 144703 180918
rect 580073 179210 580139 179213
rect 583520 179210 584960 179300
rect 580073 179208 584960 179210
rect 580073 179152 580078 179208
rect 580134 179152 584960 179208
rect 580073 179150 584960 179152
rect 580073 179147 580139 179150
rect 583520 179060 584960 179150
rect 142838 178876 142844 178940
rect 142908 178938 142914 178940
rect 144085 178938 144151 178941
rect 142908 178936 144151 178938
rect 142908 178880 144090 178936
rect 144146 178880 144151 178936
rect 142908 178878 144151 178880
rect 142908 178876 142914 178878
rect 144085 178875 144151 178878
rect 140998 178740 141004 178804
rect 141068 178802 141074 178804
rect 141601 178802 141667 178805
rect 141785 178804 141851 178805
rect 141068 178800 141667 178802
rect 141068 178744 141606 178800
rect 141662 178744 141667 178800
rect 141068 178742 141667 178744
rect 141068 178740 141074 178742
rect 141601 178739 141667 178742
rect 141734 178740 141740 178804
rect 141804 178802 141851 178804
rect 141804 178800 141896 178802
rect 141846 178744 141896 178800
rect 141804 178742 141896 178744
rect 141804 178740 141851 178742
rect 141785 178739 141851 178740
rect 140814 178604 140820 178668
rect 140884 178666 140890 178668
rect 142061 178666 142127 178669
rect 140884 178664 142127 178666
rect 140884 178608 142066 178664
rect 142122 178608 142127 178664
rect 140884 178606 142127 178608
rect 140884 178604 140890 178606
rect 142061 178603 142127 178606
rect 145046 177380 145052 177444
rect 145116 177442 145122 177444
rect 145465 177442 145531 177445
rect 145116 177440 145531 177442
rect 145116 177384 145470 177440
rect 145526 177384 145531 177440
rect 145116 177382 145531 177384
rect 145116 177380 145122 177382
rect 145465 177379 145531 177382
rect 158662 176428 158668 176492
rect 158732 176490 158738 176492
rect 158805 176490 158871 176493
rect 158732 176488 158871 176490
rect 158732 176432 158810 176488
rect 158866 176432 158871 176488
rect 158732 176430 158871 176432
rect 158732 176428 158738 176430
rect 158805 176427 158871 176430
rect -960 175796 480 176036
rect 149237 175810 149303 175813
rect 159173 175810 159239 175813
rect 149237 175808 159239 175810
rect 149237 175752 149242 175808
rect 149298 175752 159178 175808
rect 159234 175752 159239 175808
rect 149237 175750 159239 175752
rect 149237 175747 149303 175750
rect 159173 175747 159239 175750
rect 164233 175810 164299 175813
rect 166993 175810 167059 175813
rect 164233 175808 167059 175810
rect 164233 175752 164238 175808
rect 164294 175752 166998 175808
rect 167054 175752 167059 175808
rect 164233 175750 167059 175752
rect 164233 175747 164299 175750
rect 166993 175747 167059 175750
rect 149329 175402 149395 175405
rect 159081 175402 159147 175405
rect 149329 175400 159147 175402
rect 149329 175344 149334 175400
rect 149390 175344 159086 175400
rect 159142 175344 159147 175400
rect 149329 175342 159147 175344
rect 149329 175339 149395 175342
rect 159081 175339 159147 175342
rect 148685 175266 148751 175269
rect 154573 175266 154639 175269
rect 148685 175264 154639 175266
rect 148685 175208 148690 175264
rect 148746 175208 154578 175264
rect 154634 175208 154639 175264
rect 148685 175206 154639 175208
rect 148685 175203 148751 175206
rect 154573 175203 154639 175206
rect 142521 172956 142587 172957
rect 142470 172954 142476 172956
rect 142430 172894 142476 172954
rect 142540 172952 142587 172956
rect 142582 172896 142587 172952
rect 142470 172892 142476 172894
rect 142540 172892 142587 172896
rect 142521 172891 142587 172892
rect 158437 172954 158503 172957
rect 158662 172954 158668 172956
rect 158437 172952 158668 172954
rect 158437 172896 158442 172952
rect 158498 172896 158668 172952
rect 158437 172894 158668 172896
rect 158437 172891 158503 172894
rect 158662 172892 158668 172894
rect 158732 172892 158738 172956
rect 152590 169492 152596 169556
rect 152660 169554 152666 169556
rect 154481 169554 154547 169557
rect 152660 169552 154547 169554
rect 152660 169496 154486 169552
rect 154542 169496 154547 169552
rect 152660 169494 154547 169496
rect 152660 169492 152666 169494
rect 154481 169491 154547 169494
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 146150 157932 146156 157996
rect 146220 157994 146226 157996
rect 171133 157994 171199 157997
rect 146220 157992 171199 157994
rect 146220 157936 171138 157992
rect 171194 157936 171199 157992
rect 146220 157934 171199 157936
rect 146220 157932 146226 157934
rect 171133 157931 171199 157934
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 117313 137186 117379 137189
rect 118141 137186 118207 137189
rect 117313 137184 120090 137186
rect 117313 137128 117318 137184
rect 117374 137128 118146 137184
rect 118202 137128 120090 137184
rect 117313 137126 120090 137128
rect 117313 137123 117379 137126
rect 118141 137123 118207 137126
rect 120030 137088 120090 137126
rect -960 136778 480 136868
rect 3417 136778 3483 136781
rect -960 136776 3483 136778
rect -960 136720 3422 136776
rect 3478 136720 3483 136776
rect -960 136718 3483 136720
rect -960 136628 480 136718
rect 3417 136715 3483 136718
rect 120625 136234 120691 136237
rect 120582 136232 120691 136234
rect 120582 136176 120630 136232
rect 120686 136176 120691 136232
rect 120582 136171 120691 136176
rect 118233 135554 118299 135557
rect 120582 135554 120642 136171
rect 118233 135552 120642 135554
rect 118233 135496 118238 135552
rect 118294 135496 120642 135552
rect 118233 135494 120642 135496
rect 118233 135491 118299 135494
rect 179830 135418 179890 135592
rect 180885 135418 180951 135421
rect 179830 135416 180951 135418
rect 179830 135360 180890 135416
rect 180946 135360 180951 135416
rect 179830 135358 180951 135360
rect 180885 135355 180951 135358
rect 117313 134058 117379 134061
rect 120030 134058 120090 134096
rect 117313 134056 120090 134058
rect 117313 134000 117318 134056
rect 117374 134000 120090 134056
rect 117313 133998 120090 134000
rect 117313 133995 117379 133998
rect 179830 133922 179890 134096
rect 183001 133922 183067 133925
rect 179830 133920 183067 133922
rect 179830 133864 183006 133920
rect 183062 133864 183067 133920
rect 179830 133862 183067 133864
rect 183001 133859 183067 133862
rect 182173 133242 182239 133245
rect 179830 133240 182239 133242
rect 179830 133184 182178 133240
rect 182234 133184 182239 133240
rect 179830 133182 182239 133184
rect 179830 132600 179890 133182
rect 182173 133179 182239 133182
rect 117313 132562 117379 132565
rect 120030 132562 120090 132600
rect 117313 132560 120090 132562
rect 117313 132504 117318 132560
rect 117374 132504 120090 132560
rect 117313 132502 120090 132504
rect 117313 132499 117379 132502
rect 179505 131746 179571 131749
rect 179462 131744 179571 131746
rect 179462 131688 179510 131744
rect 179566 131688 179571 131744
rect 179462 131683 179571 131688
rect 117313 131202 117379 131205
rect 117313 131200 120090 131202
rect 117313 131144 117318 131200
rect 117374 131144 120090 131200
rect 117313 131142 120090 131144
rect 117313 131139 117379 131142
rect 120030 131104 120090 131142
rect 179462 131104 179522 131683
rect 117313 129706 117379 129709
rect 180977 129706 181043 129709
rect 117313 129704 120090 129706
rect 117313 129648 117318 129704
rect 117374 129648 120090 129704
rect 117313 129646 120090 129648
rect 117313 129643 117379 129646
rect 120030 129608 120090 129646
rect 179830 129704 181043 129706
rect 179830 129648 180982 129704
rect 181038 129648 181043 129704
rect 179830 129646 181043 129648
rect 179830 129608 179890 129646
rect 180977 129643 181043 129646
rect 182357 128346 182423 128349
rect 179830 128344 182423 128346
rect 179830 128288 182362 128344
rect 182418 128288 182423 128344
rect 179830 128286 182423 128288
rect 117313 128210 117379 128213
rect 117313 128208 120090 128210
rect 117313 128152 117318 128208
rect 117374 128152 120090 128208
rect 117313 128150 120090 128152
rect 117313 128147 117379 128150
rect 120030 128112 120090 128150
rect 179830 128112 179890 128286
rect 182357 128283 182423 128286
rect 182909 126986 182975 126989
rect 179830 126984 182975 126986
rect 179830 126928 182914 126984
rect 182970 126928 182975 126984
rect 179830 126926 182975 126928
rect 117313 126850 117379 126853
rect 117313 126848 120090 126850
rect 117313 126792 117318 126848
rect 117374 126792 120090 126848
rect 117313 126790 120090 126792
rect 117313 126787 117379 126790
rect 120030 126616 120090 126790
rect 179830 126616 179890 126926
rect 182909 126923 182975 126926
rect 580073 126034 580139 126037
rect 583520 126034 584960 126124
rect 580073 126032 584960 126034
rect 580073 125976 580078 126032
rect 580134 125976 584960 126032
rect 580073 125974 584960 125976
rect 580073 125971 580139 125974
rect 583520 125884 584960 125974
rect 118141 125490 118207 125493
rect 118141 125488 120090 125490
rect 118141 125432 118146 125488
rect 118202 125432 120090 125488
rect 118141 125430 120090 125432
rect 118141 125427 118207 125430
rect 120030 125120 120090 125430
rect 182725 125354 182791 125357
rect 179830 125352 182791 125354
rect 179830 125296 182730 125352
rect 182786 125296 182791 125352
rect 179830 125294 182791 125296
rect 179830 125120 179890 125294
rect 182725 125291 182791 125294
rect 182265 124130 182331 124133
rect 179830 124128 182331 124130
rect 179830 124072 182270 124128
rect 182326 124072 182331 124128
rect 179830 124070 182331 124072
rect 117313 123858 117379 123861
rect 117313 123856 120090 123858
rect -960 123572 480 123812
rect 117313 123800 117318 123856
rect 117374 123800 120090 123856
rect 117313 123798 120090 123800
rect 117313 123795 117379 123798
rect 120030 123624 120090 123798
rect 179830 123624 179890 124070
rect 182265 124067 182331 124070
rect 117313 122770 117379 122773
rect 180793 122770 180859 122773
rect 117313 122768 120090 122770
rect 117313 122712 117318 122768
rect 117374 122712 120090 122768
rect 117313 122710 120090 122712
rect 117313 122707 117379 122710
rect 120030 122128 120090 122710
rect 179830 122768 180859 122770
rect 179830 122712 180798 122768
rect 180854 122712 180859 122768
rect 179830 122710 180859 122712
rect 179830 122128 179890 122710
rect 180793 122707 180859 122710
rect 117313 121274 117379 121277
rect 182817 121274 182883 121277
rect 117313 121272 120090 121274
rect 117313 121216 117318 121272
rect 117374 121216 120090 121272
rect 117313 121214 120090 121216
rect 117313 121211 117379 121214
rect 120030 120632 120090 121214
rect 179830 121272 182883 121274
rect 179830 121216 182822 121272
rect 182878 121216 182883 121272
rect 179830 121214 182883 121216
rect 179830 120632 179890 121214
rect 182817 121211 182883 121214
rect 117313 119778 117379 119781
rect 182633 119778 182699 119781
rect 117313 119776 120090 119778
rect 117313 119720 117318 119776
rect 117374 119720 120090 119776
rect 117313 119718 120090 119720
rect 117313 119715 117379 119718
rect 120030 119136 120090 119718
rect 179830 119776 182699 119778
rect 179830 119720 182638 119776
rect 182694 119720 182699 119776
rect 179830 119718 182699 119720
rect 179830 119136 179890 119718
rect 182633 119715 182699 119718
rect 117313 118282 117379 118285
rect 179597 118282 179663 118285
rect 117313 118280 120090 118282
rect 117313 118224 117318 118280
rect 117374 118224 120090 118280
rect 117313 118222 120090 118224
rect 117313 118219 117379 118222
rect 120030 117640 120090 118222
rect 179597 118280 179706 118282
rect 179597 118224 179602 118280
rect 179658 118224 179706 118280
rect 179597 118219 179706 118224
rect 179646 117640 179706 118219
rect 117313 116786 117379 116789
rect 182541 116786 182607 116789
rect 117313 116784 120090 116786
rect 117313 116728 117318 116784
rect 117374 116728 120090 116784
rect 117313 116726 120090 116728
rect 117313 116723 117379 116726
rect 120030 116144 120090 116726
rect 179830 116784 182607 116786
rect 179830 116728 182546 116784
rect 182602 116728 182607 116784
rect 179830 116726 182607 116728
rect 179830 116144 179890 116726
rect 182541 116723 182607 116726
rect 117313 115290 117379 115293
rect 181069 115290 181135 115293
rect 117313 115288 120090 115290
rect 117313 115232 117318 115288
rect 117374 115232 120090 115288
rect 117313 115230 120090 115232
rect 117313 115227 117379 115230
rect 120030 114648 120090 115230
rect 179830 115288 181135 115290
rect 179830 115232 181074 115288
rect 181130 115232 181135 115288
rect 179830 115230 181135 115232
rect 179830 114648 179890 115230
rect 181069 115227 181135 115230
rect 117313 113114 117379 113117
rect 120030 113114 120090 113152
rect 117313 113112 120090 113114
rect 117313 113056 117318 113112
rect 117374 113056 120090 113112
rect 117313 113054 120090 113056
rect 179830 113114 179890 113152
rect 181161 113114 181227 113117
rect 179830 113112 181227 113114
rect 179830 113056 181166 113112
rect 181222 113056 181227 113112
rect 179830 113054 181227 113056
rect 117313 113051 117379 113054
rect 181161 113051 181227 113054
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect 179413 111890 179479 111893
rect 179413 111888 179522 111890
rect 179413 111832 179418 111888
rect 179474 111832 179522 111888
rect 179413 111827 179522 111832
rect 117313 111754 117379 111757
rect 117313 111752 120090 111754
rect 117313 111696 117318 111752
rect 117374 111696 120090 111752
rect 117313 111694 120090 111696
rect 117313 111691 117379 111694
rect 120030 111656 120090 111694
rect 179462 111656 179522 111827
rect -960 110666 480 110756
rect 3233 110666 3299 110669
rect -960 110664 3299 110666
rect -960 110608 3238 110664
rect 3294 110608 3299 110664
rect -960 110606 3299 110608
rect -960 110516 480 110606
rect 3233 110603 3299 110606
rect 182449 110394 182515 110397
rect 179830 110392 182515 110394
rect 179830 110336 182454 110392
rect 182510 110336 182515 110392
rect 179830 110334 182515 110336
rect 117313 110258 117379 110261
rect 117313 110256 120090 110258
rect 117313 110200 117318 110256
rect 117374 110200 120090 110256
rect 117313 110198 120090 110200
rect 117313 110195 117379 110198
rect 120030 110160 120090 110198
rect 179830 110160 179890 110334
rect 182449 110331 182515 110334
rect 117313 108898 117379 108901
rect 183461 108898 183527 108901
rect 117313 108896 120090 108898
rect 117313 108840 117318 108896
rect 117374 108840 120090 108896
rect 117313 108838 120090 108840
rect 117313 108835 117379 108838
rect 120030 108664 120090 108838
rect 179830 108896 183527 108898
rect 179830 108840 183466 108896
rect 183522 108840 183527 108896
rect 179830 108838 183527 108840
rect 179830 108664 179890 108838
rect 183461 108835 183527 108838
rect 117313 107538 117379 107541
rect 117313 107536 120090 107538
rect 117313 107480 117318 107536
rect 117374 107480 120090 107536
rect 117313 107478 120090 107480
rect 117313 107475 117379 107478
rect 120030 107168 120090 107478
rect 183461 107402 183527 107405
rect 179830 107400 183527 107402
rect 179830 107344 183466 107400
rect 183522 107344 183527 107400
rect 179830 107342 183527 107344
rect 179830 107168 179890 107342
rect 183461 107339 183527 107342
rect 118601 106178 118667 106181
rect 118601 106176 120090 106178
rect 118601 106120 118606 106176
rect 118662 106120 120090 106176
rect 118601 106118 120090 106120
rect 118601 106115 118667 106118
rect 120030 105672 120090 106118
rect 183461 106042 183527 106045
rect 179830 106040 183527 106042
rect 179830 105984 183466 106040
rect 183522 105984 183527 106040
rect 179830 105982 183527 105984
rect 179830 105672 179890 105982
rect 183461 105979 183527 105982
rect 119337 104818 119403 104821
rect 119337 104816 120090 104818
rect 119337 104760 119342 104816
rect 119398 104760 120090 104816
rect 119337 104758 120090 104760
rect 119337 104755 119403 104758
rect 120030 104176 120090 104758
rect 183461 104546 183527 104549
rect 179830 104544 183527 104546
rect 179830 104488 183466 104544
rect 183522 104488 183527 104544
rect 179830 104486 183527 104488
rect 179830 104176 179890 104486
rect 183461 104483 183527 104486
rect 119061 103186 119127 103189
rect 119061 103184 120090 103186
rect 119061 103128 119066 103184
rect 119122 103128 120090 103184
rect 119061 103126 120090 103128
rect 119061 103123 119127 103126
rect 120030 102680 120090 103126
rect 183461 103050 183527 103053
rect 179830 103048 183527 103050
rect 179830 102992 183466 103048
rect 183522 102992 183527 103048
rect 179830 102990 183527 102992
rect 179830 102680 179890 102990
rect 183461 102987 183527 102990
rect 120625 101826 120691 101829
rect 120582 101824 120691 101826
rect 120582 101768 120630 101824
rect 120686 101768 120691 101824
rect 120582 101763 120691 101768
rect 120582 101184 120642 101763
rect 183461 101690 183527 101693
rect 179830 101688 183527 101690
rect 179830 101632 183466 101688
rect 183522 101632 183527 101688
rect 179830 101630 183527 101632
rect 179830 101184 179890 101630
rect 183461 101627 183527 101630
rect 118969 100330 119035 100333
rect 118969 100328 120090 100330
rect 118969 100272 118974 100328
rect 119030 100272 120090 100328
rect 118969 100270 120090 100272
rect 118969 100267 119035 100270
rect 120030 99688 120090 100270
rect 182817 100194 182883 100197
rect 179830 100192 182883 100194
rect 179830 100136 182822 100192
rect 182878 100136 182883 100192
rect 179830 100134 182883 100136
rect 179830 99688 179890 100134
rect 182817 100131 182883 100134
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 119153 98834 119219 98837
rect 182817 98834 182883 98837
rect 119153 98832 120090 98834
rect 119153 98776 119158 98832
rect 119214 98776 120090 98832
rect 119153 98774 120090 98776
rect 119153 98771 119219 98774
rect 120030 98192 120090 98774
rect 179830 98832 182883 98834
rect 179830 98776 182822 98832
rect 182878 98776 182883 98832
rect 179830 98774 182883 98776
rect 179830 98192 179890 98774
rect 182817 98771 182883 98774
rect -960 97610 480 97700
rect 3325 97610 3391 97613
rect -960 97608 3391 97610
rect -960 97552 3330 97608
rect 3386 97552 3391 97608
rect -960 97550 3391 97552
rect -960 97460 480 97550
rect 3325 97547 3391 97550
rect 119245 97338 119311 97341
rect 183461 97338 183527 97341
rect 119245 97336 120090 97338
rect 119245 97280 119250 97336
rect 119306 97280 120090 97336
rect 119245 97278 120090 97280
rect 119245 97275 119311 97278
rect 120030 96696 120090 97278
rect 179830 97336 183527 97338
rect 179830 97280 183466 97336
rect 183522 97280 183527 97336
rect 179830 97278 183527 97280
rect 179830 96696 179890 97278
rect 183461 97275 183527 97278
rect 118233 95162 118299 95165
rect 120030 95162 120090 95200
rect 118233 95160 120090 95162
rect 118233 95104 118238 95160
rect 118294 95104 120090 95160
rect 118233 95102 120090 95104
rect 179830 95162 179890 95200
rect 183461 95162 183527 95165
rect 179830 95160 183527 95162
rect 179830 95104 183466 95160
rect 183522 95104 183527 95160
rect 179830 95102 183527 95104
rect 118233 95099 118299 95102
rect 183461 95099 183527 95102
rect 118877 93802 118943 93805
rect 183461 93802 183527 93805
rect 118877 93800 120090 93802
rect 118877 93744 118882 93800
rect 118938 93744 120090 93800
rect 118877 93742 120090 93744
rect 118877 93739 118943 93742
rect 120030 93704 120090 93742
rect 179830 93800 183527 93802
rect 179830 93744 183466 93800
rect 183522 93744 183527 93800
rect 179830 93742 183527 93744
rect 179830 93704 179890 93742
rect 183461 93739 183527 93742
rect 118693 92442 118759 92445
rect 118693 92440 120090 92442
rect 118693 92384 118698 92440
rect 118754 92384 120090 92440
rect 118693 92382 120090 92384
rect 118693 92379 118759 92382
rect 120030 92208 120090 92382
rect 183461 92306 183527 92309
rect 179830 92304 183527 92306
rect 179830 92248 183466 92304
rect 183522 92248 183527 92304
rect 179830 92246 183527 92248
rect 179830 92208 179890 92246
rect 183461 92243 183527 92246
rect 118325 91082 118391 91085
rect 118325 91080 120090 91082
rect 118325 91024 118330 91080
rect 118386 91024 120090 91080
rect 118325 91022 120090 91024
rect 118325 91019 118391 91022
rect 120030 90712 120090 91022
rect 183461 90946 183527 90949
rect 179830 90944 183527 90946
rect 179830 90888 183466 90944
rect 183522 90888 183527 90944
rect 179830 90886 183527 90888
rect 179830 90712 179890 90886
rect 183461 90883 183527 90886
rect 118417 89722 118483 89725
rect 118417 89720 120090 89722
rect 118417 89664 118422 89720
rect 118478 89664 120090 89720
rect 118417 89662 120090 89664
rect 118417 89659 118483 89662
rect 120030 89216 120090 89662
rect 182265 89450 182331 89453
rect 179830 89448 182331 89450
rect 179830 89392 182270 89448
rect 182326 89392 182331 89448
rect 179830 89390 182331 89392
rect 179830 89216 179890 89390
rect 182265 89387 182331 89390
rect 118509 88226 118575 88229
rect 118509 88224 120090 88226
rect 118509 88168 118514 88224
rect 118570 88168 120090 88224
rect 118509 88166 120090 88168
rect 118509 88163 118575 88166
rect 120030 87720 120090 88166
rect 183461 88090 183527 88093
rect 179830 88088 183527 88090
rect 179830 88032 183466 88088
rect 183522 88032 183527 88088
rect 179830 88030 183527 88032
rect 179830 87720 179890 88030
rect 183461 88027 183527 88030
rect 118141 86866 118207 86869
rect 118141 86864 120090 86866
rect 118141 86808 118146 86864
rect 118202 86808 120090 86864
rect 118141 86806 120090 86808
rect 118141 86803 118207 86806
rect 120030 86224 120090 86806
rect 183461 86594 183527 86597
rect 179830 86592 183527 86594
rect 179830 86536 183466 86592
rect 183522 86536 183527 86592
rect 179830 86534 183527 86536
rect 179830 86224 179890 86534
rect 183461 86531 183527 86534
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 118785 85370 118851 85373
rect 118785 85368 120090 85370
rect 118785 85312 118790 85368
rect 118846 85312 120090 85368
rect 118785 85310 120090 85312
rect 118785 85307 118851 85310
rect -960 84690 480 84780
rect 120030 84728 120090 85310
rect 182173 85098 182239 85101
rect 179830 85096 182239 85098
rect 179830 85040 182178 85096
rect 182234 85040 182239 85096
rect 179830 85038 182239 85040
rect 179830 84728 179890 85038
rect 182173 85035 182239 85038
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 182265 83874 182331 83877
rect 179830 83872 182331 83874
rect 179830 83816 182270 83872
rect 182326 83816 182331 83872
rect 179830 83814 182331 83816
rect 117865 83738 117931 83741
rect 117865 83736 120090 83738
rect 117865 83680 117870 83736
rect 117926 83680 120090 83736
rect 117865 83678 120090 83680
rect 117865 83675 117931 83678
rect 120030 83232 120090 83678
rect 179830 83232 179890 83814
rect 182265 83811 182331 83814
rect 120582 81565 120642 81736
rect 120582 81560 120691 81565
rect 120582 81504 120630 81560
rect 120686 81504 120691 81560
rect 120582 81502 120691 81504
rect 179830 81562 179890 81736
rect 182817 81562 182883 81565
rect 179830 81560 182883 81562
rect 179830 81504 182822 81560
rect 182878 81504 182883 81560
rect 179830 81502 182883 81504
rect 120625 81499 120691 81502
rect 182817 81499 182883 81502
rect 118509 80202 118575 80205
rect 120030 80202 120090 80240
rect 118509 80200 120090 80202
rect 118509 80144 118514 80200
rect 118570 80144 120090 80200
rect 118509 80142 120090 80144
rect 179830 80202 179890 80240
rect 183461 80202 183527 80205
rect 179830 80200 183527 80202
rect 179830 80144 183466 80200
rect 183522 80144 183527 80200
rect 179830 80142 183527 80144
rect 118509 80139 118575 80142
rect 183461 80139 183527 80142
rect 118417 78706 118483 78709
rect 120030 78706 120090 78744
rect 118417 78704 120090 78706
rect 118417 78648 118422 78704
rect 118478 78648 120090 78704
rect 118417 78646 120090 78648
rect 118417 78643 118483 78646
rect 153510 78508 153516 78572
rect 153580 78570 153586 78572
rect 163998 78570 164004 78572
rect 153580 78510 164004 78570
rect 153580 78508 153586 78510
rect 163998 78508 164004 78510
rect 164068 78508 164074 78572
rect 165286 78508 165292 78572
rect 165356 78570 165362 78572
rect 173566 78570 173572 78572
rect 165356 78510 173572 78570
rect 165356 78508 165362 78510
rect 173566 78508 173572 78510
rect 173636 78508 173642 78572
rect 178953 78570 179019 78573
rect 174678 78568 179019 78570
rect 174678 78512 178958 78568
rect 179014 78512 179019 78568
rect 174678 78510 179019 78512
rect 162158 78372 162164 78436
rect 162228 78434 162234 78436
rect 171358 78434 171364 78436
rect 162228 78374 171364 78434
rect 162228 78372 162234 78374
rect 171358 78372 171364 78374
rect 171428 78372 171434 78436
rect 171542 78372 171548 78436
rect 171612 78434 171618 78436
rect 174678 78434 174738 78510
rect 178953 78507 179019 78510
rect 171612 78374 174738 78434
rect 174813 78434 174879 78437
rect 180149 78434 180215 78437
rect 174813 78432 180215 78434
rect 174813 78376 174818 78432
rect 174874 78376 180154 78432
rect 180210 78376 180215 78432
rect 174813 78374 180215 78376
rect 171612 78372 171618 78374
rect 174813 78371 174879 78374
rect 180149 78371 180215 78374
rect 144870 78238 154590 78298
rect 6913 78162 6979 78165
rect 144870 78162 144930 78238
rect 145414 78162 145420 78164
rect 6913 78160 144930 78162
rect 6913 78104 6918 78160
rect 6974 78104 144930 78160
rect 6913 78102 144930 78104
rect 145054 78102 145420 78162
rect 6913 78099 6979 78102
rect 3693 78026 3759 78029
rect 130694 78026 130700 78028
rect 3693 78024 130700 78026
rect 3693 77968 3698 78024
rect 3754 77968 130700 78024
rect 3693 77966 130700 77968
rect 3693 77963 3759 77966
rect 130694 77964 130700 77966
rect 130764 77964 130770 78028
rect 131062 77964 131068 78028
rect 131132 78026 131138 78028
rect 144862 78026 144868 78028
rect 131132 77966 144868 78026
rect 131132 77964 131138 77966
rect 144862 77964 144868 77966
rect 144932 77964 144938 78028
rect 3366 77828 3372 77892
rect 3436 77890 3442 77892
rect 123753 77890 123819 77893
rect 126007 77890 126073 77893
rect 3436 77830 118710 77890
rect 3436 77828 3442 77830
rect 118650 77618 118710 77830
rect 123753 77888 126073 77890
rect 123753 77832 123758 77888
rect 123814 77832 126012 77888
rect 126068 77832 126073 77888
rect 123753 77830 126073 77832
rect 123753 77827 123819 77830
rect 126007 77827 126073 77830
rect 126283 77888 126349 77893
rect 126283 77832 126288 77888
rect 126344 77832 126349 77888
rect 126283 77827 126349 77832
rect 126646 77828 126652 77892
rect 126716 77890 126722 77892
rect 127571 77890 127637 77893
rect 128031 77890 128097 77893
rect 126716 77888 127637 77890
rect 126716 77832 127576 77888
rect 127632 77832 127637 77888
rect 126716 77830 127637 77832
rect 126716 77828 126722 77830
rect 127571 77827 127637 77830
rect 127758 77888 128097 77890
rect 127758 77832 128036 77888
rect 128092 77832 128097 77888
rect 127758 77830 128097 77832
rect 126286 77757 126346 77827
rect 126237 77752 126346 77757
rect 126237 77696 126242 77752
rect 126298 77696 126346 77752
rect 126237 77694 126346 77696
rect 127525 77754 127591 77757
rect 127758 77754 127818 77830
rect 128031 77827 128097 77830
rect 128670 77828 128676 77892
rect 128740 77890 128746 77892
rect 129043 77890 129109 77893
rect 128740 77888 129109 77890
rect 128740 77832 129048 77888
rect 129104 77832 129109 77888
rect 128740 77830 129109 77832
rect 128740 77828 128746 77830
rect 129043 77827 129109 77830
rect 129590 77828 129596 77892
rect 129660 77890 129666 77892
rect 129871 77890 129937 77893
rect 130515 77892 130581 77893
rect 130510 77890 130516 77892
rect 129660 77888 129937 77890
rect 129660 77832 129876 77888
rect 129932 77832 129937 77888
rect 129660 77830 129937 77832
rect 130424 77830 130516 77890
rect 129660 77828 129666 77830
rect 129871 77827 129937 77830
rect 130510 77828 130516 77830
rect 130580 77828 130586 77892
rect 131430 77828 131436 77892
rect 131500 77890 131506 77892
rect 131711 77890 131777 77893
rect 131987 77892 132053 77893
rect 131982 77890 131988 77892
rect 131500 77888 131777 77890
rect 131500 77832 131716 77888
rect 131772 77832 131777 77888
rect 131500 77830 131777 77832
rect 131896 77830 131988 77890
rect 131500 77828 131506 77830
rect 130515 77827 130581 77828
rect 131711 77827 131777 77830
rect 131982 77828 131988 77830
rect 132052 77828 132058 77892
rect 132355 77888 132421 77893
rect 132539 77892 132605 77893
rect 132907 77892 132973 77893
rect 132355 77832 132360 77888
rect 132416 77832 132421 77888
rect 131987 77827 132053 77828
rect 132355 77827 132421 77832
rect 132534 77828 132540 77892
rect 132604 77890 132610 77892
rect 132902 77890 132908 77892
rect 132604 77830 132696 77890
rect 132816 77830 132908 77890
rect 132604 77828 132610 77830
rect 132902 77828 132908 77830
rect 132972 77828 132978 77892
rect 133183 77890 133249 77893
rect 133140 77888 133249 77890
rect 133140 77832 133188 77888
rect 133244 77832 133249 77888
rect 132539 77827 132605 77828
rect 132907 77827 132973 77828
rect 133140 77827 133249 77832
rect 133643 77888 133709 77893
rect 133827 77890 133893 77893
rect 133643 77832 133648 77888
rect 133704 77832 133709 77888
rect 133643 77827 133709 77832
rect 133784 77888 133893 77890
rect 133784 77832 133832 77888
rect 133888 77832 133893 77888
rect 133784 77827 133893 77832
rect 134190 77828 134196 77892
rect 134260 77890 134266 77892
rect 134379 77890 134445 77893
rect 134260 77888 134445 77890
rect 134260 77832 134384 77888
rect 134440 77832 134445 77888
rect 134260 77830 134445 77832
rect 134260 77828 134266 77830
rect 134379 77827 134445 77830
rect 134747 77888 134813 77893
rect 136035 77892 136101 77893
rect 136030 77890 136036 77892
rect 134747 77832 134752 77888
rect 134808 77832 134813 77888
rect 134747 77827 134813 77832
rect 135944 77830 136036 77890
rect 136030 77828 136036 77830
rect 136100 77828 136106 77892
rect 136219 77888 136285 77893
rect 136403 77892 136469 77893
rect 136219 77832 136224 77888
rect 136280 77832 136285 77888
rect 136035 77827 136101 77828
rect 136219 77827 136285 77832
rect 136398 77828 136404 77892
rect 136468 77890 136474 77892
rect 136679 77890 136745 77893
rect 136468 77830 136560 77890
rect 136636 77888 136745 77890
rect 136636 77832 136684 77888
rect 136740 77832 136745 77888
rect 136468 77828 136474 77830
rect 136403 77827 136469 77828
rect 136636 77827 136745 77832
rect 136863 77890 136929 77893
rect 137415 77890 137481 77893
rect 144678 77890 144684 77892
rect 136863 77888 137202 77890
rect 136863 77832 136868 77888
rect 136924 77832 137202 77888
rect 136863 77830 137202 77832
rect 136863 77827 136929 77830
rect 127525 77752 127818 77754
rect 127525 77696 127530 77752
rect 127586 77696 127818 77752
rect 127525 77694 127818 77696
rect 126237 77691 126303 77694
rect 127525 77691 127591 77694
rect 130694 77692 130700 77756
rect 130764 77754 130770 77756
rect 130837 77754 130903 77757
rect 130764 77752 130903 77754
rect 130764 77696 130842 77752
rect 130898 77696 130903 77752
rect 130764 77694 130903 77696
rect 130764 77692 130770 77694
rect 130837 77691 130903 77694
rect 131941 77754 132007 77757
rect 132358 77754 132418 77827
rect 133140 77756 133200 77827
rect 131941 77752 132418 77754
rect 131941 77696 131946 77752
rect 132002 77696 132418 77752
rect 131941 77694 132418 77696
rect 131941 77691 132007 77694
rect 133086 77692 133092 77756
rect 133156 77694 133200 77756
rect 133505 77754 133571 77757
rect 133646 77754 133706 77827
rect 133784 77757 133844 77827
rect 133505 77752 133706 77754
rect 133505 77696 133510 77752
rect 133566 77696 133706 77752
rect 133505 77694 133706 77696
rect 133781 77752 133847 77757
rect 133781 77696 133786 77752
rect 133842 77696 133847 77752
rect 133156 77692 133162 77694
rect 133505 77691 133571 77694
rect 133781 77691 133847 77696
rect 134517 77754 134583 77757
rect 134750 77754 134810 77827
rect 135391 77788 135457 77791
rect 135348 77786 135457 77788
rect 135348 77756 135396 77786
rect 134517 77752 134810 77754
rect 134517 77696 134522 77752
rect 134578 77696 134810 77752
rect 134517 77694 134810 77696
rect 134517 77691 134583 77694
rect 135294 77692 135300 77756
rect 135364 77730 135396 77756
rect 135452 77730 135457 77786
rect 136222 77757 136282 77827
rect 135364 77725 135457 77730
rect 136173 77752 136282 77757
rect 135364 77694 135408 77725
rect 136173 77696 136178 77752
rect 136234 77696 136282 77752
rect 136173 77694 136282 77696
rect 136636 77754 136696 77827
rect 136817 77754 136883 77757
rect 136636 77752 136883 77754
rect 136636 77696 136822 77752
rect 136878 77696 136883 77752
rect 136636 77694 136883 77696
rect 135364 77692 135370 77694
rect 136173 77691 136239 77694
rect 136817 77691 136883 77694
rect 136950 77692 136956 77756
rect 137020 77754 137026 77756
rect 137142 77754 137202 77830
rect 137415 77888 137754 77890
rect 137415 77832 137420 77888
rect 137476 77832 137754 77888
rect 137415 77830 137754 77832
rect 137415 77827 137481 77830
rect 137020 77694 137202 77754
rect 137369 77754 137435 77757
rect 137694 77754 137754 77830
rect 137369 77752 137754 77754
rect 137369 77696 137374 77752
rect 137430 77696 137754 77752
rect 137369 77694 137754 77696
rect 137970 77830 144684 77890
rect 137020 77692 137026 77694
rect 137369 77691 137435 77694
rect 137970 77618 138030 77830
rect 144678 77828 144684 77830
rect 144748 77828 144754 77892
rect 144867 77890 144933 77893
rect 145054 77890 145114 78102
rect 145414 78100 145420 78102
rect 145484 78100 145490 78164
rect 154530 78162 154590 78238
rect 155166 78236 155172 78300
rect 155236 78298 155242 78300
rect 163814 78298 163820 78300
rect 155236 78238 163820 78298
rect 155236 78236 155242 78238
rect 163814 78236 163820 78238
rect 163884 78236 163890 78300
rect 163998 78236 164004 78300
rect 164068 78298 164074 78300
rect 164068 78238 173266 78298
rect 164068 78236 164074 78238
rect 169334 78162 169340 78164
rect 154530 78102 169340 78162
rect 169334 78100 169340 78102
rect 169404 78100 169410 78164
rect 145230 77964 145236 78028
rect 145300 78026 145306 78028
rect 155166 78026 155172 78028
rect 145300 77966 155172 78026
rect 145300 77964 145306 77966
rect 155166 77964 155172 77966
rect 155236 77964 155242 78028
rect 167310 78026 167316 78028
rect 167088 77966 167316 78026
rect 155907 77922 155973 77927
rect 144867 77888 145114 77890
rect 144867 77832 144872 77888
rect 144928 77832 145114 77888
rect 144867 77830 145114 77832
rect 144867 77827 144933 77830
rect 145230 77828 145236 77892
rect 145300 77890 145306 77892
rect 145300 77830 149714 77890
rect 145300 77828 145306 77830
rect 138606 77692 138612 77756
rect 138676 77754 138682 77756
rect 138841 77754 138907 77757
rect 138676 77752 138907 77754
rect 138676 77696 138846 77752
rect 138902 77696 138907 77752
rect 138676 77694 138907 77696
rect 138676 77692 138682 77694
rect 138841 77691 138907 77694
rect 139899 77752 139965 77757
rect 143119 77754 143185 77757
rect 139899 77696 139904 77752
rect 139960 77696 139965 77752
rect 139899 77691 139965 77696
rect 142846 77752 143185 77754
rect 142846 77696 143124 77752
rect 143180 77696 143185 77752
rect 142846 77694 143185 77696
rect 118650 77558 138030 77618
rect 131389 77484 131455 77485
rect 132033 77484 132099 77485
rect 131389 77482 131436 77484
rect 131344 77480 131436 77482
rect 131344 77424 131394 77480
rect 131344 77422 131436 77424
rect 131389 77420 131436 77422
rect 131500 77420 131506 77484
rect 131982 77420 131988 77484
rect 132052 77482 132099 77484
rect 132052 77480 132144 77482
rect 132094 77424 132144 77480
rect 132052 77422 132144 77424
rect 132052 77420 132099 77422
rect 136398 77420 136404 77484
rect 136468 77482 136474 77484
rect 136541 77482 136607 77485
rect 136468 77480 136607 77482
rect 136468 77424 136546 77480
rect 136602 77424 136607 77480
rect 136468 77422 136607 77424
rect 136468 77420 136474 77422
rect 131389 77419 131455 77420
rect 132033 77419 132099 77420
rect 136541 77419 136607 77422
rect 137686 77420 137692 77484
rect 137756 77482 137762 77484
rect 138105 77482 138171 77485
rect 137756 77480 138171 77482
rect 137756 77424 138110 77480
rect 138166 77424 138171 77480
rect 137756 77422 138171 77424
rect 137756 77420 137762 77422
rect 138105 77419 138171 77422
rect 138381 77482 138447 77485
rect 138565 77482 138631 77485
rect 138381 77480 138631 77482
rect 138381 77424 138386 77480
rect 138442 77424 138570 77480
rect 138626 77424 138631 77480
rect 138381 77422 138631 77424
rect 139902 77482 139962 77691
rect 140497 77618 140563 77621
rect 140630 77618 140636 77620
rect 140497 77616 140636 77618
rect 140497 77560 140502 77616
rect 140558 77560 140636 77616
rect 140497 77558 140636 77560
rect 140497 77555 140563 77558
rect 140630 77556 140636 77558
rect 140700 77556 140706 77620
rect 142846 77618 142906 77694
rect 143119 77691 143185 77694
rect 143579 77754 143645 77757
rect 144545 77754 144611 77757
rect 145046 77754 145052 77756
rect 143579 77752 143688 77754
rect 143579 77696 143584 77752
rect 143640 77696 143688 77752
rect 143579 77691 143688 77696
rect 144545 77752 145052 77754
rect 144545 77696 144550 77752
rect 144606 77696 145052 77752
rect 144545 77694 145052 77696
rect 144545 77691 144611 77694
rect 145046 77692 145052 77694
rect 145116 77692 145122 77756
rect 145230 77692 145236 77756
rect 145300 77754 145306 77756
rect 145603 77754 145669 77757
rect 145300 77752 145669 77754
rect 145300 77696 145608 77752
rect 145664 77696 145669 77752
rect 145300 77694 145669 77696
rect 145300 77692 145306 77694
rect 145603 77691 145669 77694
rect 145833 77754 145899 77757
rect 146247 77754 146313 77757
rect 145833 77752 146034 77754
rect 145833 77696 145838 77752
rect 145894 77696 146034 77752
rect 145833 77694 146034 77696
rect 145833 77691 145899 77694
rect 143073 77618 143139 77621
rect 142846 77616 143139 77618
rect 142846 77560 143078 77616
rect 143134 77560 143139 77616
rect 142846 77558 143139 77560
rect 143628 77618 143688 77691
rect 144862 77618 144868 77620
rect 143628 77558 144868 77618
rect 143073 77555 143139 77558
rect 144862 77556 144868 77558
rect 144932 77556 144938 77620
rect 145833 77618 145899 77621
rect 145054 77616 145899 77618
rect 145054 77560 145838 77616
rect 145894 77560 145899 77616
rect 145054 77558 145899 77560
rect 140497 77482 140563 77485
rect 139902 77480 140563 77482
rect 139902 77424 140502 77480
rect 140558 77424 140563 77480
rect 139902 77422 140563 77424
rect 138381 77419 138447 77422
rect 138565 77419 138631 77422
rect 140497 77419 140563 77422
rect 144862 77420 144868 77484
rect 144932 77482 144938 77484
rect 145054 77482 145114 77558
rect 145833 77555 145899 77558
rect 145974 77485 146034 77694
rect 146112 77752 146313 77754
rect 146112 77696 146252 77752
rect 146308 77696 146313 77752
rect 146112 77694 146313 77696
rect 146112 77618 146172 77694
rect 146247 77691 146313 77694
rect 146891 77752 146957 77757
rect 146891 77696 146896 77752
rect 146952 77696 146957 77752
rect 146891 77691 146957 77696
rect 148685 77754 148751 77757
rect 148685 77752 148794 77754
rect 148685 77696 148690 77752
rect 148746 77696 148794 77752
rect 148685 77691 148794 77696
rect 146293 77618 146359 77621
rect 146112 77616 146359 77618
rect 146112 77560 146298 77616
rect 146354 77560 146359 77616
rect 146112 77558 146359 77560
rect 146293 77555 146359 77558
rect 146661 77618 146727 77621
rect 146894 77618 146954 77691
rect 147029 77618 147095 77621
rect 146661 77616 146770 77618
rect 146661 77560 146666 77616
rect 146722 77560 146770 77616
rect 146661 77555 146770 77560
rect 146894 77616 147095 77618
rect 146894 77560 147034 77616
rect 147090 77560 147095 77616
rect 146894 77558 147095 77560
rect 147029 77555 147095 77558
rect 148593 77618 148659 77621
rect 148734 77618 148794 77691
rect 148593 77616 148794 77618
rect 148593 77560 148598 77616
rect 148654 77560 148794 77616
rect 148593 77558 148794 77560
rect 149654 77618 149714 77830
rect 150939 77888 151005 77893
rect 150939 77832 150944 77888
rect 151000 77832 151005 77888
rect 150939 77827 151005 77832
rect 151486 77828 151492 77892
rect 151556 77890 151562 77892
rect 151675 77890 151741 77893
rect 152043 77892 152109 77893
rect 151556 77888 151741 77890
rect 151556 77832 151680 77888
rect 151736 77832 151741 77888
rect 151556 77830 151741 77832
rect 151556 77828 151562 77830
rect 151675 77827 151741 77830
rect 152038 77828 152044 77892
rect 152108 77890 152114 77892
rect 152319 77890 152385 77893
rect 152108 77830 152200 77890
rect 152276 77888 152385 77890
rect 152276 77832 152324 77888
rect 152380 77832 152385 77888
rect 152108 77828 152114 77830
rect 152043 77827 152109 77828
rect 152276 77827 152385 77832
rect 152595 77888 152661 77893
rect 152779 77892 152845 77893
rect 153423 77892 153489 77893
rect 153699 77892 153765 77893
rect 154067 77892 154133 77893
rect 152595 77832 152600 77888
rect 152656 77832 152661 77888
rect 152595 77827 152661 77832
rect 152774 77828 152780 77892
rect 152844 77890 152850 77892
rect 153372 77890 153378 77892
rect 152844 77830 152936 77890
rect 153332 77830 153378 77890
rect 153442 77888 153489 77892
rect 153694 77890 153700 77892
rect 153484 77832 153489 77888
rect 152844 77828 152850 77830
rect 153372 77828 153378 77830
rect 153442 77828 153489 77832
rect 153608 77830 153700 77890
rect 153694 77828 153700 77830
rect 153764 77828 153770 77892
rect 154062 77890 154068 77892
rect 153976 77830 154068 77890
rect 154062 77828 154068 77830
rect 154132 77828 154138 77892
rect 154246 77828 154252 77892
rect 154316 77890 154322 77892
rect 154527 77890 154593 77893
rect 154987 77892 155053 77893
rect 154982 77890 154988 77892
rect 154316 77888 154593 77890
rect 154316 77832 154532 77888
rect 154588 77832 154593 77888
rect 154316 77830 154593 77832
rect 154896 77830 154988 77890
rect 154316 77828 154322 77830
rect 152779 77827 152845 77828
rect 153423 77827 153489 77828
rect 153699 77827 153765 77828
rect 154067 77827 154133 77828
rect 154527 77827 154593 77830
rect 154982 77828 154988 77830
rect 155052 77828 155058 77892
rect 155907 77866 155912 77922
rect 155968 77866 155973 77922
rect 155907 77861 155973 77866
rect 156183 77924 156249 77927
rect 157103 77924 157169 77927
rect 156183 77922 156430 77924
rect 156183 77866 156188 77922
rect 156244 77866 156430 77922
rect 157103 77922 157212 77924
rect 156183 77864 156430 77866
rect 156183 77861 156249 77864
rect 154987 77827 155053 77828
rect 150942 77754 151002 77827
rect 151077 77754 151143 77757
rect 150942 77752 151143 77754
rect 150942 77696 151082 77752
rect 151138 77696 151143 77752
rect 150942 77694 151143 77696
rect 152276 77754 152336 77827
rect 152406 77754 152412 77756
rect 152276 77694 152412 77754
rect 151077 77691 151143 77694
rect 152406 77692 152412 77694
rect 152476 77692 152482 77756
rect 152598 77754 152658 77827
rect 152733 77754 152799 77757
rect 152598 77752 152799 77754
rect 152598 77696 152738 77752
rect 152794 77696 152799 77752
rect 152598 77694 152799 77696
rect 152733 77691 152799 77694
rect 152966 77694 155602 77754
rect 152966 77618 153026 77694
rect 153193 77620 153259 77621
rect 149654 77558 153026 77618
rect 148593 77555 148659 77558
rect 153142 77556 153148 77620
rect 153212 77618 153259 77620
rect 154205 77620 154271 77621
rect 154205 77618 154252 77620
rect 153212 77616 153304 77618
rect 153254 77560 153304 77616
rect 153212 77558 153304 77560
rect 154160 77616 154252 77618
rect 154160 77560 154210 77616
rect 154160 77558 154252 77560
rect 153212 77556 153259 77558
rect 153193 77555 153259 77556
rect 154205 77556 154252 77558
rect 154316 77556 154322 77620
rect 154205 77555 154271 77556
rect 145465 77484 145531 77485
rect 144932 77422 145114 77482
rect 144932 77420 144938 77422
rect 145414 77420 145420 77484
rect 145484 77482 145531 77484
rect 145484 77480 145576 77482
rect 145526 77424 145576 77480
rect 145484 77422 145576 77424
rect 145925 77480 146034 77485
rect 145925 77424 145930 77480
rect 145986 77424 146034 77480
rect 145925 77422 146034 77424
rect 146569 77482 146635 77485
rect 146710 77482 146770 77555
rect 146569 77480 146770 77482
rect 146569 77424 146574 77480
rect 146630 77424 146770 77480
rect 146569 77422 146770 77424
rect 149329 77482 149395 77485
rect 155309 77482 155375 77485
rect 149329 77480 155375 77482
rect 149329 77424 149334 77480
rect 149390 77424 155314 77480
rect 155370 77424 155375 77480
rect 149329 77422 155375 77424
rect 155542 77482 155602 77694
rect 155910 77621 155970 77861
rect 156086 77692 156092 77756
rect 156156 77754 156162 77756
rect 156370 77754 156430 77864
rect 156822 77828 156828 77892
rect 156892 77890 156898 77892
rect 157103 77890 157108 77922
rect 156892 77866 157108 77890
rect 157164 77866 157212 77922
rect 157747 77922 157813 77927
rect 156892 77830 157212 77866
rect 157379 77888 157445 77893
rect 157379 77832 157384 77888
rect 157440 77832 157445 77888
rect 157747 77866 157752 77922
rect 157808 77866 157813 77922
rect 162715 77922 162781 77927
rect 157747 77861 157813 77866
rect 156892 77828 156898 77830
rect 157379 77827 157445 77832
rect 157382 77757 157442 77827
rect 156156 77694 156430 77754
rect 156156 77692 156162 77694
rect 156638 77692 156644 77756
rect 156708 77754 156714 77756
rect 157241 77754 157307 77757
rect 156708 77752 157307 77754
rect 156708 77696 157246 77752
rect 157302 77696 157307 77752
rect 156708 77694 157307 77696
rect 157382 77752 157491 77757
rect 157382 77696 157430 77752
rect 157486 77696 157491 77752
rect 157382 77694 157491 77696
rect 157750 77754 157810 77861
rect 158110 77828 158116 77892
rect 158180 77890 158186 77892
rect 158483 77890 158549 77893
rect 158667 77892 158733 77893
rect 158180 77888 158549 77890
rect 158180 77832 158488 77888
rect 158544 77832 158549 77888
rect 158180 77830 158549 77832
rect 158180 77828 158186 77830
rect 158483 77827 158549 77830
rect 158662 77828 158668 77892
rect 158732 77890 158738 77892
rect 162158 77890 162164 77892
rect 158732 77830 158824 77890
rect 159038 77830 162164 77890
rect 158732 77828 158738 77830
rect 158667 77827 158733 77828
rect 157885 77754 157951 77757
rect 158529 77756 158595 77757
rect 158478 77754 158484 77756
rect 157750 77752 157951 77754
rect 157750 77696 157890 77752
rect 157946 77696 157951 77752
rect 157750 77694 157951 77696
rect 158438 77694 158484 77754
rect 158548 77752 158595 77756
rect 158590 77696 158595 77752
rect 156708 77692 156714 77694
rect 157241 77691 157307 77694
rect 157425 77691 157491 77694
rect 157885 77691 157951 77694
rect 158478 77692 158484 77694
rect 158548 77692 158595 77696
rect 158529 77691 158595 77692
rect 155910 77616 156019 77621
rect 155910 77560 155958 77616
rect 156014 77560 156019 77616
rect 155910 77558 156019 77560
rect 155953 77555 156019 77558
rect 156270 77556 156276 77620
rect 156340 77618 156346 77620
rect 156689 77618 156755 77621
rect 156340 77616 156755 77618
rect 156340 77560 156694 77616
rect 156750 77560 156755 77616
rect 156340 77558 156755 77560
rect 156340 77556 156346 77558
rect 156689 77555 156755 77558
rect 158253 77620 158319 77621
rect 158253 77616 158300 77620
rect 158364 77618 158370 77620
rect 158253 77560 158258 77616
rect 158253 77556 158300 77560
rect 158364 77558 158410 77618
rect 158364 77556 158370 77558
rect 158253 77555 158319 77556
rect 159038 77482 159098 77830
rect 162158 77828 162164 77830
rect 162228 77828 162234 77892
rect 162347 77888 162413 77893
rect 162715 77892 162720 77922
rect 162776 77892 162781 77922
rect 164003 77922 164069 77927
rect 163083 77892 163149 77893
rect 162347 77832 162352 77888
rect 162408 77832 162413 77888
rect 162347 77827 162413 77832
rect 162710 77828 162716 77892
rect 162780 77890 162786 77892
rect 163078 77890 163084 77892
rect 162780 77830 162838 77890
rect 162992 77830 163084 77890
rect 162780 77828 162786 77830
rect 163078 77828 163084 77830
rect 163148 77828 163154 77892
rect 163262 77828 163268 77892
rect 163332 77890 163338 77892
rect 163451 77890 163517 77893
rect 163332 77888 163517 77890
rect 163332 77832 163456 77888
rect 163512 77832 163517 77888
rect 163332 77830 163517 77832
rect 163332 77828 163338 77830
rect 163083 77827 163149 77828
rect 163451 77827 163517 77830
rect 163630 77828 163636 77892
rect 163700 77890 163706 77892
rect 164003 77890 164008 77922
rect 163700 77866 164008 77890
rect 164064 77866 164069 77922
rect 164831 77924 164897 77927
rect 164831 77922 164940 77924
rect 163700 77861 164069 77866
rect 164187 77890 164253 77893
rect 164366 77890 164372 77892
rect 164187 77888 164372 77890
rect 163700 77830 164066 77861
rect 164187 77832 164192 77888
rect 164248 77832 164372 77888
rect 164187 77830 164372 77832
rect 163700 77828 163706 77830
rect 164187 77827 164253 77830
rect 164366 77828 164372 77830
rect 164436 77828 164442 77892
rect 164831 77866 164836 77922
rect 164892 77892 164940 77922
rect 165475 77922 165541 77927
rect 164892 77866 164924 77892
rect 164831 77861 164924 77866
rect 164880 77830 164924 77861
rect 164918 77828 164924 77830
rect 164988 77828 164994 77892
rect 165102 77828 165108 77892
rect 165172 77890 165178 77892
rect 165291 77890 165357 77893
rect 165475 77892 165480 77922
rect 165536 77892 165541 77922
rect 165843 77892 165909 77893
rect 165172 77888 165357 77890
rect 165172 77832 165296 77888
rect 165352 77832 165357 77888
rect 165172 77830 165357 77832
rect 165172 77828 165178 77830
rect 165291 77827 165357 77830
rect 165470 77828 165476 77892
rect 165540 77890 165546 77892
rect 165838 77890 165844 77892
rect 165540 77830 165598 77890
rect 165752 77830 165844 77890
rect 165540 77828 165546 77830
rect 165838 77828 165844 77830
rect 165908 77828 165914 77892
rect 166758 77828 166764 77892
rect 166828 77890 166834 77892
rect 166947 77890 167013 77893
rect 166828 77888 167013 77890
rect 166828 77832 166952 77888
rect 167008 77832 167013 77888
rect 166828 77830 167013 77832
rect 167088 77890 167148 77966
rect 167310 77964 167316 77966
rect 167380 77964 167386 78028
rect 167678 77964 167684 78028
rect 167748 77964 167754 78028
rect 168330 77966 169770 78026
rect 167499 77922 167565 77927
rect 167223 77890 167289 77893
rect 167499 77892 167504 77922
rect 167560 77892 167565 77922
rect 167088 77888 167289 77890
rect 167088 77832 167228 77888
rect 167284 77832 167289 77888
rect 167088 77830 167289 77832
rect 166828 77828 166834 77830
rect 165843 77827 165909 77828
rect 166947 77827 167013 77830
rect 167223 77827 167289 77830
rect 167494 77828 167500 77892
rect 167564 77890 167570 77892
rect 167686 77890 167746 77964
rect 168051 77890 168117 77893
rect 167564 77830 167622 77890
rect 167686 77888 168117 77890
rect 167686 77832 168056 77888
rect 168112 77832 168117 77888
rect 167686 77830 168117 77832
rect 167564 77828 167570 77830
rect 168051 77827 168117 77830
rect 159219 77752 159285 77757
rect 159219 77696 159224 77752
rect 159280 77696 159285 77752
rect 159219 77691 159285 77696
rect 159725 77754 159791 77757
rect 160691 77756 160757 77757
rect 160318 77754 160324 77756
rect 159725 77752 160324 77754
rect 159725 77696 159730 77752
rect 159786 77696 160324 77752
rect 159725 77694 160324 77696
rect 159725 77691 159791 77694
rect 160318 77692 160324 77694
rect 160388 77692 160394 77756
rect 160686 77692 160692 77756
rect 160756 77754 160762 77756
rect 161238 77754 161244 77756
rect 160756 77694 160848 77754
rect 161062 77723 161244 77754
rect 161013 77718 161244 77723
rect 160756 77692 160762 77694
rect 160691 77691 160757 77692
rect 159222 77618 159282 77691
rect 161013 77662 161018 77718
rect 161074 77694 161244 77718
rect 161074 77662 161122 77694
rect 161238 77692 161244 77694
rect 161308 77692 161314 77756
rect 161013 77660 161122 77662
rect 161013 77657 161079 77660
rect 160461 77618 160527 77621
rect 159222 77616 160527 77618
rect 159222 77560 160466 77616
rect 160522 77560 160527 77616
rect 159222 77558 160527 77560
rect 160461 77555 160527 77558
rect 161473 77618 161539 77621
rect 162350 77618 162410 77827
rect 162577 77754 162643 77757
rect 162710 77754 162716 77756
rect 162577 77752 162716 77754
rect 162577 77696 162582 77752
rect 162638 77696 162716 77752
rect 162577 77694 162716 77696
rect 162577 77691 162643 77694
rect 162710 77692 162716 77694
rect 162780 77692 162786 77756
rect 163814 77692 163820 77756
rect 163884 77754 163890 77756
rect 168330 77754 168390 77966
rect 168603 77892 168669 77893
rect 168598 77890 168604 77892
rect 168512 77830 168604 77890
rect 168598 77828 168604 77830
rect 168668 77828 168674 77892
rect 169155 77890 169221 77893
rect 169112 77888 169221 77890
rect 169112 77832 169160 77888
rect 169216 77832 169221 77888
rect 168603 77827 168669 77828
rect 169112 77827 169221 77832
rect 169339 77888 169405 77893
rect 169339 77832 169344 77888
rect 169400 77832 169405 77888
rect 169339 77827 169405 77832
rect 169523 77888 169589 77893
rect 169523 77832 169528 77888
rect 169584 77832 169589 77888
rect 169523 77827 169589 77832
rect 163884 77694 168390 77754
rect 163884 77692 163890 77694
rect 169112 77621 169172 77827
rect 169342 77621 169402 77827
rect 169526 77621 169586 77827
rect 161473 77616 162410 77618
rect 161473 77560 161478 77616
rect 161534 77560 162410 77616
rect 161473 77558 162410 77560
rect 164417 77618 164483 77621
rect 164550 77618 164556 77620
rect 164417 77616 164556 77618
rect 164417 77560 164422 77616
rect 164478 77560 164556 77616
rect 164417 77558 164556 77560
rect 161473 77555 161539 77558
rect 164417 77555 164483 77558
rect 164550 77556 164556 77558
rect 164620 77556 164626 77620
rect 166022 77556 166028 77620
rect 166092 77618 166098 77620
rect 166165 77618 166231 77621
rect 166092 77616 166231 77618
rect 166092 77560 166170 77616
rect 166226 77560 166231 77616
rect 166092 77558 166231 77560
rect 166092 77556 166098 77558
rect 166165 77555 166231 77558
rect 166574 77556 166580 77620
rect 166644 77618 166650 77620
rect 166901 77618 166967 77621
rect 166644 77616 166967 77618
rect 166644 77560 166906 77616
rect 166962 77560 166967 77616
rect 166644 77558 166967 77560
rect 166644 77556 166650 77558
rect 166901 77555 166967 77558
rect 168373 77618 168439 77621
rect 168557 77618 168623 77621
rect 168373 77616 168623 77618
rect 168373 77560 168378 77616
rect 168434 77560 168562 77616
rect 168618 77560 168623 77616
rect 168373 77558 168623 77560
rect 168373 77555 168439 77558
rect 168557 77555 168623 77558
rect 169109 77616 169175 77621
rect 169109 77560 169114 77616
rect 169170 77560 169175 77616
rect 169109 77555 169175 77560
rect 169293 77616 169402 77621
rect 169293 77560 169298 77616
rect 169354 77560 169402 77616
rect 169293 77558 169402 77560
rect 169477 77616 169586 77621
rect 169477 77560 169482 77616
rect 169538 77560 169586 77616
rect 169477 77558 169586 77560
rect 169710 77618 169770 77966
rect 170259 77922 170325 77927
rect 170075 77892 170141 77893
rect 170259 77892 170264 77922
rect 170320 77892 170325 77922
rect 172375 77924 172441 77927
rect 172375 77922 172484 77924
rect 170627 77892 170693 77893
rect 170995 77892 171061 77893
rect 170070 77890 170076 77892
rect 169984 77830 170076 77890
rect 170070 77828 170076 77830
rect 170140 77828 170146 77892
rect 170254 77828 170260 77892
rect 170324 77890 170330 77892
rect 170622 77890 170628 77892
rect 170324 77830 170382 77890
rect 170536 77830 170628 77890
rect 170324 77828 170330 77830
rect 170622 77828 170628 77830
rect 170692 77828 170698 77892
rect 170990 77890 170996 77892
rect 170904 77830 170996 77890
rect 170990 77828 170996 77830
rect 171060 77828 171066 77892
rect 171639 77890 171705 77893
rect 171910 77890 171916 77892
rect 171639 77888 171916 77890
rect 171639 77832 171644 77888
rect 171700 77832 171916 77888
rect 171639 77830 171916 77832
rect 170075 77827 170141 77828
rect 170627 77827 170693 77828
rect 170995 77827 171061 77828
rect 171639 77827 171705 77830
rect 171910 77828 171916 77830
rect 171980 77828 171986 77892
rect 172191 77890 172257 77893
rect 172056 77888 172257 77890
rect 172056 77832 172196 77888
rect 172252 77832 172257 77888
rect 172375 77866 172380 77922
rect 172436 77892 172484 77922
rect 172436 77866 172468 77892
rect 172375 77861 172468 77866
rect 172056 77830 172257 77832
rect 172424 77830 172468 77861
rect 170443 77754 170509 77757
rect 170806 77754 170812 77756
rect 170443 77752 170812 77754
rect 170443 77696 170448 77752
rect 170504 77696 170812 77752
rect 170443 77694 170812 77696
rect 170443 77691 170509 77694
rect 170806 77692 170812 77694
rect 170876 77692 170882 77756
rect 172056 77754 172116 77830
rect 172191 77827 172257 77830
rect 172462 77828 172468 77830
rect 172532 77828 172538 77892
rect 172743 77890 172809 77893
rect 173014 77890 173020 77892
rect 172743 77888 173020 77890
rect 172743 77832 172748 77888
rect 172804 77832 173020 77888
rect 172743 77830 173020 77832
rect 172743 77827 172809 77830
rect 173014 77828 173020 77830
rect 173084 77828 173090 77892
rect 173206 77890 173266 78238
rect 173479 77890 173545 77893
rect 173206 77888 173545 77890
rect 173206 77832 173484 77888
rect 173540 77832 173545 77888
rect 173206 77830 173545 77832
rect 173479 77827 173545 77830
rect 173847 77890 173913 77893
rect 174353 77890 174419 77893
rect 173847 77888 174419 77890
rect 173847 77832 173852 77888
rect 173908 77832 174358 77888
rect 174414 77832 174419 77888
rect 173847 77830 174419 77832
rect 173847 77827 173913 77830
rect 174353 77827 174419 77830
rect 176285 77890 176351 77893
rect 181437 77890 181503 77893
rect 176285 77888 181503 77890
rect 176285 77832 176290 77888
rect 176346 77832 181442 77888
rect 181498 77832 181503 77888
rect 176285 77830 181503 77832
rect 176285 77827 176351 77830
rect 181437 77827 181503 77830
rect 175641 77754 175707 77757
rect 172056 77752 175707 77754
rect 172056 77696 175646 77752
rect 175702 77696 175707 77752
rect 172056 77694 175707 77696
rect 175641 77691 175707 77694
rect 175825 77754 175891 77757
rect 396574 77754 396580 77756
rect 175825 77752 396580 77754
rect 175825 77696 175830 77752
rect 175886 77696 396580 77752
rect 175825 77694 396580 77696
rect 175825 77691 175891 77694
rect 396574 77692 396580 77694
rect 396644 77692 396650 77756
rect 173341 77618 173407 77621
rect 173617 77620 173683 77621
rect 173566 77618 173572 77620
rect 169710 77616 173407 77618
rect 169710 77560 173346 77616
rect 173402 77560 173407 77616
rect 169710 77558 173407 77560
rect 173526 77558 173572 77618
rect 173636 77616 173683 77620
rect 173678 77560 173683 77616
rect 169293 77555 169359 77558
rect 169477 77555 169543 77558
rect 173341 77555 173407 77558
rect 173566 77556 173572 77558
rect 173636 77556 173683 77560
rect 173617 77555 173683 77556
rect 175825 77618 175891 77621
rect 396809 77618 396875 77621
rect 175825 77616 396875 77618
rect 175825 77560 175830 77616
rect 175886 77560 396814 77616
rect 396870 77560 396875 77616
rect 175825 77558 396875 77560
rect 175825 77555 175891 77558
rect 396809 77555 396875 77558
rect 155542 77422 159098 77482
rect 159541 77482 159607 77485
rect 162945 77482 163011 77485
rect 159541 77480 163011 77482
rect 159541 77424 159546 77480
rect 159602 77424 162950 77480
rect 163006 77424 163011 77480
rect 159541 77422 163011 77424
rect 145484 77420 145531 77422
rect 145465 77419 145531 77420
rect 145925 77419 145991 77422
rect 146569 77419 146635 77422
rect 149329 77419 149395 77422
rect 155309 77419 155375 77422
rect 159541 77419 159607 77422
rect 162945 77419 163011 77422
rect 164233 77482 164299 77485
rect 164366 77482 164372 77484
rect 164233 77480 164372 77482
rect 164233 77424 164238 77480
rect 164294 77424 164372 77480
rect 164233 77422 164372 77424
rect 164233 77419 164299 77422
rect 164366 77420 164372 77422
rect 164436 77420 164442 77484
rect 164877 77482 164943 77485
rect 165286 77482 165292 77484
rect 164877 77480 165292 77482
rect 164877 77424 164882 77480
rect 164938 77424 165292 77480
rect 164877 77422 165292 77424
rect 164877 77419 164943 77422
rect 165286 77420 165292 77422
rect 165356 77420 165362 77484
rect 165889 77482 165955 77485
rect 166441 77482 166507 77485
rect 165889 77480 166507 77482
rect 165889 77424 165894 77480
rect 165950 77424 166446 77480
rect 166502 77424 166507 77480
rect 165889 77422 166507 77424
rect 165889 77419 165955 77422
rect 166441 77419 166507 77422
rect 166993 77482 167059 77485
rect 166993 77480 168390 77482
rect 166993 77424 166998 77480
rect 167054 77424 168390 77480
rect 166993 77422 168390 77424
rect 166993 77419 167059 77422
rect 134149 77346 134215 77349
rect 138565 77346 138631 77349
rect 134149 77344 138631 77346
rect 134149 77288 134154 77344
rect 134210 77288 138570 77344
rect 138626 77288 138631 77344
rect 134149 77286 138631 77288
rect 134149 77283 134215 77286
rect 138565 77283 138631 77286
rect 144545 77346 144611 77349
rect 149053 77346 149119 77349
rect 144545 77344 149119 77346
rect 144545 77288 144550 77344
rect 144606 77288 149058 77344
rect 149114 77288 149119 77344
rect 144545 77286 149119 77288
rect 144545 77283 144611 77286
rect 149053 77283 149119 77286
rect 150433 77346 150499 77349
rect 167545 77346 167611 77349
rect 150433 77344 167611 77346
rect 150433 77288 150438 77344
rect 150494 77288 167550 77344
rect 167606 77288 167611 77344
rect 150433 77286 167611 77288
rect 168330 77346 168390 77422
rect 169334 77420 169340 77484
rect 169404 77482 169410 77484
rect 171961 77482 172027 77485
rect 172145 77484 172211 77485
rect 169404 77480 172027 77482
rect 169404 77424 171966 77480
rect 172022 77424 172027 77480
rect 169404 77422 172027 77424
rect 169404 77420 169410 77422
rect 171961 77419 172027 77422
rect 172094 77420 172100 77484
rect 172164 77482 172211 77484
rect 172421 77482 172487 77485
rect 175825 77482 175891 77485
rect 181437 77482 181503 77485
rect 396993 77482 397059 77485
rect 172164 77480 172256 77482
rect 172206 77424 172256 77480
rect 172164 77422 172256 77424
rect 172421 77480 175520 77482
rect 172421 77424 172426 77480
rect 172482 77424 175520 77480
rect 172421 77422 175520 77424
rect 172164 77420 172211 77422
rect 172145 77419 172211 77420
rect 172421 77419 172487 77422
rect 171133 77346 171199 77349
rect 171501 77348 171567 77349
rect 171501 77346 171548 77348
rect 168330 77344 171199 77346
rect 168330 77288 171138 77344
rect 171194 77288 171199 77344
rect 168330 77286 171199 77288
rect 171456 77344 171548 77346
rect 171456 77288 171506 77344
rect 171456 77286 171548 77288
rect 150433 77283 150499 77286
rect 167545 77283 167611 77286
rect 171133 77283 171199 77286
rect 171501 77284 171548 77286
rect 171612 77284 171618 77348
rect 172053 77346 172119 77349
rect 172973 77346 173039 77349
rect 172053 77344 173039 77346
rect 172053 77288 172058 77344
rect 172114 77288 172978 77344
rect 173034 77288 173039 77344
rect 172053 77286 173039 77288
rect 175460 77346 175520 77422
rect 175825 77480 180810 77482
rect 175825 77424 175830 77480
rect 175886 77424 180810 77480
rect 175825 77422 180810 77424
rect 175825 77419 175891 77422
rect 180750 77346 180810 77422
rect 181437 77480 397059 77482
rect 181437 77424 181442 77480
rect 181498 77424 396998 77480
rect 397054 77424 397059 77480
rect 181437 77422 397059 77424
rect 181437 77419 181503 77422
rect 396993 77419 397059 77422
rect 527173 77346 527239 77349
rect 175460 77286 179430 77346
rect 180750 77344 527239 77346
rect 180750 77288 527178 77344
rect 527234 77288 527239 77344
rect 180750 77286 527239 77288
rect 171501 77283 171567 77284
rect 172053 77283 172119 77286
rect 172973 77283 173039 77286
rect 124765 77210 124831 77213
rect 129273 77210 129339 77213
rect 132493 77212 132559 77213
rect 132493 77210 132540 77212
rect 124765 77208 129339 77210
rect 124765 77152 124770 77208
rect 124826 77152 129278 77208
rect 129334 77152 129339 77208
rect 124765 77150 129339 77152
rect 132448 77208 132540 77210
rect 132448 77152 132498 77208
rect 132448 77150 132540 77152
rect 124765 77147 124831 77150
rect 129273 77147 129339 77150
rect 132493 77148 132540 77150
rect 132604 77148 132610 77212
rect 139577 77210 139643 77213
rect 153837 77212 153903 77213
rect 153510 77210 153516 77212
rect 139577 77208 153516 77210
rect 139577 77152 139582 77208
rect 139638 77152 153516 77208
rect 139577 77150 153516 77152
rect 132493 77147 132559 77148
rect 139577 77147 139643 77150
rect 153510 77148 153516 77150
rect 153580 77148 153586 77212
rect 153837 77210 153884 77212
rect 153792 77208 153884 77210
rect 153792 77152 153842 77208
rect 153792 77150 153884 77152
rect 153837 77148 153884 77150
rect 153948 77148 153954 77212
rect 163037 77210 163103 77213
rect 154070 77208 163103 77210
rect 154070 77152 163042 77208
rect 163098 77152 163103 77208
rect 154070 77150 163103 77152
rect 153837 77147 153903 77148
rect 143625 77074 143691 77077
rect 154070 77074 154130 77150
rect 163037 77147 163103 77150
rect 167085 77210 167151 77213
rect 168005 77210 168071 77213
rect 167085 77208 168071 77210
rect 167085 77152 167090 77208
rect 167146 77152 168010 77208
rect 168066 77152 168071 77208
rect 167085 77150 168071 77152
rect 167085 77147 167151 77150
rect 168005 77147 168071 77150
rect 170990 77148 170996 77212
rect 171060 77210 171066 77212
rect 178401 77210 178467 77213
rect 171060 77208 178467 77210
rect 171060 77152 178406 77208
rect 178462 77152 178467 77208
rect 171060 77150 178467 77152
rect 179370 77210 179430 77286
rect 527173 77283 527239 77286
rect 397453 77210 397519 77213
rect 179370 77208 397519 77210
rect 179370 77152 397458 77208
rect 397514 77152 397519 77208
rect 179370 77150 397519 77152
rect 171060 77148 171066 77150
rect 178401 77147 178467 77150
rect 397453 77147 397519 77150
rect 143625 77072 154130 77074
rect 143625 77016 143630 77072
rect 143686 77016 154130 77072
rect 143625 77014 154130 77016
rect 154849 77074 154915 77077
rect 154982 77074 154988 77076
rect 154849 77072 154988 77074
rect 154849 77016 154854 77072
rect 154910 77016 154988 77072
rect 154849 77014 154988 77016
rect 143625 77011 143691 77014
rect 154849 77011 154915 77014
rect 154982 77012 154988 77014
rect 155052 77012 155058 77076
rect 156086 77012 156092 77076
rect 156156 77074 156162 77076
rect 156321 77074 156387 77077
rect 156156 77072 156387 77074
rect 156156 77016 156326 77072
rect 156382 77016 156387 77072
rect 156156 77014 156387 77016
rect 156156 77012 156162 77014
rect 156321 77011 156387 77014
rect 158529 77074 158595 77077
rect 159541 77074 159607 77077
rect 158529 77072 159607 77074
rect 158529 77016 158534 77072
rect 158590 77016 159546 77072
rect 159602 77016 159607 77072
rect 158529 77014 159607 77016
rect 158529 77011 158595 77014
rect 159541 77011 159607 77014
rect 164918 77012 164924 77076
rect 164988 77074 164994 77076
rect 165337 77074 165403 77077
rect 164988 77072 165403 77074
rect 164988 77016 165342 77072
rect 165398 77016 165403 77072
rect 164988 77014 165403 77016
rect 164988 77012 164994 77014
rect 165337 77011 165403 77014
rect 166390 77012 166396 77076
rect 166460 77074 166466 77076
rect 166625 77074 166691 77077
rect 166460 77072 166691 77074
rect 166460 77016 166630 77072
rect 166686 77016 166691 77072
rect 166460 77014 166691 77016
rect 166460 77012 166466 77014
rect 166625 77011 166691 77014
rect 166901 77074 166967 77077
rect 167085 77074 167151 77077
rect 166901 77072 167151 77074
rect 166901 77016 166906 77072
rect 166962 77016 167090 77072
rect 167146 77016 167151 77072
rect 166901 77014 167151 77016
rect 166901 77011 166967 77014
rect 167085 77011 167151 77014
rect 171593 77074 171659 77077
rect 176285 77074 176351 77077
rect 396717 77074 396783 77077
rect 171593 77072 176351 77074
rect 171593 77016 171598 77072
rect 171654 77016 176290 77072
rect 176346 77016 176351 77072
rect 171593 77014 176351 77016
rect 171593 77011 171659 77014
rect 176285 77011 176351 77014
rect 186270 77072 396783 77074
rect 186270 77016 396722 77072
rect 396778 77016 396783 77072
rect 186270 77014 396783 77016
rect 3969 76938 4035 76941
rect 173525 76938 173591 76941
rect 3969 76936 173591 76938
rect 3969 76880 3974 76936
rect 4030 76880 173530 76936
rect 173586 76880 173591 76936
rect 3969 76878 173591 76880
rect 3969 76875 4035 76878
rect 173525 76875 173591 76878
rect 127249 76804 127315 76805
rect 127198 76802 127204 76804
rect 127158 76742 127204 76802
rect 127268 76800 127315 76804
rect 127310 76744 127315 76800
rect 127198 76740 127204 76742
rect 127268 76740 127315 76744
rect 127249 76739 127315 76740
rect 128445 76802 128511 76805
rect 147305 76804 147371 76805
rect 129038 76802 129044 76804
rect 128445 76800 129044 76802
rect 128445 76744 128450 76800
rect 128506 76744 129044 76800
rect 128445 76742 129044 76744
rect 128445 76739 128511 76742
rect 129038 76740 129044 76742
rect 129108 76740 129114 76804
rect 147254 76802 147260 76804
rect 147214 76742 147260 76802
rect 147324 76800 147371 76804
rect 147366 76744 147371 76800
rect 147254 76740 147260 76742
rect 147324 76740 147371 76744
rect 147305 76739 147371 76740
rect 153193 76802 153259 76805
rect 153326 76802 153332 76804
rect 153193 76800 153332 76802
rect 153193 76744 153198 76800
rect 153254 76744 153332 76800
rect 153193 76742 153332 76744
rect 153193 76739 153259 76742
rect 153326 76740 153332 76742
rect 153396 76740 153402 76804
rect 154113 76802 154179 76805
rect 155677 76804 155743 76805
rect 154430 76802 154436 76804
rect 154113 76800 154436 76802
rect 154113 76744 154118 76800
rect 154174 76744 154436 76800
rect 154113 76742 154436 76744
rect 154113 76739 154179 76742
rect 154430 76740 154436 76742
rect 154500 76740 154506 76804
rect 155677 76800 155724 76804
rect 155788 76802 155794 76804
rect 162669 76802 162735 76805
rect 165521 76802 165587 76805
rect 155677 76744 155682 76800
rect 155677 76740 155724 76744
rect 155788 76742 155834 76802
rect 162669 76800 165587 76802
rect 162669 76744 162674 76800
rect 162730 76744 165526 76800
rect 165582 76744 165587 76800
rect 162669 76742 165587 76744
rect 155788 76740 155794 76742
rect 155677 76739 155743 76740
rect 162669 76739 162735 76742
rect 165521 76739 165587 76742
rect 166901 76802 166967 76805
rect 168097 76804 168163 76805
rect 167494 76802 167500 76804
rect 166901 76800 167500 76802
rect 166901 76744 166906 76800
rect 166962 76744 167500 76800
rect 166901 76742 167500 76744
rect 166901 76739 166967 76742
rect 167494 76740 167500 76742
rect 167564 76740 167570 76804
rect 168046 76802 168052 76804
rect 168006 76742 168052 76802
rect 168116 76800 168163 76804
rect 168158 76744 168163 76800
rect 168046 76740 168052 76742
rect 168116 76740 168163 76744
rect 168097 76739 168163 76740
rect 171777 76802 171843 76805
rect 186270 76802 186330 77014
rect 396717 77011 396783 77014
rect 171777 76800 186330 76802
rect 171777 76744 171782 76800
rect 171838 76744 186330 76800
rect 171777 76742 186330 76744
rect 171777 76739 171843 76742
rect 3785 76666 3851 76669
rect 173433 76666 173499 76669
rect 3785 76664 173499 76666
rect 3785 76608 3790 76664
rect 3846 76608 173438 76664
rect 173494 76608 173499 76664
rect 3785 76606 173499 76608
rect 3785 76603 3851 76606
rect 173433 76603 173499 76606
rect 3509 76530 3575 76533
rect 173157 76530 173223 76533
rect 3509 76528 173223 76530
rect 3509 76472 3514 76528
rect 3570 76472 173162 76528
rect 173218 76472 173223 76528
rect 3509 76470 173223 76472
rect 3509 76467 3575 76470
rect 173157 76467 173223 76470
rect 127065 76394 127131 76397
rect 127382 76394 127388 76396
rect 127065 76392 127388 76394
rect 127065 76336 127070 76392
rect 127126 76336 127388 76392
rect 127065 76334 127388 76336
rect 127065 76331 127131 76334
rect 127382 76332 127388 76334
rect 127452 76332 127458 76396
rect 128445 76394 128511 76397
rect 129733 76396 129799 76397
rect 130009 76396 130075 76397
rect 128670 76394 128676 76396
rect 128445 76392 128676 76394
rect 128445 76336 128450 76392
rect 128506 76336 128676 76392
rect 128445 76334 128676 76336
rect 128445 76331 128511 76334
rect 128670 76332 128676 76334
rect 128740 76332 128746 76396
rect 129733 76394 129780 76396
rect 129688 76392 129780 76394
rect 129688 76336 129738 76392
rect 129688 76334 129780 76336
rect 129733 76332 129780 76334
rect 129844 76332 129850 76396
rect 129958 76394 129964 76396
rect 129918 76334 129964 76394
rect 130028 76392 130075 76396
rect 130070 76336 130075 76392
rect 129958 76332 129964 76334
rect 130028 76332 130075 76336
rect 129733 76331 129799 76332
rect 130009 76331 130075 76332
rect 132585 76394 132651 76397
rect 134333 76396 134399 76397
rect 139025 76396 139091 76397
rect 132902 76394 132908 76396
rect 132585 76392 132908 76394
rect 132585 76336 132590 76392
rect 132646 76336 132908 76392
rect 132585 76334 132908 76336
rect 132585 76331 132651 76334
rect 132902 76332 132908 76334
rect 132972 76332 132978 76396
rect 134333 76392 134380 76396
rect 134444 76394 134450 76396
rect 138974 76394 138980 76396
rect 134333 76336 134338 76392
rect 134333 76332 134380 76336
rect 134444 76334 134490 76394
rect 138934 76334 138980 76394
rect 139044 76392 139091 76396
rect 139086 76336 139091 76392
rect 134444 76332 134450 76334
rect 138974 76332 138980 76334
rect 139044 76332 139091 76336
rect 139158 76332 139164 76396
rect 139228 76394 139234 76396
rect 139301 76394 139367 76397
rect 139228 76392 139367 76394
rect 139228 76336 139306 76392
rect 139362 76336 139367 76392
rect 139228 76334 139367 76336
rect 139228 76332 139234 76334
rect 134333 76331 134399 76332
rect 139025 76331 139091 76332
rect 139301 76331 139367 76334
rect 145598 76332 145604 76396
rect 145668 76394 145674 76396
rect 146109 76394 146175 76397
rect 145668 76392 146175 76394
rect 145668 76336 146114 76392
rect 146170 76336 146175 76392
rect 145668 76334 146175 76336
rect 145668 76332 145674 76334
rect 146109 76331 146175 76334
rect 153326 76332 153332 76396
rect 153396 76394 153402 76396
rect 154021 76394 154087 76397
rect 162577 76396 162643 76397
rect 162526 76394 162532 76396
rect 153396 76392 154087 76394
rect 153396 76336 154026 76392
rect 154082 76336 154087 76392
rect 153396 76334 154087 76336
rect 162486 76334 162532 76394
rect 162596 76392 162643 76396
rect 162638 76336 162643 76392
rect 153396 76332 153402 76334
rect 154021 76331 154087 76334
rect 162526 76332 162532 76334
rect 162596 76332 162643 76336
rect 167494 76332 167500 76396
rect 167564 76394 167570 76396
rect 168281 76394 168347 76397
rect 167564 76392 168347 76394
rect 167564 76336 168286 76392
rect 168342 76336 168347 76392
rect 167564 76334 168347 76336
rect 167564 76332 167570 76334
rect 162577 76331 162643 76332
rect 168281 76331 168347 76334
rect 168465 76394 168531 76397
rect 168598 76394 168604 76396
rect 168465 76392 168604 76394
rect 168465 76336 168470 76392
rect 168526 76336 168604 76392
rect 168465 76334 168604 76336
rect 168465 76331 168531 76334
rect 168598 76332 168604 76334
rect 168668 76332 168674 76396
rect 169334 76332 169340 76396
rect 169404 76394 169410 76396
rect 169661 76394 169727 76397
rect 169404 76392 169727 76394
rect 169404 76336 169666 76392
rect 169722 76336 169727 76392
rect 169404 76334 169727 76336
rect 169404 76332 169410 76334
rect 169661 76331 169727 76334
rect 171358 76332 171364 76396
rect 171428 76394 171434 76396
rect 173065 76394 173131 76397
rect 171428 76392 173131 76394
rect 171428 76336 173070 76392
rect 173126 76336 173131 76392
rect 171428 76334 173131 76336
rect 171428 76332 171434 76334
rect 173065 76331 173131 76334
rect 132861 76258 132927 76261
rect 133086 76258 133092 76260
rect 132861 76256 133092 76258
rect 132861 76200 132866 76256
rect 132922 76200 133092 76256
rect 132861 76198 133092 76200
rect 132861 76195 132927 76198
rect 133086 76196 133092 76198
rect 133156 76196 133162 76260
rect 145414 76196 145420 76260
rect 145484 76258 145490 76260
rect 145833 76258 145899 76261
rect 145484 76256 145899 76258
rect 145484 76200 145838 76256
rect 145894 76200 145899 76256
rect 145484 76198 145899 76200
rect 145484 76196 145490 76198
rect 145833 76195 145899 76198
rect 149830 76196 149836 76260
rect 149900 76258 149906 76260
rect 150157 76258 150223 76261
rect 149900 76256 150223 76258
rect 149900 76200 150162 76256
rect 150218 76200 150223 76256
rect 149900 76198 150223 76200
rect 149900 76196 149906 76198
rect 150157 76195 150223 76198
rect 153653 76258 153719 76261
rect 154062 76258 154068 76260
rect 153653 76256 154068 76258
rect 153653 76200 153658 76256
rect 153714 76200 154068 76256
rect 153653 76198 154068 76200
rect 153653 76195 153719 76198
rect 154062 76196 154068 76198
rect 154132 76196 154138 76260
rect 162342 76196 162348 76260
rect 162412 76258 162418 76260
rect 162485 76258 162551 76261
rect 162412 76256 162551 76258
rect 162412 76200 162490 76256
rect 162546 76200 162551 76256
rect 162412 76198 162551 76200
rect 162412 76196 162418 76198
rect 162485 76195 162551 76198
rect 163446 76196 163452 76260
rect 163516 76258 163522 76260
rect 164049 76258 164115 76261
rect 163516 76256 164115 76258
rect 163516 76200 164054 76256
rect 164110 76200 164115 76256
rect 163516 76198 164115 76200
rect 163516 76196 163522 76198
rect 164049 76195 164115 76198
rect 166206 76196 166212 76260
rect 166276 76258 166282 76260
rect 166717 76258 166783 76261
rect 166276 76256 166783 76258
rect 166276 76200 166722 76256
rect 166778 76200 166783 76256
rect 166276 76198 166783 76200
rect 166276 76196 166282 76198
rect 166717 76195 166783 76198
rect 167269 76258 167335 76261
rect 167545 76258 167611 76261
rect 172973 76260 173039 76261
rect 172973 76258 173020 76260
rect 167269 76256 167611 76258
rect 167269 76200 167274 76256
rect 167330 76200 167550 76256
rect 167606 76200 167611 76256
rect 167269 76198 167611 76200
rect 172928 76256 173020 76258
rect 172928 76200 172978 76256
rect 172928 76198 173020 76200
rect 167269 76195 167335 76198
rect 167545 76195 167611 76198
rect 172973 76196 173020 76198
rect 173084 76196 173090 76260
rect 172973 76195 173039 76196
rect 128486 76060 128492 76124
rect 128556 76122 128562 76124
rect 128813 76122 128879 76125
rect 128556 76120 128879 76122
rect 128556 76064 128818 76120
rect 128874 76064 128879 76120
rect 128556 76062 128879 76064
rect 128556 76060 128562 76062
rect 128813 76059 128879 76062
rect 152590 76060 152596 76124
rect 152660 76122 152666 76124
rect 152825 76122 152891 76125
rect 152660 76120 152891 76122
rect 152660 76064 152830 76120
rect 152886 76064 152891 76120
rect 152660 76062 152891 76064
rect 152660 76060 152666 76062
rect 152825 76059 152891 76062
rect 157926 76060 157932 76124
rect 157996 76122 158002 76124
rect 158345 76122 158411 76125
rect 157996 76120 158411 76122
rect 157996 76064 158350 76120
rect 158406 76064 158411 76120
rect 157996 76062 158411 76064
rect 157996 76060 158002 76062
rect 158345 76059 158411 76062
rect 161749 76122 161815 76125
rect 166717 76122 166783 76125
rect 161749 76120 166783 76122
rect 161749 76064 161754 76120
rect 161810 76064 166722 76120
rect 166778 76064 166783 76120
rect 161749 76062 166783 76064
rect 161749 76059 161815 76062
rect 166717 76059 166783 76062
rect 172462 76060 172468 76124
rect 172532 76122 172538 76124
rect 176193 76122 176259 76125
rect 172532 76120 176259 76122
rect 172532 76064 176198 76120
rect 176254 76064 176259 76120
rect 172532 76062 176259 76064
rect 172532 76060 172538 76062
rect 176193 76059 176259 76062
rect 152406 75924 152412 75988
rect 152476 75986 152482 75988
rect 152825 75986 152891 75989
rect 152476 75984 152891 75986
rect 152476 75928 152830 75984
rect 152886 75928 152891 75984
rect 152476 75926 152891 75928
rect 152476 75924 152482 75926
rect 152825 75923 152891 75926
rect 160686 75924 160692 75988
rect 160756 75986 160762 75988
rect 161381 75986 161447 75989
rect 160756 75984 161447 75986
rect 160756 75928 161386 75984
rect 161442 75928 161447 75984
rect 160756 75926 161447 75928
rect 160756 75924 160762 75926
rect 161381 75923 161447 75926
rect 163078 75924 163084 75988
rect 163148 75986 163154 75988
rect 163405 75986 163471 75989
rect 163148 75984 163471 75986
rect 163148 75928 163410 75984
rect 163466 75928 163471 75984
rect 163148 75926 163471 75928
rect 163148 75924 163154 75926
rect 163405 75923 163471 75926
rect 128537 75850 128603 75853
rect 128854 75850 128860 75852
rect 128537 75848 128860 75850
rect 128537 75792 128542 75848
rect 128598 75792 128860 75848
rect 128537 75790 128860 75792
rect 128537 75787 128603 75790
rect 128854 75788 128860 75790
rect 128924 75788 128930 75852
rect 151169 75850 151235 75853
rect 151126 75848 151235 75850
rect 151126 75792 151174 75848
rect 151230 75792 151235 75848
rect 151126 75787 151235 75792
rect 152273 75848 152339 75853
rect 152273 75792 152278 75848
rect 152334 75792 152339 75848
rect 152273 75787 152339 75792
rect 153878 75788 153884 75852
rect 153948 75850 153954 75852
rect 154205 75850 154271 75853
rect 154849 75850 154915 75853
rect 153948 75848 154271 75850
rect 153948 75792 154210 75848
rect 154266 75792 154271 75848
rect 153948 75790 154271 75792
rect 153948 75788 153954 75790
rect 154205 75787 154271 75790
rect 154806 75848 154915 75850
rect 154806 75792 154854 75848
rect 154910 75792 154915 75848
rect 154806 75787 154915 75792
rect 156045 75850 156111 75853
rect 166901 75850 166967 75853
rect 156045 75848 166967 75850
rect 156045 75792 156050 75848
rect 156106 75792 166906 75848
rect 166962 75792 166967 75848
rect 156045 75790 166967 75792
rect 156045 75787 156111 75790
rect 166901 75787 166967 75790
rect 167862 75788 167868 75852
rect 167932 75850 167938 75852
rect 168189 75850 168255 75853
rect 167932 75848 168255 75850
rect 167932 75792 168194 75848
rect 168250 75792 168255 75848
rect 167932 75790 168255 75792
rect 167932 75788 167938 75790
rect 168189 75787 168255 75790
rect 130561 75714 130627 75717
rect 148869 75716 148935 75717
rect 130694 75714 130700 75716
rect 130561 75712 130700 75714
rect 130561 75656 130566 75712
rect 130622 75656 130700 75712
rect 130561 75654 130700 75656
rect 130561 75651 130627 75654
rect 130694 75652 130700 75654
rect 130764 75652 130770 75716
rect 148869 75712 148916 75716
rect 148980 75714 148986 75716
rect 148869 75656 148874 75712
rect 148869 75652 148916 75656
rect 148980 75654 149026 75714
rect 148980 75652 148986 75654
rect 149646 75652 149652 75716
rect 149716 75714 149722 75716
rect 149973 75714 150039 75717
rect 149716 75712 150039 75714
rect 149716 75656 149978 75712
rect 150034 75656 150039 75712
rect 149716 75654 150039 75656
rect 149716 75652 149722 75654
rect 148869 75651 148935 75652
rect 149973 75651 150039 75654
rect 128721 75580 128787 75581
rect 128670 75578 128676 75580
rect 128630 75518 128676 75578
rect 128740 75576 128787 75580
rect 128782 75520 128787 75576
rect 128670 75516 128676 75518
rect 128740 75516 128787 75520
rect 151126 75578 151186 75787
rect 151302 75652 151308 75716
rect 151372 75714 151378 75716
rect 151537 75714 151603 75717
rect 151372 75712 151603 75714
rect 151372 75656 151542 75712
rect 151598 75656 151603 75712
rect 151372 75654 151603 75656
rect 151372 75652 151378 75654
rect 151537 75651 151603 75654
rect 152276 75581 152336 75787
rect 152406 75652 152412 75716
rect 152476 75714 152482 75716
rect 152917 75714 152983 75717
rect 154297 75716 154363 75717
rect 154246 75714 154252 75716
rect 152476 75712 152983 75714
rect 152476 75656 152922 75712
rect 152978 75656 152983 75712
rect 152476 75654 152983 75656
rect 154206 75654 154252 75714
rect 154316 75712 154363 75716
rect 154358 75656 154363 75712
rect 152476 75652 152482 75654
rect 152917 75651 152983 75654
rect 154246 75652 154252 75654
rect 154316 75652 154363 75656
rect 154297 75651 154363 75652
rect 154806 75581 154866 75787
rect 156045 75714 156111 75717
rect 156270 75714 156276 75716
rect 156045 75712 156276 75714
rect 156045 75656 156050 75712
rect 156106 75656 156276 75712
rect 156045 75654 156276 75656
rect 156045 75651 156111 75654
rect 156270 75652 156276 75654
rect 156340 75652 156346 75716
rect 157006 75652 157012 75716
rect 157076 75714 157082 75716
rect 157425 75714 157491 75717
rect 157076 75712 157491 75714
rect 157076 75656 157430 75712
rect 157486 75656 157491 75712
rect 157076 75654 157491 75656
rect 157076 75652 157082 75654
rect 157425 75651 157491 75654
rect 158662 75652 158668 75716
rect 158732 75714 158738 75716
rect 158732 75654 169034 75714
rect 158732 75652 158738 75654
rect 151537 75578 151603 75581
rect 151126 75576 151603 75578
rect 151126 75520 151542 75576
rect 151598 75520 151603 75576
rect 151126 75518 151603 75520
rect 128721 75515 128787 75516
rect 151537 75515 151603 75518
rect 152273 75576 152339 75581
rect 152273 75520 152278 75576
rect 152334 75520 152339 75576
rect 152273 75515 152339 75520
rect 154062 75516 154068 75580
rect 154132 75578 154138 75580
rect 154481 75578 154547 75581
rect 154132 75576 154547 75578
rect 154132 75520 154486 75576
rect 154542 75520 154547 75576
rect 154132 75518 154547 75520
rect 154132 75516 154138 75518
rect 154481 75515 154547 75518
rect 154757 75576 154866 75581
rect 154757 75520 154762 75576
rect 154818 75520 154866 75576
rect 154757 75518 154866 75520
rect 160737 75578 160803 75581
rect 160870 75578 160876 75580
rect 160737 75576 160876 75578
rect 160737 75520 160742 75576
rect 160798 75520 160876 75576
rect 160737 75518 160876 75520
rect 154757 75515 154823 75518
rect 160737 75515 160803 75518
rect 160870 75516 160876 75518
rect 160940 75516 160946 75580
rect 161054 75516 161060 75580
rect 161124 75578 161130 75580
rect 161289 75578 161355 75581
rect 161124 75576 161355 75578
rect 161124 75520 161294 75576
rect 161350 75520 161355 75576
rect 161124 75518 161355 75520
rect 161124 75516 161130 75518
rect 161289 75515 161355 75518
rect 163262 75516 163268 75580
rect 163332 75578 163338 75580
rect 163589 75578 163655 75581
rect 163332 75576 163655 75578
rect 163332 75520 163594 75576
rect 163650 75520 163655 75576
rect 163332 75518 163655 75520
rect 168974 75578 169034 75654
rect 170070 75652 170076 75716
rect 170140 75714 170146 75716
rect 170305 75714 170371 75717
rect 170140 75712 170371 75714
rect 170140 75656 170310 75712
rect 170366 75656 170371 75712
rect 170140 75654 170371 75656
rect 170140 75652 170146 75654
rect 170305 75651 170371 75654
rect 170581 75714 170647 75717
rect 170990 75714 170996 75716
rect 170581 75712 170996 75714
rect 170581 75656 170586 75712
rect 170642 75656 170996 75712
rect 170581 75654 170996 75656
rect 170581 75651 170647 75654
rect 170990 75652 170996 75654
rect 171060 75652 171066 75716
rect 174537 75578 174603 75581
rect 168974 75576 174603 75578
rect 168974 75520 174542 75576
rect 174598 75520 174603 75576
rect 168974 75518 174603 75520
rect 163332 75516 163338 75518
rect 163589 75515 163655 75518
rect 174537 75515 174603 75518
rect 126605 75442 126671 75445
rect 130510 75442 130516 75444
rect 126605 75440 130516 75442
rect 126605 75384 126610 75440
rect 126666 75384 130516 75440
rect 126605 75382 130516 75384
rect 126605 75379 126671 75382
rect 130510 75380 130516 75382
rect 130580 75380 130586 75444
rect 157057 75442 157123 75445
rect 172329 75442 172395 75445
rect 157057 75440 172395 75442
rect 157057 75384 157062 75440
rect 157118 75384 172334 75440
rect 172390 75384 172395 75440
rect 157057 75382 172395 75384
rect 157057 75379 157123 75382
rect 172329 75379 172395 75382
rect 153285 75308 153351 75309
rect 164509 75308 164575 75309
rect 153285 75306 153332 75308
rect 153240 75304 153332 75306
rect 153240 75248 153290 75304
rect 153240 75246 153332 75248
rect 153285 75244 153332 75246
rect 153396 75244 153402 75308
rect 164509 75306 164556 75308
rect 164464 75304 164556 75306
rect 164464 75248 164514 75304
rect 164464 75246 164556 75248
rect 164509 75244 164556 75246
rect 164620 75244 164626 75308
rect 153285 75243 153351 75244
rect 164509 75243 164575 75244
rect 125317 75170 125383 75173
rect 125910 75170 125916 75172
rect 125317 75168 125916 75170
rect 125317 75112 125322 75168
rect 125378 75112 125916 75168
rect 125317 75110 125916 75112
rect 125317 75107 125383 75110
rect 125910 75108 125916 75110
rect 125980 75108 125986 75172
rect 144126 75108 144132 75172
rect 144196 75170 144202 75172
rect 144913 75170 144979 75173
rect 144196 75168 144979 75170
rect 144196 75112 144918 75168
rect 144974 75112 144979 75168
rect 144196 75110 144979 75112
rect 144196 75108 144202 75110
rect 144913 75107 144979 75110
rect 158897 75170 158963 75173
rect 159030 75170 159036 75172
rect 158897 75168 159036 75170
rect 158897 75112 158902 75168
rect 158958 75112 159036 75168
rect 158897 75110 159036 75112
rect 158897 75107 158963 75110
rect 159030 75108 159036 75110
rect 159100 75108 159106 75172
rect 164734 75108 164740 75172
rect 164804 75170 164810 75172
rect 164969 75170 165035 75173
rect 164804 75168 165035 75170
rect 164804 75112 164974 75168
rect 165030 75112 165035 75168
rect 164804 75110 165035 75112
rect 164804 75108 164810 75110
rect 164969 75107 165035 75110
rect 166073 75170 166139 75173
rect 518893 75170 518959 75173
rect 166073 75168 518959 75170
rect 166073 75112 166078 75168
rect 166134 75112 518898 75168
rect 518954 75112 518959 75168
rect 166073 75110 518959 75112
rect 166073 75107 166139 75110
rect 518893 75107 518959 75110
rect 132677 75034 132743 75037
rect 134057 75036 134123 75037
rect 133086 75034 133092 75036
rect 132677 75032 133092 75034
rect 132677 74976 132682 75032
rect 132738 74976 133092 75032
rect 132677 74974 133092 74976
rect 132677 74971 132743 74974
rect 133086 74972 133092 74974
rect 133156 74972 133162 75036
rect 134006 75034 134012 75036
rect 133966 74974 134012 75034
rect 134076 75032 134123 75036
rect 134118 74976 134123 75032
rect 134006 74972 134012 74974
rect 134076 74972 134123 74976
rect 134057 74971 134123 74972
rect 135437 75034 135503 75037
rect 136081 75036 136147 75037
rect 137921 75036 137987 75037
rect 135662 75034 135668 75036
rect 135437 75032 135668 75034
rect 135437 74976 135442 75032
rect 135498 74976 135668 75032
rect 135437 74974 135668 74976
rect 135437 74971 135503 74974
rect 135662 74972 135668 74974
rect 135732 74972 135738 75036
rect 136030 74972 136036 75036
rect 136100 75034 136147 75036
rect 137870 75034 137876 75036
rect 136100 75032 136192 75034
rect 136142 74976 136192 75032
rect 136100 74974 136192 74976
rect 137830 74974 137876 75034
rect 137940 75032 137987 75036
rect 137982 74976 137987 75032
rect 136100 74972 136147 74974
rect 137870 74972 137876 74974
rect 137940 74972 137987 74976
rect 138790 74972 138796 75036
rect 138860 75034 138866 75036
rect 138933 75034 138999 75037
rect 138860 75032 138999 75034
rect 138860 74976 138938 75032
rect 138994 74976 138999 75032
rect 138860 74974 138999 74976
rect 138860 74972 138866 74974
rect 136081 74971 136147 74972
rect 137921 74971 137987 74972
rect 138933 74971 138999 74974
rect 139853 75034 139919 75037
rect 140078 75034 140084 75036
rect 139853 75032 140084 75034
rect 139853 74976 139858 75032
rect 139914 74976 140084 75032
rect 139853 74974 140084 74976
rect 139853 74971 139919 74974
rect 140078 74972 140084 74974
rect 140148 74972 140154 75036
rect 140446 74972 140452 75036
rect 140516 75034 140522 75036
rect 140589 75034 140655 75037
rect 140516 75032 140655 75034
rect 140516 74976 140594 75032
rect 140650 74976 140655 75032
rect 140516 74974 140655 74976
rect 140516 74972 140522 74974
rect 140589 74971 140655 74974
rect 144494 74972 144500 75036
rect 144564 75034 144570 75036
rect 144637 75034 144703 75037
rect 144564 75032 144703 75034
rect 144564 74976 144642 75032
rect 144698 74976 144703 75032
rect 144564 74974 144703 74976
rect 144564 74972 144570 74974
rect 144637 74971 144703 74974
rect 145097 75034 145163 75037
rect 148777 75036 148843 75037
rect 145230 75034 145236 75036
rect 145097 75032 145236 75034
rect 145097 74976 145102 75032
rect 145158 74976 145236 75032
rect 145097 74974 145236 74976
rect 145097 74971 145163 74974
rect 145230 74972 145236 74974
rect 145300 74972 145306 75036
rect 148726 75034 148732 75036
rect 148686 74974 148732 75034
rect 148796 75032 148843 75036
rect 148838 74976 148843 75032
rect 148726 74972 148732 74974
rect 148796 74972 148843 74976
rect 152038 74972 152044 75036
rect 152108 75034 152114 75036
rect 154021 75034 154087 75037
rect 152108 75032 154087 75034
rect 152108 74976 154026 75032
rect 154082 74976 154087 75032
rect 152108 74974 154087 74976
rect 152108 74972 152114 74974
rect 148777 74971 148843 74972
rect 154021 74971 154087 74974
rect 158846 74972 158852 75036
rect 158916 75034 158922 75036
rect 160001 75034 160067 75037
rect 170213 75036 170279 75037
rect 170213 75034 170260 75036
rect 158916 75032 160067 75034
rect 158916 74976 160006 75032
rect 160062 74976 160067 75032
rect 158916 74974 160067 74976
rect 170168 75032 170260 75034
rect 170168 74976 170218 75032
rect 170168 74974 170260 74976
rect 158916 74972 158922 74974
rect 160001 74971 160067 74974
rect 170213 74972 170260 74974
rect 170324 74972 170330 75036
rect 170213 74971 170279 74972
rect 131113 74898 131179 74901
rect 131430 74898 131436 74900
rect 131113 74896 131436 74898
rect 131113 74840 131118 74896
rect 131174 74840 131436 74896
rect 131113 74838 131436 74840
rect 131113 74835 131179 74838
rect 131430 74836 131436 74838
rect 131500 74836 131506 74900
rect 140262 74836 140268 74900
rect 140332 74898 140338 74900
rect 140681 74898 140747 74901
rect 140332 74896 140747 74898
rect 140332 74840 140686 74896
rect 140742 74840 140747 74896
rect 140332 74838 140747 74840
rect 140332 74836 140338 74838
rect 140681 74835 140747 74838
rect 142838 74836 142844 74900
rect 142908 74898 142914 74900
rect 143257 74898 143323 74901
rect 142908 74896 143323 74898
rect 142908 74840 143262 74896
rect 143318 74840 143323 74896
rect 142908 74838 143323 74840
rect 142908 74836 142914 74838
rect 143257 74835 143323 74838
rect 131062 74700 131068 74764
rect 131132 74762 131138 74764
rect 131205 74762 131271 74765
rect 131132 74760 131271 74762
rect 131132 74704 131210 74760
rect 131266 74704 131271 74760
rect 131132 74702 131271 74704
rect 131132 74700 131138 74702
rect 131205 74699 131271 74702
rect 143022 74700 143028 74764
rect 143092 74762 143098 74764
rect 143165 74762 143231 74765
rect 143441 74764 143507 74765
rect 143390 74762 143396 74764
rect 143092 74760 143231 74762
rect 143092 74704 143170 74760
rect 143226 74704 143231 74760
rect 143092 74702 143231 74704
rect 143350 74702 143396 74762
rect 143460 74760 143507 74764
rect 143502 74704 143507 74760
rect 143092 74700 143098 74702
rect 143165 74699 143231 74702
rect 143390 74700 143396 74702
rect 143460 74700 143507 74704
rect 167310 74700 167316 74764
rect 167380 74762 167386 74764
rect 167821 74762 167887 74765
rect 170765 74762 170831 74765
rect 171726 74762 171732 74764
rect 167380 74760 167887 74762
rect 167380 74704 167826 74760
rect 167882 74704 167887 74760
rect 167380 74702 167887 74704
rect 167380 74700 167386 74702
rect 143441 74699 143507 74700
rect 167821 74699 167887 74702
rect 169158 74702 169954 74762
rect 131297 74628 131363 74629
rect 131246 74626 131252 74628
rect 131206 74566 131252 74626
rect 131316 74624 131363 74628
rect 131358 74568 131363 74624
rect 131246 74564 131252 74566
rect 131316 74564 131363 74568
rect 140998 74564 141004 74628
rect 141068 74626 141074 74628
rect 142061 74626 142127 74629
rect 141068 74624 142127 74626
rect 141068 74568 142066 74624
rect 142122 74568 142127 74624
rect 141068 74566 142127 74568
rect 141068 74564 141074 74566
rect 131297 74563 131363 74564
rect 142061 74563 142127 74566
rect 143206 74564 143212 74628
rect 143276 74626 143282 74628
rect 143349 74626 143415 74629
rect 143276 74624 143415 74626
rect 143276 74568 143354 74624
rect 143410 74568 143415 74624
rect 143276 74566 143415 74568
rect 143276 74564 143282 74566
rect 143349 74563 143415 74566
rect 148542 74564 148548 74628
rect 148612 74626 148618 74628
rect 148961 74626 149027 74629
rect 148612 74624 149027 74626
rect 148612 74568 148966 74624
rect 149022 74568 149027 74624
rect 148612 74566 149027 74568
rect 148612 74564 148618 74566
rect 148961 74563 149027 74566
rect 159633 74626 159699 74629
rect 169158 74626 169218 74702
rect 159633 74624 169218 74626
rect 159633 74568 159638 74624
rect 159694 74568 169218 74624
rect 159633 74566 169218 74568
rect 169894 74626 169954 74702
rect 170765 74760 171732 74762
rect 170765 74704 170770 74760
rect 170826 74704 171732 74760
rect 170765 74702 171732 74704
rect 170765 74699 170831 74702
rect 171726 74700 171732 74702
rect 171796 74700 171802 74764
rect 175641 74762 175707 74765
rect 504357 74762 504423 74765
rect 175641 74760 504423 74762
rect 175641 74704 175646 74760
rect 175702 74704 504362 74760
rect 504418 74704 504423 74760
rect 175641 74702 504423 74704
rect 175641 74699 175707 74702
rect 504357 74699 504423 74702
rect 171685 74626 171751 74629
rect 169894 74566 170506 74626
rect 159633 74563 159699 74566
rect 132769 74490 132835 74493
rect 160461 74492 160527 74493
rect 133270 74490 133276 74492
rect 132769 74488 133276 74490
rect 132769 74432 132774 74488
rect 132830 74432 133276 74488
rect 132769 74430 133276 74432
rect 132769 74427 132835 74430
rect 133270 74428 133276 74430
rect 133340 74428 133346 74492
rect 160461 74490 160508 74492
rect 160416 74488 160508 74490
rect 160416 74432 160466 74488
rect 160416 74430 160508 74432
rect 160461 74428 160508 74430
rect 160572 74428 160578 74492
rect 170446 74490 170506 74566
rect 170814 74624 171751 74626
rect 170814 74568 171690 74624
rect 171746 74568 171751 74624
rect 170814 74566 171751 74568
rect 170814 74490 170874 74566
rect 171685 74563 171751 74566
rect 170446 74430 170874 74490
rect 160461 74427 160527 74428
rect 134149 74354 134215 74357
rect 118650 74352 134215 74354
rect 118650 74296 134154 74352
rect 134210 74296 134215 74352
rect 118650 74294 134215 74296
rect 111793 74082 111859 74085
rect 118650 74082 118710 74294
rect 134149 74291 134215 74294
rect 166993 74354 167059 74357
rect 169385 74354 169451 74357
rect 166993 74352 169451 74354
rect 166993 74296 166998 74352
rect 167054 74296 169390 74352
rect 169446 74296 169451 74352
rect 166993 74294 169451 74296
rect 166993 74291 167059 74294
rect 169385 74291 169451 74294
rect 128629 74218 128695 74221
rect 132585 74218 132651 74221
rect 128629 74216 132651 74218
rect 128629 74160 128634 74216
rect 128690 74160 132590 74216
rect 132646 74160 132651 74216
rect 128629 74158 132651 74160
rect 128629 74155 128695 74158
rect 132585 74155 132651 74158
rect 141969 74218 142035 74221
rect 166993 74218 167059 74221
rect 141969 74216 167059 74218
rect 141969 74160 141974 74216
rect 142030 74160 166998 74216
rect 167054 74160 167059 74216
rect 141969 74158 167059 74160
rect 141969 74155 142035 74158
rect 166993 74155 167059 74158
rect 111793 74080 118710 74082
rect 111793 74024 111798 74080
rect 111854 74024 118710 74080
rect 111793 74022 118710 74024
rect 144729 74082 144795 74085
rect 247033 74082 247099 74085
rect 144729 74080 247099 74082
rect 144729 74024 144734 74080
rect 144790 74024 247038 74080
rect 247094 74024 247099 74080
rect 144729 74022 247099 74024
rect 111793 74019 111859 74022
rect 144729 74019 144795 74022
rect 247033 74019 247099 74022
rect 20713 73946 20779 73949
rect 121361 73946 121427 73949
rect 20713 73944 121427 73946
rect 20713 73888 20718 73944
rect 20774 73888 121366 73944
rect 121422 73888 121427 73944
rect 20713 73886 121427 73888
rect 20713 73883 20779 73886
rect 121361 73883 121427 73886
rect 138289 73946 138355 73949
rect 138606 73946 138612 73948
rect 138289 73944 138612 73946
rect 138289 73888 138294 73944
rect 138350 73888 138612 73944
rect 138289 73886 138612 73888
rect 138289 73883 138355 73886
rect 138606 73884 138612 73886
rect 138676 73884 138682 73948
rect 147581 73946 147647 73949
rect 282913 73946 282979 73949
rect 147581 73944 282979 73946
rect 147581 73888 147586 73944
rect 147642 73888 282918 73944
rect 282974 73888 282979 73944
rect 147581 73886 282979 73888
rect 147581 73883 147647 73886
rect 282913 73883 282979 73886
rect 1393 73810 1459 73813
rect 125501 73810 125567 73813
rect 1393 73808 125567 73810
rect 1393 73752 1398 73808
rect 1454 73752 125506 73808
rect 125562 73752 125567 73808
rect 1393 73750 125567 73752
rect 1393 73747 1459 73750
rect 125501 73747 125567 73750
rect 136398 73748 136404 73812
rect 136468 73810 136474 73812
rect 138013 73810 138079 73813
rect 136468 73808 138079 73810
rect 136468 73752 138018 73808
rect 138074 73752 138079 73808
rect 136468 73750 138079 73752
rect 136468 73748 136474 73750
rect 138013 73747 138079 73750
rect 166993 73810 167059 73813
rect 171961 73810 172027 73813
rect 565813 73810 565879 73813
rect 166993 73808 172027 73810
rect 166993 73752 166998 73808
rect 167054 73752 171966 73808
rect 172022 73752 172027 73808
rect 166993 73750 172027 73752
rect 166993 73747 167059 73750
rect 171961 73747 172027 73750
rect 176610 73808 565879 73810
rect 176610 73752 565818 73808
rect 565874 73752 565879 73808
rect 176610 73750 565879 73752
rect 169569 73674 169635 73677
rect 176610 73674 176670 73750
rect 565813 73747 565879 73750
rect 169569 73672 176670 73674
rect 169569 73616 169574 73672
rect 169630 73616 176670 73672
rect 169569 73614 176670 73616
rect 169569 73611 169635 73614
rect 147070 73476 147076 73540
rect 147140 73538 147146 73540
rect 147397 73538 147463 73541
rect 147140 73536 147463 73538
rect 147140 73480 147402 73536
rect 147458 73480 147463 73536
rect 147140 73478 147463 73480
rect 147140 73476 147146 73478
rect 147397 73475 147463 73478
rect 165705 73538 165771 73541
rect 166022 73538 166028 73540
rect 165705 73536 166028 73538
rect 165705 73480 165710 73536
rect 165766 73480 166028 73536
rect 165705 73478 166028 73480
rect 165705 73475 165771 73478
rect 166022 73476 166028 73478
rect 166092 73476 166098 73540
rect 136582 73340 136588 73404
rect 136652 73402 136658 73404
rect 137277 73402 137343 73405
rect 136652 73400 137343 73402
rect 136652 73344 137282 73400
rect 137338 73344 137343 73400
rect 136652 73342 137343 73344
rect 136652 73340 136658 73342
rect 137277 73339 137343 73342
rect 170857 73266 170923 73269
rect 171910 73266 171916 73268
rect 170857 73264 171916 73266
rect 170857 73208 170862 73264
rect 170918 73208 171916 73264
rect 170857 73206 171916 73208
rect 170857 73203 170923 73206
rect 171910 73204 171916 73206
rect 171980 73204 171986 73268
rect 160318 73068 160324 73132
rect 160388 73130 160394 73132
rect 163865 73130 163931 73133
rect 160388 73128 163931 73130
rect 160388 73072 163870 73128
rect 163926 73072 163931 73128
rect 160388 73070 163931 73072
rect 160388 73068 160394 73070
rect 163865 73067 163931 73070
rect 139117 72994 139183 72997
rect 173893 72994 173959 72997
rect 139117 72992 173959 72994
rect 139117 72936 139122 72992
rect 139178 72936 173898 72992
rect 173954 72936 173959 72992
rect 139117 72934 173959 72936
rect 139117 72931 139183 72934
rect 173893 72931 173959 72934
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 151721 72860 151787 72861
rect 151670 72858 151676 72860
rect 151630 72798 151676 72858
rect 151740 72856 151787 72860
rect 151782 72800 151787 72856
rect 151670 72796 151676 72798
rect 151740 72796 151787 72800
rect 151721 72795 151787 72796
rect 155769 72858 155835 72861
rect 389173 72858 389239 72861
rect 155769 72856 389239 72858
rect 155769 72800 155774 72856
rect 155830 72800 389178 72856
rect 389234 72800 389239 72856
rect 583520 72844 584960 72934
rect 155769 72798 389239 72800
rect 155769 72795 155835 72798
rect 389173 72795 389239 72798
rect 57973 72722 58039 72725
rect 129825 72722 129891 72725
rect 57973 72720 129891 72722
rect 57973 72664 57978 72720
rect 58034 72664 129830 72720
rect 129886 72664 129891 72720
rect 57973 72662 129891 72664
rect 57973 72659 58039 72662
rect 129825 72659 129891 72662
rect 157149 72722 157215 72725
rect 402973 72722 403039 72725
rect 157149 72720 403039 72722
rect 157149 72664 157154 72720
rect 157210 72664 402978 72720
rect 403034 72664 403039 72720
rect 157149 72662 403039 72664
rect 157149 72659 157215 72662
rect 402973 72659 403039 72662
rect 53833 72586 53899 72589
rect 129774 72586 129780 72588
rect 53833 72584 129780 72586
rect 53833 72528 53838 72584
rect 53894 72528 129780 72584
rect 53833 72526 129780 72528
rect 53833 72523 53899 72526
rect 129774 72524 129780 72526
rect 129844 72524 129850 72588
rect 165337 72586 165403 72589
rect 496813 72586 496879 72589
rect 165337 72584 496879 72586
rect 165337 72528 165342 72584
rect 165398 72528 496818 72584
rect 496874 72528 496879 72584
rect 165337 72526 496879 72528
rect 165337 72523 165403 72526
rect 496813 72523 496879 72526
rect 2773 72450 2839 72453
rect 125685 72450 125751 72453
rect 2773 72448 125751 72450
rect 2773 72392 2778 72448
rect 2834 72392 125690 72448
rect 125746 72392 125751 72448
rect 2773 72390 125751 72392
rect 2773 72387 2839 72390
rect 125685 72387 125751 72390
rect 170489 72450 170555 72453
rect 514753 72450 514819 72453
rect 170489 72448 514819 72450
rect 170489 72392 170494 72448
rect 170550 72392 514758 72448
rect 514814 72392 514819 72448
rect 170489 72390 514819 72392
rect 170489 72387 170555 72390
rect 514753 72387 514819 72390
rect 126237 71906 126303 71909
rect 131430 71906 131436 71908
rect 126237 71904 131436 71906
rect 126237 71848 126242 71904
rect 126298 71848 131436 71904
rect 126237 71846 131436 71848
rect 126237 71843 126303 71846
rect 131430 71844 131436 71846
rect 131500 71844 131506 71908
rect 130377 71770 130443 71773
rect 135294 71770 135300 71772
rect 130377 71768 135300 71770
rect -960 71634 480 71724
rect 130377 71712 130382 71768
rect 130438 71712 135300 71768
rect 130377 71710 135300 71712
rect 130377 71707 130443 71710
rect 135294 71708 135300 71710
rect 135364 71708 135370 71772
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 143390 71436 143396 71500
rect 143460 71498 143466 71500
rect 230473 71498 230539 71501
rect 143460 71496 230539 71498
rect 143460 71440 230478 71496
rect 230534 71440 230539 71496
rect 143460 71438 230539 71440
rect 143460 71436 143466 71438
rect 230473 71435 230539 71438
rect 126605 71364 126671 71365
rect 126605 71362 126652 71364
rect 126560 71360 126652 71362
rect 126560 71304 126610 71360
rect 126560 71302 126652 71304
rect 126605 71300 126652 71302
rect 126716 71300 126722 71364
rect 144862 71300 144868 71364
rect 144932 71362 144938 71364
rect 244273 71362 244339 71365
rect 144932 71360 244339 71362
rect 144932 71304 244278 71360
rect 244334 71304 244339 71360
rect 144932 71302 244339 71304
rect 144932 71300 144938 71302
rect 126605 71299 126671 71300
rect 244273 71299 244339 71302
rect 89713 71226 89779 71229
rect 132493 71226 132559 71229
rect 89713 71224 132559 71226
rect 89713 71168 89718 71224
rect 89774 71168 132498 71224
rect 132554 71168 132559 71224
rect 89713 71166 132559 71168
rect 89713 71163 89779 71166
rect 132493 71163 132559 71166
rect 146201 71226 146267 71229
rect 266353 71226 266419 71229
rect 146201 71224 266419 71226
rect 146201 71168 146206 71224
rect 146262 71168 266358 71224
rect 266414 71168 266419 71224
rect 146201 71166 266419 71168
rect 146201 71163 146267 71166
rect 266353 71163 266419 71166
rect 35893 71090 35959 71093
rect 129038 71090 129044 71092
rect 35893 71088 129044 71090
rect 35893 71032 35898 71088
rect 35954 71032 129044 71088
rect 35893 71030 129044 71032
rect 35893 71027 35959 71030
rect 129038 71028 129044 71030
rect 129108 71028 129114 71092
rect 170990 71028 170996 71092
rect 171060 71090 171066 71092
rect 578233 71090 578299 71093
rect 171060 71088 578299 71090
rect 171060 71032 578238 71088
rect 578294 71032 578299 71088
rect 171060 71030 578299 71032
rect 171060 71028 171066 71030
rect 578233 71027 578299 71030
rect 165838 70892 165844 70956
rect 165908 70954 165914 70956
rect 166073 70954 166139 70957
rect 165908 70952 166139 70954
rect 165908 70896 166078 70952
rect 166134 70896 166139 70952
rect 165908 70894 166139 70896
rect 165908 70892 165914 70894
rect 166073 70891 166139 70894
rect 164926 70486 173266 70546
rect 164926 70412 164986 70486
rect 173206 70413 173266 70486
rect 164918 70348 164924 70412
rect 164988 70348 164994 70412
rect 173206 70408 173315 70413
rect 173206 70352 173254 70408
rect 173310 70352 173315 70408
rect 173206 70350 173315 70352
rect 173249 70347 173315 70350
rect 162710 69940 162716 70004
rect 162780 70002 162786 70004
rect 172145 70002 172211 70005
rect 162780 70000 172211 70002
rect 162780 69944 172150 70000
rect 172206 69944 172211 70000
rect 162780 69942 172211 69944
rect 162780 69940 162786 69942
rect 172145 69939 172211 69942
rect 150157 69866 150223 69869
rect 284385 69866 284451 69869
rect 150157 69864 284451 69866
rect 150157 69808 150162 69864
rect 150218 69808 284390 69864
rect 284446 69808 284451 69864
rect 150157 69806 284451 69808
rect 150157 69803 150223 69806
rect 284385 69803 284451 69806
rect 149053 69730 149119 69733
rect 298093 69730 298159 69733
rect 149053 69728 298159 69730
rect 149053 69672 149058 69728
rect 149114 69672 298098 69728
rect 298154 69672 298159 69728
rect 149053 69670 298159 69672
rect 149053 69667 149119 69670
rect 298093 69667 298159 69670
rect 150341 69594 150407 69597
rect 318793 69594 318859 69597
rect 150341 69592 318859 69594
rect 150341 69536 150346 69592
rect 150402 69536 318798 69592
rect 318854 69536 318859 69592
rect 150341 69534 318859 69536
rect 150341 69531 150407 69534
rect 318793 69531 318859 69534
rect 154430 68172 154436 68236
rect 154500 68234 154506 68236
rect 367093 68234 367159 68237
rect 154500 68232 367159 68234
rect 154500 68176 367098 68232
rect 367154 68176 367159 68232
rect 154500 68174 367159 68176
rect 154500 68172 154506 68174
rect 367093 68171 367159 68174
rect 152958 66812 152964 66876
rect 153028 66874 153034 66876
rect 353293 66874 353359 66877
rect 153028 66872 353359 66874
rect 153028 66816 353298 66872
rect 353354 66816 353359 66872
rect 153028 66814 353359 66816
rect 153028 66812 153034 66814
rect 353293 66811 353359 66814
rect 138790 65452 138796 65516
rect 138860 65514 138866 65516
rect 172513 65514 172579 65517
rect 138860 65512 172579 65514
rect 138860 65456 172518 65512
rect 172574 65456 172579 65512
rect 138860 65454 172579 65456
rect 138860 65452 138866 65454
rect 172513 65451 172579 65454
rect 138974 63004 138980 63068
rect 139044 63066 139050 63068
rect 175273 63066 175339 63069
rect 139044 63064 175339 63066
rect 139044 63008 175278 63064
rect 175334 63008 175339 63064
rect 139044 63006 175339 63008
rect 139044 63004 139050 63006
rect 175273 63003 175339 63006
rect 140078 62868 140084 62932
rect 140148 62930 140154 62932
rect 193213 62930 193279 62933
rect 140148 62928 193279 62930
rect 140148 62872 193218 62928
rect 193274 62872 193279 62928
rect 140148 62870 193279 62872
rect 140148 62868 140154 62870
rect 193213 62867 193279 62870
rect 166206 62732 166212 62796
rect 166276 62794 166282 62796
rect 529933 62794 529999 62797
rect 166276 62792 529999 62794
rect 166276 62736 529938 62792
rect 529994 62736 529999 62792
rect 166276 62734 529999 62736
rect 166276 62732 166282 62734
rect 529933 62731 529999 62734
rect 158846 59876 158852 59940
rect 158916 59938 158922 59940
rect 441613 59938 441679 59941
rect 158916 59936 441679 59938
rect 158916 59880 441618 59936
rect 441674 59880 441679 59936
rect 158916 59878 441679 59880
rect 158916 59876 158922 59878
rect 441613 59875 441679 59878
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3601 58578 3667 58581
rect -960 58576 3667 58578
rect -960 58520 3606 58576
rect 3662 58520 3667 58576
rect -960 58518 3667 58520
rect -960 58428 480 58518
rect 3601 58515 3667 58518
rect 140262 57292 140268 57356
rect 140332 57354 140338 57356
rect 194593 57354 194659 57357
rect 140332 57352 194659 57354
rect 140332 57296 194598 57352
rect 194654 57296 194659 57352
rect 140332 57294 194659 57296
rect 140332 57292 140338 57294
rect 194593 57291 194659 57294
rect 144494 57156 144500 57220
rect 144564 57218 144570 57220
rect 245653 57218 245719 57221
rect 144564 57216 245719 57218
rect 144564 57160 245658 57216
rect 245714 57160 245719 57216
rect 144564 57158 245719 57160
rect 144564 57156 144570 57158
rect 245653 57155 245719 57158
rect 156822 54436 156828 54500
rect 156892 54498 156898 54500
rect 405733 54498 405799 54501
rect 156892 54496 405799 54498
rect 156892 54440 405738 54496
rect 405794 54440 405799 54496
rect 156892 54438 405799 54440
rect 156892 54436 156898 54438
rect 405733 54435 405799 54438
rect 171910 50220 171916 50284
rect 171980 50282 171986 50284
rect 582373 50282 582439 50285
rect 171980 50280 582439 50282
rect 171980 50224 582378 50280
rect 582434 50224 582439 50280
rect 171980 50222 582439 50224
rect 171980 50220 171986 50222
rect 582373 50219 582439 50222
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 162342 39204 162348 39268
rect 162412 39266 162418 39268
rect 476113 39266 476179 39269
rect 162412 39264 476179 39266
rect 162412 39208 476118 39264
rect 476174 39208 476179 39264
rect 162412 39206 476179 39208
rect 162412 39204 162418 39206
rect 476113 39203 476179 39206
rect 157926 36484 157932 36548
rect 157996 36546 158002 36548
rect 422293 36546 422359 36549
rect 157996 36544 422359 36546
rect 157996 36488 422298 36544
rect 422354 36488 422359 36544
rect 157996 36486 422359 36488
rect 157996 36484 158002 36486
rect 422293 36483 422359 36486
rect 147254 35260 147260 35324
rect 147324 35322 147330 35324
rect 280153 35322 280219 35325
rect 147324 35320 280219 35322
rect 147324 35264 280158 35320
rect 280214 35264 280219 35320
rect 147324 35262 280219 35264
rect 147324 35260 147330 35262
rect 280153 35259 280219 35262
rect 149830 35124 149836 35188
rect 149900 35186 149906 35188
rect 316125 35186 316191 35189
rect 149900 35184 316191 35186
rect 149900 35128 316130 35184
rect 316186 35128 316191 35184
rect 149900 35126 316191 35128
rect 149900 35124 149906 35126
rect 316125 35123 316191 35126
rect 139158 33900 139164 33964
rect 139228 33962 139234 33964
rect 176653 33962 176719 33965
rect 139228 33960 176719 33962
rect 139228 33904 176658 33960
rect 176714 33904 176719 33960
rect 139228 33902 176719 33904
rect 139228 33900 139234 33902
rect 176653 33899 176719 33902
rect 143022 33764 143028 33828
rect 143092 33826 143098 33828
rect 226425 33826 226491 33829
rect 143092 33824 226491 33826
rect 143092 33768 226430 33824
rect 226486 33768 226491 33824
rect 143092 33766 226491 33768
rect 143092 33764 143098 33766
rect 226425 33763 226491 33766
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect 166390 32676 166396 32740
rect 166460 32738 166466 32740
rect 528553 32738 528619 32741
rect 166460 32736 528619 32738
rect 166460 32680 528558 32736
rect 528614 32680 528619 32736
rect 166460 32678 528619 32680
rect 166460 32676 166466 32678
rect 528553 32675 528619 32678
rect -960 32466 480 32556
rect 167678 32540 167684 32604
rect 167748 32602 167754 32604
rect 546493 32602 546559 32605
rect 167748 32600 546559 32602
rect 167748 32544 546498 32600
rect 546554 32544 546559 32600
rect 167748 32542 546559 32544
rect 167748 32540 167754 32542
rect 546493 32539 546559 32542
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 167494 32404 167500 32468
rect 167564 32466 167570 32468
rect 549253 32466 549319 32469
rect 167564 32464 549319 32466
rect 167564 32408 549258 32464
rect 549314 32408 549319 32464
rect 167564 32406 549319 32408
rect 167564 32404 167570 32406
rect 549253 32403 549319 32406
rect 160686 30908 160692 30972
rect 160756 30970 160762 30972
rect 460933 30970 460999 30973
rect 160756 30968 460999 30970
rect 160756 30912 460938 30968
rect 460994 30912 460999 30968
rect 160756 30910 460999 30912
rect 160756 30908 160762 30910
rect 460933 30907 460999 30910
rect 162526 29548 162532 29612
rect 162596 29610 162602 29612
rect 473353 29610 473419 29613
rect 162596 29608 473419 29610
rect 162596 29552 473358 29608
rect 473414 29552 473419 29608
rect 162596 29550 473419 29552
rect 162596 29548 162602 29550
rect 473353 29547 473419 29550
rect 143206 28188 143212 28252
rect 143276 28250 143282 28252
rect 229093 28250 229159 28253
rect 143276 28248 229159 28250
rect 143276 28192 229098 28248
rect 229154 28192 229159 28248
rect 143276 28190 229159 28192
rect 143276 28188 143282 28190
rect 229093 28187 229159 28190
rect 140446 26964 140452 27028
rect 140516 27026 140522 27028
rect 193305 27026 193371 27029
rect 140516 27024 193371 27026
rect 140516 26968 193310 27024
rect 193366 26968 193371 27024
rect 140516 26966 193371 26968
rect 140516 26964 140522 26966
rect 193305 26963 193371 26966
rect 169334 26828 169340 26892
rect 169404 26890 169410 26892
rect 567193 26890 567259 26893
rect 169404 26888 567259 26890
rect 169404 26832 567198 26888
rect 567254 26832 567259 26888
rect 169404 26830 567259 26832
rect 169404 26828 169410 26830
rect 567193 26827 567259 26830
rect 149646 25468 149652 25532
rect 149716 25530 149722 25532
rect 317413 25530 317479 25533
rect 149716 25528 317479 25530
rect 149716 25472 317418 25528
rect 317474 25472 317479 25528
rect 149716 25470 317479 25472
rect 149716 25468 149722 25470
rect 317413 25467 317479 25470
rect 167862 24244 167868 24308
rect 167932 24306 167938 24308
rect 547873 24306 547939 24309
rect 167932 24304 547939 24306
rect 167932 24248 547878 24304
rect 547934 24248 547939 24304
rect 167932 24246 547939 24248
rect 167932 24244 167938 24246
rect 547873 24243 547939 24246
rect 170806 24108 170812 24172
rect 170876 24170 170882 24172
rect 576853 24170 576919 24173
rect 170876 24168 576919 24170
rect 170876 24112 576858 24168
rect 576914 24112 576919 24168
rect 170876 24110 576919 24112
rect 170876 24108 170882 24110
rect 576853 24107 576919 24110
rect 166574 22612 166580 22676
rect 166644 22674 166650 22676
rect 531313 22674 531379 22677
rect 166644 22672 531379 22674
rect 166644 22616 531318 22672
rect 531374 22616 531379 22672
rect 166644 22614 531379 22616
rect 166644 22612 166650 22614
rect 531313 22611 531379 22614
rect 159030 21388 159036 21452
rect 159100 21450 159106 21452
rect 442993 21450 443059 21453
rect 159100 21448 443059 21450
rect 159100 21392 442998 21448
rect 443054 21392 443059 21448
rect 159100 21390 443059 21392
rect 159100 21388 159106 21390
rect 442993 21387 443059 21390
rect 165286 21252 165292 21316
rect 165356 21314 165362 21316
rect 513373 21314 513439 21317
rect 165356 21312 513439 21314
rect 165356 21256 513378 21312
rect 513434 21256 513439 21312
rect 165356 21254 513439 21256
rect 165356 21252 165362 21254
rect 513373 21251 513439 21254
rect 144126 20028 144132 20092
rect 144196 20090 144202 20092
rect 248413 20090 248479 20093
rect 144196 20088 248479 20090
rect 144196 20032 248418 20088
rect 248474 20032 248479 20088
rect 144196 20030 248479 20032
rect 144196 20028 144202 20030
rect 248413 20027 248479 20030
rect 148542 19892 148548 19956
rect 148612 19954 148618 19956
rect 300853 19954 300919 19957
rect 148612 19952 300919 19954
rect 148612 19896 300858 19952
rect 300914 19896 300919 19952
rect 148612 19894 300919 19896
rect 148612 19892 148618 19894
rect 300853 19891 300919 19894
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 140630 18668 140636 18732
rect 140700 18730 140706 18732
rect 191833 18730 191899 18733
rect 140700 18728 191899 18730
rect 140700 18672 191838 18728
rect 191894 18672 191899 18728
rect 140700 18670 191899 18672
rect 140700 18668 140706 18670
rect 191833 18667 191899 18670
rect 160870 18532 160876 18596
rect 160940 18594 160946 18596
rect 458173 18594 458239 18597
rect 160940 18592 458239 18594
rect 160940 18536 458178 18592
rect 458234 18536 458239 18592
rect 160940 18534 458239 18536
rect 160940 18532 160946 18534
rect 458173 18531 458239 18534
rect 152590 17308 152596 17372
rect 152660 17370 152666 17372
rect 350533 17370 350599 17373
rect 152660 17368 350599 17370
rect 152660 17312 350538 17368
rect 350594 17312 350599 17368
rect 152660 17310 350599 17312
rect 152660 17308 152666 17310
rect 350533 17307 350599 17310
rect 161054 17172 161060 17236
rect 161124 17234 161130 17236
rect 459553 17234 459619 17237
rect 161124 17232 459619 17234
rect 161124 17176 459558 17232
rect 459614 17176 459619 17232
rect 161124 17174 459619 17176
rect 161124 17172 161130 17174
rect 459553 17171 459619 17174
rect 137686 16356 137692 16420
rect 137756 16418 137762 16420
rect 158897 16418 158963 16421
rect 137756 16416 158963 16418
rect 137756 16360 158902 16416
rect 158958 16360 158963 16416
rect 137756 16358 158963 16360
rect 137756 16356 137762 16358
rect 158897 16355 158963 16358
rect 154062 16220 154068 16284
rect 154132 16282 154138 16284
rect 371233 16282 371299 16285
rect 154132 16280 371299 16282
rect 154132 16224 371238 16280
rect 371294 16224 371299 16280
rect 154132 16222 371299 16224
rect 154132 16220 154138 16222
rect 371233 16219 371299 16222
rect 157006 16084 157012 16148
rect 157076 16146 157082 16148
rect 407113 16146 407179 16149
rect 157076 16144 407179 16146
rect 157076 16088 407118 16144
rect 407174 16088 407179 16144
rect 157076 16086 407179 16088
rect 157076 16084 157082 16086
rect 407113 16083 407179 16086
rect 158294 15948 158300 16012
rect 158364 16010 158370 16012
rect 420913 16010 420979 16013
rect 158364 16008 420979 16010
rect 158364 15952 420918 16008
rect 420974 15952 420979 16008
rect 158364 15950 420979 15952
rect 158364 15948 158370 15950
rect 420913 15947 420979 15950
rect 158110 15812 158116 15876
rect 158180 15874 158186 15876
rect 423765 15874 423831 15877
rect 158180 15872 423831 15874
rect 158180 15816 423770 15872
rect 423826 15816 423831 15872
rect 158180 15814 423831 15816
rect 158180 15812 158186 15814
rect 423765 15811 423831 15814
rect 152774 14860 152780 14924
rect 152844 14922 152850 14924
rect 349153 14922 349219 14925
rect 152844 14920 349219 14922
rect 152844 14864 349158 14920
rect 349214 14864 349219 14920
rect 152844 14862 349219 14864
rect 152844 14860 152850 14862
rect 349153 14859 349219 14862
rect 155718 14724 155724 14788
rect 155788 14786 155794 14788
rect 387793 14786 387859 14789
rect 155788 14784 387859 14786
rect 155788 14728 387798 14784
rect 387854 14728 387859 14784
rect 155788 14726 387859 14728
rect 155788 14724 155794 14726
rect 387793 14723 387859 14726
rect 156638 14588 156644 14652
rect 156708 14650 156714 14652
rect 407205 14650 407271 14653
rect 156708 14648 407271 14650
rect 156708 14592 407210 14648
rect 407266 14592 407271 14648
rect 156708 14590 407271 14592
rect 156708 14588 156714 14590
rect 407205 14587 407271 14590
rect 163446 14452 163452 14516
rect 163516 14514 163522 14516
rect 495433 14514 495499 14517
rect 163516 14512 495499 14514
rect 163516 14456 495438 14512
rect 495494 14456 495499 14512
rect 163516 14454 495499 14456
rect 163516 14452 163522 14454
rect 495433 14451 495499 14454
rect 154246 12956 154252 13020
rect 154316 13018 154322 13020
rect 370129 13018 370195 13021
rect 154316 13016 370195 13018
rect 154316 12960 370134 13016
rect 370190 12960 370195 13016
rect 154316 12958 370195 12960
rect 154316 12956 154322 12958
rect 370129 12955 370195 12958
rect 140998 12140 141004 12204
rect 141068 12202 141074 12204
rect 213361 12202 213427 12205
rect 141068 12200 213427 12202
rect 141068 12144 213366 12200
rect 213422 12144 213427 12200
rect 141068 12142 213427 12144
rect 141068 12140 141074 12142
rect 213361 12139 213427 12142
rect 152406 12004 152412 12068
rect 152476 12066 152482 12068
rect 352833 12066 352899 12069
rect 152476 12064 352899 12066
rect 152476 12008 352838 12064
rect 352894 12008 352899 12064
rect 152476 12006 352899 12008
rect 152476 12004 152482 12006
rect 352833 12003 352899 12006
rect 153878 11868 153884 11932
rect 153948 11930 153954 11932
rect 372889 11930 372955 11933
rect 153948 11928 372955 11930
rect 153948 11872 372894 11928
rect 372950 11872 372955 11928
rect 153948 11870 372955 11872
rect 153948 11868 153954 11870
rect 372889 11867 372955 11870
rect 161238 11732 161244 11796
rect 161308 11794 161314 11796
rect 456885 11794 456951 11797
rect 161308 11792 456951 11794
rect 161308 11736 456890 11792
rect 456946 11736 456951 11792
rect 161308 11734 456951 11736
rect 161308 11732 161314 11734
rect 456885 11731 456951 11734
rect 74993 11658 75059 11661
rect 131246 11658 131252 11660
rect 74993 11656 131252 11658
rect 74993 11600 74998 11656
rect 75054 11600 131252 11656
rect 74993 11598 131252 11600
rect 74993 11595 75059 11598
rect 131246 11596 131252 11598
rect 131316 11596 131322 11660
rect 170622 11596 170628 11660
rect 170692 11658 170698 11660
rect 580993 11658 581059 11661
rect 170692 11656 581059 11658
rect 170692 11600 580998 11656
rect 581054 11600 581059 11656
rect 170692 11598 581059 11600
rect 170692 11596 170698 11598
rect 580993 11595 581059 11598
rect 114001 10570 114067 10573
rect 134190 10570 134196 10572
rect 114001 10568 134196 10570
rect 114001 10512 114006 10568
rect 114062 10512 134196 10568
rect 114001 10510 134196 10512
rect 114001 10507 114067 10510
rect 134190 10508 134196 10510
rect 134260 10508 134266 10572
rect 110505 10434 110571 10437
rect 134006 10434 134012 10436
rect 110505 10432 134012 10434
rect 110505 10376 110510 10432
rect 110566 10376 134012 10432
rect 110505 10374 134012 10376
rect 110505 10371 110571 10374
rect 134006 10372 134012 10374
rect 134076 10372 134082 10436
rect 151302 10372 151308 10436
rect 151372 10434 151378 10436
rect 334617 10434 334683 10437
rect 151372 10432 334683 10434
rect 151372 10376 334622 10432
rect 334678 10376 334683 10432
rect 151372 10374 334683 10376
rect 151372 10372 151378 10374
rect 334617 10371 334683 10374
rect 92473 10298 92539 10301
rect 133270 10298 133276 10300
rect 92473 10296 133276 10298
rect 92473 10240 92478 10296
rect 92534 10240 133276 10296
rect 92473 10238 133276 10240
rect 92473 10235 92539 10238
rect 133270 10236 133276 10238
rect 133340 10236 133346 10300
rect 151486 10236 151492 10300
rect 151556 10298 151562 10300
rect 336273 10298 336339 10301
rect 151556 10296 336339 10298
rect 151556 10240 336278 10296
rect 336334 10240 336339 10296
rect 151556 10238 336339 10240
rect 151556 10236 151562 10238
rect 336273 10235 336339 10238
rect 109309 9346 109375 9349
rect 134374 9346 134380 9348
rect 109309 9344 134380 9346
rect 109309 9288 109314 9344
rect 109370 9288 134380 9344
rect 109309 9286 134380 9288
rect 109309 9283 109375 9286
rect 134374 9284 134380 9286
rect 134444 9284 134450 9348
rect 147070 9284 147076 9348
rect 147140 9346 147146 9348
rect 281901 9346 281967 9349
rect 147140 9344 281967 9346
rect 147140 9288 281906 9344
rect 281962 9288 281967 9344
rect 147140 9286 281967 9288
rect 147140 9284 147146 9286
rect 281901 9283 281967 9286
rect 57237 9210 57303 9213
rect 129958 9210 129964 9212
rect 57237 9208 129964 9210
rect 57237 9152 57242 9208
rect 57298 9152 129964 9208
rect 57237 9150 129964 9152
rect 57237 9147 57303 9150
rect 129958 9148 129964 9150
rect 130028 9148 130034 9212
rect 148910 9148 148916 9212
rect 148980 9210 148986 9212
rect 300761 9210 300827 9213
rect 148980 9208 300827 9210
rect 148980 9152 300766 9208
rect 300822 9152 300827 9208
rect 148980 9150 300827 9152
rect 148980 9148 148986 9150
rect 300761 9147 300827 9150
rect 41873 9074 41939 9077
rect 128670 9074 128676 9076
rect 41873 9072 128676 9074
rect 41873 9016 41878 9072
rect 41934 9016 128676 9072
rect 41873 9014 128676 9016
rect 41873 9011 41939 9014
rect 128670 9012 128676 9014
rect 128740 9012 128746 9076
rect 148726 9012 148732 9076
rect 148796 9074 148802 9076
rect 299657 9074 299723 9077
rect 148796 9072 299723 9074
rect 148796 9016 299662 9072
rect 299718 9016 299723 9072
rect 148796 9014 299723 9016
rect 148796 9012 148802 9014
rect 299657 9011 299723 9014
rect 38377 8938 38443 8941
rect 128854 8938 128860 8940
rect 38377 8936 128860 8938
rect 38377 8880 38382 8936
rect 38438 8880 128860 8936
rect 38377 8878 128860 8880
rect 38377 8875 38443 8878
rect 128854 8876 128860 8878
rect 128924 8876 128930 8940
rect 165102 8876 165108 8940
rect 165172 8938 165178 8940
rect 511257 8938 511323 8941
rect 165172 8936 511323 8938
rect 165172 8880 511262 8936
rect 511318 8880 511323 8936
rect 165172 8878 511323 8880
rect 165172 8876 165178 8878
rect 511257 8875 511323 8878
rect 145414 8060 145420 8124
rect 145484 8122 145490 8124
rect 264145 8122 264211 8125
rect 145484 8120 264211 8122
rect 145484 8064 264150 8120
rect 264206 8064 264211 8120
rect 145484 8062 264211 8064
rect 145484 8060 145490 8062
rect 264145 8059 264211 8062
rect 145598 7924 145604 7988
rect 145668 7986 145674 7988
rect 265341 7986 265407 7989
rect 145668 7984 265407 7986
rect 145668 7928 265346 7984
rect 265402 7928 265407 7984
rect 145668 7926 265407 7928
rect 145668 7924 145674 7926
rect 265341 7923 265407 7926
rect 151670 7788 151676 7852
rect 151740 7850 151746 7852
rect 337469 7850 337535 7853
rect 151740 7848 337535 7850
rect 151740 7792 337474 7848
rect 337530 7792 337535 7848
rect 151740 7790 337535 7792
rect 151740 7788 151746 7790
rect 337469 7787 337535 7790
rect 91553 7714 91619 7717
rect 133086 7714 133092 7716
rect 91553 7712 133092 7714
rect 91553 7656 91558 7712
rect 91614 7656 133092 7712
rect 91553 7654 133092 7656
rect 91553 7651 91619 7654
rect 133086 7652 133092 7654
rect 133156 7652 133162 7716
rect 158478 7652 158484 7716
rect 158548 7714 158554 7716
rect 424961 7714 425027 7717
rect 158548 7712 425027 7714
rect 158548 7656 424966 7712
rect 425022 7656 425027 7712
rect 158548 7654 425027 7656
rect 158548 7652 158554 7654
rect 424961 7651 425027 7654
rect 56041 7578 56107 7581
rect 130142 7578 130148 7580
rect 56041 7576 130148 7578
rect 56041 7520 56046 7576
rect 56102 7520 130148 7576
rect 56041 7518 130148 7520
rect 56041 7515 56107 7518
rect 130142 7516 130148 7518
rect 130212 7516 130218 7580
rect 162158 7516 162164 7580
rect 162228 7578 162234 7580
rect 478229 7578 478295 7581
rect 162228 7576 478295 7578
rect 162228 7520 478234 7576
rect 478290 7520 478295 7576
rect 162228 7518 478295 7520
rect 162228 7516 162234 7518
rect 478229 7515 478295 7518
rect 88149 6626 88215 6629
rect 127198 6626 127204 6628
rect 88149 6624 127204 6626
rect -960 6490 480 6580
rect 88149 6568 88154 6624
rect 88210 6568 127204 6624
rect 88149 6566 127204 6568
rect 88149 6563 88215 6566
rect 127198 6564 127204 6566
rect 127268 6564 127274 6628
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3509 6490 3575 6493
rect -960 6488 3575 6490
rect -960 6432 3514 6488
rect 3570 6432 3575 6488
rect -960 6430 3575 6432
rect -960 6340 480 6430
rect 3509 6427 3575 6430
rect 73797 6490 73863 6493
rect 131062 6490 131068 6492
rect 73797 6488 131068 6490
rect 73797 6432 73802 6488
rect 73858 6432 131068 6488
rect 73797 6430 131068 6432
rect 73797 6427 73863 6430
rect 131062 6428 131068 6430
rect 131132 6428 131138 6492
rect 583520 6476 584960 6566
rect 40677 6354 40743 6357
rect 128670 6354 128676 6356
rect 40677 6352 128676 6354
rect 40677 6296 40682 6352
rect 40738 6296 128676 6352
rect 40677 6294 128676 6296
rect 40677 6291 40743 6294
rect 128670 6292 128676 6294
rect 128740 6292 128746 6356
rect 20621 6218 20687 6221
rect 127382 6218 127388 6220
rect 20621 6216 127388 6218
rect 20621 6160 20626 6216
rect 20682 6160 127388 6216
rect 20621 6158 127388 6160
rect 20621 6155 20687 6158
rect 127382 6156 127388 6158
rect 127452 6156 127458 6220
rect 142838 6156 142844 6220
rect 142908 6218 142914 6220
rect 228725 6218 228791 6221
rect 142908 6216 228791 6218
rect 142908 6160 228730 6216
rect 228786 6160 228791 6216
rect 142908 6158 228791 6160
rect 142908 6156 142914 6158
rect 228725 6155 228791 6158
rect 166758 4932 166764 4996
rect 166828 4994 166834 4996
rect 532509 4994 532575 4997
rect 166828 4992 532575 4994
rect 166828 4936 532514 4992
rect 532570 4936 532575 4992
rect 166828 4934 532575 4936
rect 166828 4932 166834 4934
rect 532509 4931 532575 4934
rect 137870 4796 137876 4860
rect 137940 4858 137946 4860
rect 160093 4858 160159 4861
rect 137940 4856 160159 4858
rect 137940 4800 160098 4856
rect 160154 4800 160159 4856
rect 137940 4798 160159 4800
rect 137940 4796 137946 4798
rect 160093 4795 160159 4798
rect 168046 4796 168052 4860
rect 168116 4858 168122 4860
rect 547873 4858 547939 4861
rect 168116 4856 547939 4858
rect 168116 4800 547878 4856
rect 547934 4800 547939 4856
rect 168116 4798 547939 4800
rect 168116 4796 168122 4798
rect 547873 4795 547939 4798
rect 163630 3436 163636 3500
rect 163700 3498 163706 3500
rect 494697 3498 494763 3501
rect 163700 3496 494763 3498
rect 163700 3440 494702 3496
rect 494758 3440 494763 3496
rect 163700 3438 494763 3440
rect 163700 3436 163706 3438
rect 494697 3435 494763 3438
rect 4061 3362 4127 3365
rect 125910 3362 125916 3364
rect 4061 3360 125916 3362
rect 4061 3304 4066 3360
rect 4122 3304 125916 3360
rect 4061 3302 125916 3304
rect 4061 3299 4127 3302
rect 125910 3300 125916 3302
rect 125980 3300 125986 3364
rect 128169 3362 128235 3365
rect 135662 3362 135668 3364
rect 128169 3360 135668 3362
rect 128169 3304 128174 3360
rect 128230 3304 135668 3360
rect 128169 3302 135668 3304
rect 128169 3299 128235 3302
rect 135662 3300 135668 3302
rect 135732 3300 135738 3364
rect 136398 3300 136404 3364
rect 136468 3362 136474 3364
rect 161289 3362 161355 3365
rect 136468 3360 161355 3362
rect 136468 3304 161294 3360
rect 161350 3304 161355 3360
rect 136468 3302 161355 3304
rect 136468 3300 136474 3302
rect 161289 3299 161355 3302
rect 171726 3300 171732 3364
rect 171796 3362 171802 3364
rect 554957 3362 555023 3365
rect 171796 3360 555023 3362
rect 171796 3304 554962 3360
rect 555018 3304 555023 3360
rect 171796 3302 555023 3304
rect 171796 3300 171802 3302
rect 554957 3299 555023 3302
<< via3 >>
rect 3372 658140 3436 658204
rect 396764 643724 396828 643788
rect 396580 643180 396644 643244
rect 396764 227700 396828 227764
rect 144868 190980 144932 191044
rect 141004 190300 141068 190364
rect 146156 188532 146220 188596
rect 141740 184316 141804 184380
rect 140820 184240 140884 184244
rect 140820 184184 140834 184240
rect 140834 184184 140884 184240
rect 140820 184180 140884 184184
rect 142844 184044 142908 184108
rect 144868 182200 144932 182204
rect 144868 182144 144918 182200
rect 144918 182144 144932 182200
rect 144868 182140 144932 182144
rect 145052 181188 145116 181252
rect 152596 181188 152660 181252
rect 142476 180916 142540 180980
rect 142844 178876 142908 178940
rect 141004 178740 141068 178804
rect 141740 178800 141804 178804
rect 141740 178744 141790 178800
rect 141790 178744 141804 178800
rect 141740 178740 141804 178744
rect 140820 178604 140884 178668
rect 145052 177380 145116 177444
rect 158668 176428 158732 176492
rect 142476 172952 142540 172956
rect 142476 172896 142526 172952
rect 142526 172896 142540 172952
rect 142476 172892 142540 172896
rect 158668 172892 158732 172956
rect 152596 169492 152660 169556
rect 146156 157932 146220 157996
rect 153516 78508 153580 78572
rect 164004 78508 164068 78572
rect 165292 78508 165356 78572
rect 173572 78508 173636 78572
rect 162164 78372 162228 78436
rect 171364 78372 171428 78436
rect 171548 78372 171612 78436
rect 130700 77964 130764 78028
rect 131068 77964 131132 78028
rect 144868 77964 144932 78028
rect 3372 77828 3436 77892
rect 126652 77828 126716 77892
rect 128676 77828 128740 77892
rect 129596 77828 129660 77892
rect 130516 77888 130580 77892
rect 130516 77832 130520 77888
rect 130520 77832 130576 77888
rect 130576 77832 130580 77888
rect 130516 77828 130580 77832
rect 131436 77828 131500 77892
rect 131988 77888 132052 77892
rect 131988 77832 131992 77888
rect 131992 77832 132048 77888
rect 132048 77832 132052 77888
rect 131988 77828 132052 77832
rect 132540 77888 132604 77892
rect 132540 77832 132544 77888
rect 132544 77832 132600 77888
rect 132600 77832 132604 77888
rect 132540 77828 132604 77832
rect 132908 77888 132972 77892
rect 132908 77832 132912 77888
rect 132912 77832 132968 77888
rect 132968 77832 132972 77888
rect 132908 77828 132972 77832
rect 134196 77828 134260 77892
rect 136036 77888 136100 77892
rect 136036 77832 136040 77888
rect 136040 77832 136096 77888
rect 136096 77832 136100 77888
rect 136036 77828 136100 77832
rect 136404 77888 136468 77892
rect 136404 77832 136408 77888
rect 136408 77832 136464 77888
rect 136464 77832 136468 77888
rect 136404 77828 136468 77832
rect 130700 77692 130764 77756
rect 133092 77692 133156 77756
rect 135300 77692 135364 77756
rect 136956 77692 137020 77756
rect 144684 77828 144748 77892
rect 145420 78100 145484 78164
rect 155172 78236 155236 78300
rect 163820 78236 163884 78300
rect 164004 78236 164068 78300
rect 169340 78100 169404 78164
rect 145236 77964 145300 78028
rect 155172 77964 155236 78028
rect 145236 77828 145300 77892
rect 138612 77692 138676 77756
rect 131436 77480 131500 77484
rect 131436 77424 131450 77480
rect 131450 77424 131500 77480
rect 131436 77420 131500 77424
rect 131988 77480 132052 77484
rect 131988 77424 132038 77480
rect 132038 77424 132052 77480
rect 131988 77420 132052 77424
rect 136404 77420 136468 77484
rect 137692 77420 137756 77484
rect 140636 77556 140700 77620
rect 145052 77692 145116 77756
rect 145236 77692 145300 77756
rect 144868 77556 144932 77620
rect 144868 77420 144932 77484
rect 151492 77828 151556 77892
rect 152044 77888 152108 77892
rect 152044 77832 152048 77888
rect 152048 77832 152104 77888
rect 152104 77832 152108 77888
rect 152044 77828 152108 77832
rect 152780 77888 152844 77892
rect 152780 77832 152784 77888
rect 152784 77832 152840 77888
rect 152840 77832 152844 77888
rect 152780 77828 152844 77832
rect 153378 77888 153442 77892
rect 153378 77832 153428 77888
rect 153428 77832 153442 77888
rect 153378 77828 153442 77832
rect 153700 77888 153764 77892
rect 153700 77832 153704 77888
rect 153704 77832 153760 77888
rect 153760 77832 153764 77888
rect 153700 77828 153764 77832
rect 154068 77888 154132 77892
rect 154068 77832 154072 77888
rect 154072 77832 154128 77888
rect 154128 77832 154132 77888
rect 154068 77828 154132 77832
rect 154252 77828 154316 77892
rect 154988 77888 155052 77892
rect 154988 77832 154992 77888
rect 154992 77832 155048 77888
rect 155048 77832 155052 77888
rect 154988 77828 155052 77832
rect 152412 77692 152476 77756
rect 153148 77616 153212 77620
rect 153148 77560 153198 77616
rect 153198 77560 153212 77616
rect 153148 77556 153212 77560
rect 154252 77616 154316 77620
rect 154252 77560 154266 77616
rect 154266 77560 154316 77616
rect 154252 77556 154316 77560
rect 145420 77480 145484 77484
rect 145420 77424 145470 77480
rect 145470 77424 145484 77480
rect 145420 77420 145484 77424
rect 156092 77692 156156 77756
rect 156828 77828 156892 77892
rect 156644 77692 156708 77756
rect 158116 77828 158180 77892
rect 158668 77888 158732 77892
rect 158668 77832 158672 77888
rect 158672 77832 158728 77888
rect 158728 77832 158732 77888
rect 158668 77828 158732 77832
rect 158484 77752 158548 77756
rect 158484 77696 158534 77752
rect 158534 77696 158548 77752
rect 158484 77692 158548 77696
rect 156276 77556 156340 77620
rect 158300 77616 158364 77620
rect 158300 77560 158314 77616
rect 158314 77560 158364 77616
rect 158300 77556 158364 77560
rect 162164 77828 162228 77892
rect 162716 77866 162720 77892
rect 162720 77866 162776 77892
rect 162776 77866 162780 77892
rect 162716 77828 162780 77866
rect 163084 77888 163148 77892
rect 163084 77832 163088 77888
rect 163088 77832 163144 77888
rect 163144 77832 163148 77888
rect 163084 77828 163148 77832
rect 163268 77828 163332 77892
rect 163636 77828 163700 77892
rect 164372 77828 164436 77892
rect 164924 77828 164988 77892
rect 165108 77828 165172 77892
rect 165476 77866 165480 77892
rect 165480 77866 165536 77892
rect 165536 77866 165540 77892
rect 165476 77828 165540 77866
rect 165844 77888 165908 77892
rect 165844 77832 165848 77888
rect 165848 77832 165904 77888
rect 165904 77832 165908 77888
rect 165844 77828 165908 77832
rect 166764 77828 166828 77892
rect 167316 77964 167380 78028
rect 167684 77964 167748 78028
rect 167500 77866 167504 77892
rect 167504 77866 167560 77892
rect 167560 77866 167564 77892
rect 167500 77828 167564 77866
rect 160324 77692 160388 77756
rect 160692 77752 160756 77756
rect 160692 77696 160696 77752
rect 160696 77696 160752 77752
rect 160752 77696 160756 77752
rect 160692 77692 160756 77696
rect 161244 77692 161308 77756
rect 162716 77692 162780 77756
rect 163820 77692 163884 77756
rect 168604 77888 168668 77892
rect 168604 77832 168608 77888
rect 168608 77832 168664 77888
rect 168664 77832 168668 77888
rect 168604 77828 168668 77832
rect 164556 77556 164620 77620
rect 166028 77556 166092 77620
rect 166580 77556 166644 77620
rect 170076 77888 170140 77892
rect 170076 77832 170080 77888
rect 170080 77832 170136 77888
rect 170136 77832 170140 77888
rect 170076 77828 170140 77832
rect 170260 77866 170264 77892
rect 170264 77866 170320 77892
rect 170320 77866 170324 77892
rect 170260 77828 170324 77866
rect 170628 77888 170692 77892
rect 170628 77832 170632 77888
rect 170632 77832 170688 77888
rect 170688 77832 170692 77888
rect 170628 77828 170692 77832
rect 170996 77888 171060 77892
rect 170996 77832 171000 77888
rect 171000 77832 171056 77888
rect 171056 77832 171060 77888
rect 170996 77828 171060 77832
rect 171916 77828 171980 77892
rect 170812 77692 170876 77756
rect 172468 77828 172532 77892
rect 173020 77828 173084 77892
rect 396580 77692 396644 77756
rect 173572 77616 173636 77620
rect 173572 77560 173622 77616
rect 173622 77560 173636 77616
rect 173572 77556 173636 77560
rect 164372 77420 164436 77484
rect 165292 77420 165356 77484
rect 169340 77420 169404 77484
rect 172100 77480 172164 77484
rect 172100 77424 172150 77480
rect 172150 77424 172164 77480
rect 172100 77420 172164 77424
rect 171548 77344 171612 77348
rect 171548 77288 171562 77344
rect 171562 77288 171612 77344
rect 171548 77284 171612 77288
rect 132540 77208 132604 77212
rect 132540 77152 132554 77208
rect 132554 77152 132604 77208
rect 132540 77148 132604 77152
rect 153516 77148 153580 77212
rect 153884 77208 153948 77212
rect 153884 77152 153898 77208
rect 153898 77152 153948 77208
rect 153884 77148 153948 77152
rect 170996 77148 171060 77212
rect 154988 77012 155052 77076
rect 156092 77012 156156 77076
rect 164924 77012 164988 77076
rect 166396 77012 166460 77076
rect 127204 76800 127268 76804
rect 127204 76744 127254 76800
rect 127254 76744 127268 76800
rect 127204 76740 127268 76744
rect 129044 76740 129108 76804
rect 147260 76800 147324 76804
rect 147260 76744 147310 76800
rect 147310 76744 147324 76800
rect 147260 76740 147324 76744
rect 153332 76740 153396 76804
rect 154436 76740 154500 76804
rect 155724 76800 155788 76804
rect 155724 76744 155738 76800
rect 155738 76744 155788 76800
rect 155724 76740 155788 76744
rect 167500 76740 167564 76804
rect 168052 76800 168116 76804
rect 168052 76744 168102 76800
rect 168102 76744 168116 76800
rect 168052 76740 168116 76744
rect 127388 76332 127452 76396
rect 128676 76332 128740 76396
rect 129780 76392 129844 76396
rect 129780 76336 129794 76392
rect 129794 76336 129844 76392
rect 129780 76332 129844 76336
rect 129964 76392 130028 76396
rect 129964 76336 130014 76392
rect 130014 76336 130028 76392
rect 129964 76332 130028 76336
rect 132908 76332 132972 76396
rect 134380 76392 134444 76396
rect 134380 76336 134394 76392
rect 134394 76336 134444 76392
rect 134380 76332 134444 76336
rect 138980 76392 139044 76396
rect 138980 76336 139030 76392
rect 139030 76336 139044 76392
rect 138980 76332 139044 76336
rect 139164 76332 139228 76396
rect 145604 76332 145668 76396
rect 153332 76332 153396 76396
rect 162532 76392 162596 76396
rect 162532 76336 162582 76392
rect 162582 76336 162596 76392
rect 162532 76332 162596 76336
rect 167500 76332 167564 76396
rect 168604 76332 168668 76396
rect 169340 76332 169404 76396
rect 171364 76332 171428 76396
rect 133092 76196 133156 76260
rect 145420 76196 145484 76260
rect 149836 76196 149900 76260
rect 154068 76196 154132 76260
rect 162348 76196 162412 76260
rect 163452 76196 163516 76260
rect 166212 76196 166276 76260
rect 173020 76256 173084 76260
rect 173020 76200 173034 76256
rect 173034 76200 173084 76256
rect 173020 76196 173084 76200
rect 128492 76060 128556 76124
rect 152596 76060 152660 76124
rect 157932 76060 157996 76124
rect 172468 76060 172532 76124
rect 152412 75924 152476 75988
rect 160692 75924 160756 75988
rect 163084 75924 163148 75988
rect 128860 75788 128924 75852
rect 153884 75788 153948 75852
rect 167868 75788 167932 75852
rect 130700 75652 130764 75716
rect 148916 75712 148980 75716
rect 148916 75656 148930 75712
rect 148930 75656 148980 75712
rect 148916 75652 148980 75656
rect 149652 75652 149716 75716
rect 128676 75576 128740 75580
rect 128676 75520 128726 75576
rect 128726 75520 128740 75576
rect 128676 75516 128740 75520
rect 151308 75652 151372 75716
rect 152412 75652 152476 75716
rect 154252 75712 154316 75716
rect 154252 75656 154302 75712
rect 154302 75656 154316 75712
rect 154252 75652 154316 75656
rect 156276 75652 156340 75716
rect 157012 75652 157076 75716
rect 158668 75652 158732 75716
rect 154068 75516 154132 75580
rect 160876 75516 160940 75580
rect 161060 75516 161124 75580
rect 163268 75516 163332 75580
rect 170076 75652 170140 75716
rect 170996 75652 171060 75716
rect 130516 75380 130580 75444
rect 153332 75304 153396 75308
rect 153332 75248 153346 75304
rect 153346 75248 153396 75304
rect 153332 75244 153396 75248
rect 164556 75304 164620 75308
rect 164556 75248 164570 75304
rect 164570 75248 164620 75304
rect 164556 75244 164620 75248
rect 125916 75108 125980 75172
rect 144132 75108 144196 75172
rect 159036 75108 159100 75172
rect 164740 75108 164804 75172
rect 133092 74972 133156 75036
rect 134012 75032 134076 75036
rect 134012 74976 134062 75032
rect 134062 74976 134076 75032
rect 134012 74972 134076 74976
rect 135668 74972 135732 75036
rect 136036 75032 136100 75036
rect 136036 74976 136086 75032
rect 136086 74976 136100 75032
rect 136036 74972 136100 74976
rect 137876 75032 137940 75036
rect 137876 74976 137926 75032
rect 137926 74976 137940 75032
rect 137876 74972 137940 74976
rect 138796 74972 138860 75036
rect 140084 74972 140148 75036
rect 140452 74972 140516 75036
rect 144500 74972 144564 75036
rect 145236 74972 145300 75036
rect 148732 75032 148796 75036
rect 148732 74976 148782 75032
rect 148782 74976 148796 75032
rect 148732 74972 148796 74976
rect 152044 74972 152108 75036
rect 158852 74972 158916 75036
rect 170260 75032 170324 75036
rect 170260 74976 170274 75032
rect 170274 74976 170324 75032
rect 170260 74972 170324 74976
rect 131436 74836 131500 74900
rect 140268 74836 140332 74900
rect 142844 74836 142908 74900
rect 131068 74700 131132 74764
rect 143028 74700 143092 74764
rect 143396 74760 143460 74764
rect 143396 74704 143446 74760
rect 143446 74704 143460 74760
rect 143396 74700 143460 74704
rect 167316 74700 167380 74764
rect 131252 74624 131316 74628
rect 131252 74568 131302 74624
rect 131302 74568 131316 74624
rect 131252 74564 131316 74568
rect 141004 74564 141068 74628
rect 143212 74564 143276 74628
rect 148548 74564 148612 74628
rect 171732 74700 171796 74764
rect 133276 74428 133340 74492
rect 160508 74488 160572 74492
rect 160508 74432 160522 74488
rect 160522 74432 160572 74488
rect 160508 74428 160572 74432
rect 138612 73884 138676 73948
rect 136404 73748 136468 73812
rect 147076 73476 147140 73540
rect 166028 73476 166092 73540
rect 136588 73340 136652 73404
rect 171916 73204 171980 73268
rect 160324 73068 160388 73132
rect 151676 72856 151740 72860
rect 151676 72800 151726 72856
rect 151726 72800 151740 72856
rect 151676 72796 151740 72800
rect 129780 72524 129844 72588
rect 131436 71844 131500 71908
rect 135300 71708 135364 71772
rect 143396 71436 143460 71500
rect 126652 71360 126716 71364
rect 126652 71304 126666 71360
rect 126666 71304 126716 71360
rect 126652 71300 126716 71304
rect 144868 71300 144932 71364
rect 129044 71028 129108 71092
rect 170996 71028 171060 71092
rect 165844 70892 165908 70956
rect 164924 70348 164988 70412
rect 162716 69940 162780 70004
rect 154436 68172 154500 68236
rect 152964 66812 153028 66876
rect 138796 65452 138860 65516
rect 138980 63004 139044 63068
rect 140084 62868 140148 62932
rect 166212 62732 166276 62796
rect 158852 59876 158916 59940
rect 140268 57292 140332 57356
rect 144500 57156 144564 57220
rect 156828 54436 156892 54500
rect 171916 50220 171980 50284
rect 162348 39204 162412 39268
rect 157932 36484 157996 36548
rect 147260 35260 147324 35324
rect 149836 35124 149900 35188
rect 139164 33900 139228 33964
rect 143028 33764 143092 33828
rect 166396 32676 166460 32740
rect 167684 32540 167748 32604
rect 167500 32404 167564 32468
rect 160692 30908 160756 30972
rect 162532 29548 162596 29612
rect 143212 28188 143276 28252
rect 140452 26964 140516 27028
rect 169340 26828 169404 26892
rect 149652 25468 149716 25532
rect 167868 24244 167932 24308
rect 170812 24108 170876 24172
rect 166580 22612 166644 22676
rect 159036 21388 159100 21452
rect 165292 21252 165356 21316
rect 144132 20028 144196 20092
rect 148548 19892 148612 19956
rect 140636 18668 140700 18732
rect 160876 18532 160940 18596
rect 152596 17308 152660 17372
rect 161060 17172 161124 17236
rect 137692 16356 137756 16420
rect 154068 16220 154132 16284
rect 157012 16084 157076 16148
rect 158300 15948 158364 16012
rect 158116 15812 158180 15876
rect 152780 14860 152844 14924
rect 155724 14724 155788 14788
rect 156644 14588 156708 14652
rect 163452 14452 163516 14516
rect 154252 12956 154316 13020
rect 141004 12140 141068 12204
rect 152412 12004 152476 12068
rect 153884 11868 153948 11932
rect 161244 11732 161308 11796
rect 131252 11596 131316 11660
rect 170628 11596 170692 11660
rect 134196 10508 134260 10572
rect 134012 10372 134076 10436
rect 151308 10372 151372 10436
rect 133276 10236 133340 10300
rect 151492 10236 151556 10300
rect 134380 9284 134444 9348
rect 147076 9284 147140 9348
rect 129964 9148 130028 9212
rect 148916 9148 148980 9212
rect 128676 9012 128740 9076
rect 148732 9012 148796 9076
rect 128860 8876 128924 8940
rect 165108 8876 165172 8940
rect 145420 8060 145484 8124
rect 145604 7924 145668 7988
rect 151676 7788 151740 7852
rect 133092 7652 133156 7716
rect 158484 7652 158548 7716
rect 130148 7516 130212 7580
rect 162164 7516 162228 7580
rect 127204 6564 127268 6628
rect 131068 6428 131132 6492
rect 128676 6292 128740 6356
rect 127388 6156 127452 6220
rect 142844 6156 142908 6220
rect 166764 4932 166828 4996
rect 137876 4796 137940 4860
rect 168052 4796 168116 4860
rect 163636 3436 163700 3500
rect 125916 3300 125980 3364
rect 135668 3300 135732 3364
rect 136404 3300 136468 3364
rect 171732 3300 171796 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 3371 658204 3437 658205
rect 3371 658140 3372 658204
rect 3436 658140 3437 658204
rect 3371 658139 3437 658140
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 3374 77893 3434 658139
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 3371 77892 3437 77893
rect 3371 77828 3372 77892
rect 3436 77828 3437 77892
rect 3371 77827 3437 77828
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 248684 47414 263898
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 248684 51914 268398
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 248684 56414 272898
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 248684 60914 277398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 248684 65414 281898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 248684 69914 250398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 248684 74414 254898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 248684 78914 259398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 248684 83414 263898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 248684 87914 268398
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 248684 92414 272898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 248684 96914 277398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 248684 101414 281898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 248684 105914 250398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 248684 110414 254898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 248684 114914 259398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 248684 119414 263898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 248684 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 248684 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 248684 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 248684 137414 281898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 248684 141914 250398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 248684 146414 254898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 248684 150914 259398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 248684 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 248684 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 248684 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 248684 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 248684 173414 281898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 248684 177914 250398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 248684 182414 254898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 248684 186914 259398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 248684 191414 263898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 248684 195914 268398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 248684 200414 272898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 248684 204914 277398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 248684 209414 281898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 248684 213914 250398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 248684 218414 254898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 248684 222914 259398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 248684 227414 263898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 248684 231914 268398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 248684 236414 272898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 248684 240914 277398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 248684 245414 281898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 248684 249914 250398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 248684 254414 254898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 248684 258914 259398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 248684 263414 263898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 248684 267914 268398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 248684 272414 272898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 248684 276914 277398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 248684 281414 281898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 248684 285914 250398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 248684 290414 254898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 248684 294914 259398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 248684 299414 263898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 248684 303914 268398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 248684 308414 272898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 248684 312914 277398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 248684 317414 281898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 248684 321914 250398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 248684 326414 254898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 248684 330914 259398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 248684 335414 263898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 248684 339914 268398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 248684 344414 272898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 248684 348914 277398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 248684 353414 281898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 248684 357914 250398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 248684 362414 254898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 248684 366914 259398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 248684 371414 263898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 248684 375914 268398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 248684 380414 272898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 248684 384914 277398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 248684 389414 281898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 396763 643788 396829 643789
rect 396763 643724 396764 643788
rect 396828 643724 396829 643788
rect 396763 643723 396829 643724
rect 396579 643244 396645 643245
rect 396579 643180 396580 643244
rect 396644 643180 396645 643244
rect 396579 643179 396645 643180
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 248684 393914 250398
rect 65300 246303 70100 246486
rect 65300 246067 65342 246303
rect 65578 246067 65662 246303
rect 65898 246067 65982 246303
rect 66218 246067 66302 246303
rect 66538 246067 66622 246303
rect 66858 246067 66942 246303
rect 67178 246067 67262 246303
rect 67498 246067 67582 246303
rect 67818 246067 67902 246303
rect 68138 246067 68222 246303
rect 68458 246067 68542 246303
rect 68778 246067 68862 246303
rect 69098 246067 69182 246303
rect 69418 246067 69502 246303
rect 69738 246067 69822 246303
rect 70058 246067 70100 246303
rect 65300 245884 70100 246067
rect 65300 241953 71300 241984
rect 65300 241717 65462 241953
rect 65698 241717 65782 241953
rect 66018 241717 66102 241953
rect 66338 241717 66422 241953
rect 66658 241717 66742 241953
rect 66978 241717 67062 241953
rect 67298 241717 67382 241953
rect 67618 241717 67702 241953
rect 67938 241717 68022 241953
rect 68258 241717 68342 241953
rect 68578 241717 68662 241953
rect 68898 241717 68982 241953
rect 69218 241717 69302 241953
rect 69538 241717 69622 241953
rect 69858 241717 69942 241953
rect 70178 241717 70262 241953
rect 70498 241717 70582 241953
rect 70818 241717 70902 241953
rect 71138 241717 71300 241953
rect 65300 241633 71300 241717
rect 65300 241397 65462 241633
rect 65698 241397 65782 241633
rect 66018 241397 66102 241633
rect 66338 241397 66422 241633
rect 66658 241397 66742 241633
rect 66978 241397 67062 241633
rect 67298 241397 67382 241633
rect 67618 241397 67702 241633
rect 67938 241397 68022 241633
rect 68258 241397 68342 241633
rect 68578 241397 68662 241633
rect 68898 241397 68982 241633
rect 69218 241397 69302 241633
rect 69538 241397 69622 241633
rect 69858 241397 69942 241633
rect 70178 241397 70262 241633
rect 70498 241397 70582 241633
rect 70818 241397 70902 241633
rect 71138 241397 71300 241633
rect 65300 241366 71300 241397
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 228453 47414 228484
rect 46794 228217 46826 228453
rect 47062 228217 47146 228453
rect 47382 228217 47414 228453
rect 46794 228133 47414 228217
rect 46794 227897 46826 228133
rect 47062 227897 47146 228133
rect 47382 227897 47414 228133
rect 46794 192454 47414 227897
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 196954 51914 228484
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 201454 56414 228484
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 205954 60914 228484
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 210454 65414 228484
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 214954 69914 228484
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 219454 74414 228484
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 223954 78914 228484
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 228453 83414 228484
rect 82794 228217 82826 228453
rect 83062 228217 83146 228453
rect 83382 228217 83414 228453
rect 82794 228133 83414 228217
rect 82794 227897 82826 228133
rect 83062 227897 83146 228133
rect 83382 227897 83414 228133
rect 82794 192454 83414 227897
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 196954 87914 228484
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 201454 92414 228484
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 205954 96914 228484
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 210454 101414 228484
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 214954 105914 228484
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 219454 110414 228484
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 223954 114914 228484
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 118794 228453 119414 228484
rect 118794 228217 118826 228453
rect 119062 228217 119146 228453
rect 119382 228217 119414 228453
rect 118794 228133 119414 228217
rect 118794 227897 118826 228133
rect 119062 227897 119146 228133
rect 119382 227897 119414 228133
rect 118794 192454 119414 227897
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 140000 119414 155898
rect 123294 196954 123914 228484
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 140000 123914 160398
rect 127794 201454 128414 228484
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 140000 128414 164898
rect 132294 205954 132914 228484
rect 172794 210454 173414 228484
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 135914 205861 165514 205986
rect 135914 205625 136036 205861
rect 136272 205625 136356 205861
rect 136592 205625 136676 205861
rect 136912 205625 136996 205861
rect 137232 205625 137316 205861
rect 137552 205625 137636 205861
rect 137872 205625 137956 205861
rect 138192 205625 138276 205861
rect 138512 205625 138596 205861
rect 138832 205625 138916 205861
rect 139152 205625 139236 205861
rect 139472 205625 139556 205861
rect 139792 205625 139876 205861
rect 140112 205625 140196 205861
rect 140432 205625 140516 205861
rect 140752 205625 140836 205861
rect 141072 205625 141156 205861
rect 141392 205625 141476 205861
rect 141712 205625 141796 205861
rect 142032 205625 142116 205861
rect 142352 205625 142436 205861
rect 142672 205625 142756 205861
rect 142992 205625 143076 205861
rect 143312 205625 143396 205861
rect 143632 205625 143716 205861
rect 143952 205625 144036 205861
rect 144272 205625 144356 205861
rect 144592 205625 144676 205861
rect 144912 205625 144996 205861
rect 145232 205625 145316 205861
rect 145552 205625 145636 205861
rect 145872 205625 145956 205861
rect 146192 205625 146276 205861
rect 146512 205625 146596 205861
rect 146832 205625 146916 205861
rect 147152 205625 147236 205861
rect 147472 205625 147556 205861
rect 147792 205625 147876 205861
rect 148112 205625 148196 205861
rect 148432 205625 148516 205861
rect 148752 205625 148836 205861
rect 149072 205625 149156 205861
rect 149392 205625 149476 205861
rect 149712 205625 149796 205861
rect 150032 205625 150116 205861
rect 150352 205625 150436 205861
rect 150672 205625 150756 205861
rect 150992 205625 151076 205861
rect 151312 205625 151396 205861
rect 151632 205625 151716 205861
rect 151952 205625 152036 205861
rect 152272 205625 152356 205861
rect 152592 205625 152676 205861
rect 152912 205625 152996 205861
rect 153232 205625 153316 205861
rect 153552 205625 153636 205861
rect 153872 205625 153956 205861
rect 154192 205625 154276 205861
rect 154512 205625 154596 205861
rect 154832 205625 154916 205861
rect 155152 205625 155236 205861
rect 155472 205625 155556 205861
rect 155792 205625 155876 205861
rect 156112 205625 156196 205861
rect 156432 205625 156516 205861
rect 156752 205625 156836 205861
rect 157072 205625 157156 205861
rect 157392 205625 157476 205861
rect 157712 205625 157796 205861
rect 158032 205625 158116 205861
rect 158352 205625 158436 205861
rect 158672 205625 158756 205861
rect 158992 205625 159076 205861
rect 159312 205625 159396 205861
rect 159632 205625 159716 205861
rect 159952 205625 160036 205861
rect 160272 205625 160356 205861
rect 160592 205625 160676 205861
rect 160912 205625 160996 205861
rect 161232 205625 161316 205861
rect 161552 205625 161636 205861
rect 161872 205625 161956 205861
rect 162192 205625 162276 205861
rect 162512 205625 162596 205861
rect 162832 205625 162916 205861
rect 163152 205625 163236 205861
rect 163472 205625 163556 205861
rect 163792 205625 163876 205861
rect 164112 205625 164196 205861
rect 164432 205625 164516 205861
rect 164752 205625 164836 205861
rect 165072 205625 165156 205861
rect 165392 205625 165514 205861
rect 135914 205500 165514 205625
rect 132294 169954 132914 205398
rect 137314 201411 165514 201486
rect 137314 201175 137376 201411
rect 137612 201175 137696 201411
rect 137932 201175 138016 201411
rect 138252 201175 138336 201411
rect 138572 201175 138656 201411
rect 138892 201175 138976 201411
rect 139212 201175 139296 201411
rect 139532 201175 139616 201411
rect 139852 201175 139936 201411
rect 140172 201175 140256 201411
rect 140492 201175 140576 201411
rect 140812 201175 140896 201411
rect 141132 201175 141216 201411
rect 141452 201175 141536 201411
rect 141772 201175 141856 201411
rect 142092 201175 142176 201411
rect 142412 201175 142496 201411
rect 142732 201175 142816 201411
rect 143052 201175 143136 201411
rect 143372 201175 143456 201411
rect 143692 201175 143776 201411
rect 144012 201175 144096 201411
rect 144332 201175 144416 201411
rect 144652 201175 144736 201411
rect 144972 201175 145056 201411
rect 145292 201175 145376 201411
rect 145612 201175 145696 201411
rect 145932 201175 146016 201411
rect 146252 201175 146336 201411
rect 146572 201175 146656 201411
rect 146892 201175 146976 201411
rect 147212 201175 147296 201411
rect 147532 201175 147616 201411
rect 147852 201175 147936 201411
rect 148172 201175 148256 201411
rect 148492 201175 148576 201411
rect 148812 201175 148896 201411
rect 149132 201175 149216 201411
rect 149452 201175 149536 201411
rect 149772 201175 149856 201411
rect 150092 201175 150176 201411
rect 150412 201175 150496 201411
rect 150732 201175 150816 201411
rect 151052 201175 151136 201411
rect 151372 201175 151456 201411
rect 151692 201175 151776 201411
rect 152012 201175 152096 201411
rect 152332 201175 152416 201411
rect 152652 201175 152736 201411
rect 152972 201175 153056 201411
rect 153292 201175 153376 201411
rect 153612 201175 153696 201411
rect 153932 201175 154016 201411
rect 154252 201175 154336 201411
rect 154572 201175 154656 201411
rect 154892 201175 154976 201411
rect 155212 201175 155296 201411
rect 155532 201175 155616 201411
rect 155852 201175 155936 201411
rect 156172 201175 156256 201411
rect 156492 201175 156576 201411
rect 156812 201175 156896 201411
rect 157132 201175 157216 201411
rect 157452 201175 157536 201411
rect 157772 201175 157856 201411
rect 158092 201175 158176 201411
rect 158412 201175 158496 201411
rect 158732 201175 158816 201411
rect 159052 201175 159136 201411
rect 159372 201175 159456 201411
rect 159692 201175 159776 201411
rect 160012 201175 160096 201411
rect 160332 201175 160416 201411
rect 160652 201175 160736 201411
rect 160972 201175 161056 201411
rect 161292 201175 161376 201411
rect 161612 201175 161696 201411
rect 161932 201175 162016 201411
rect 162252 201175 162336 201411
rect 162572 201175 162656 201411
rect 162892 201175 162976 201411
rect 163212 201175 163296 201411
rect 163532 201175 163616 201411
rect 163852 201175 163936 201411
rect 164172 201175 164256 201411
rect 164492 201175 164576 201411
rect 164812 201175 164896 201411
rect 165132 201175 165216 201411
rect 165452 201175 165514 201411
rect 137314 201100 165514 201175
rect 144867 191044 144933 191045
rect 144867 190980 144868 191044
rect 144932 190980 144933 191044
rect 144867 190979 144933 190980
rect 141003 190364 141069 190365
rect 141003 190300 141004 190364
rect 141068 190300 141069 190364
rect 141003 190299 141069 190300
rect 140819 184244 140885 184245
rect 140819 184180 140820 184244
rect 140884 184180 140885 184244
rect 140819 184179 140885 184180
rect 140822 178669 140882 184179
rect 141006 178805 141066 190299
rect 141739 184380 141805 184381
rect 141739 184316 141740 184380
rect 141804 184316 141805 184380
rect 141739 184315 141805 184316
rect 141742 178805 141802 184315
rect 142843 184108 142909 184109
rect 142843 184044 142844 184108
rect 142908 184044 142909 184108
rect 142843 184043 142909 184044
rect 142475 180980 142541 180981
rect 142475 180916 142476 180980
rect 142540 180916 142541 180980
rect 142475 180915 142541 180916
rect 141003 178804 141069 178805
rect 141003 178740 141004 178804
rect 141068 178740 141069 178804
rect 141003 178739 141069 178740
rect 141739 178804 141805 178805
rect 141739 178740 141740 178804
rect 141804 178740 141805 178804
rect 141739 178739 141805 178740
rect 140819 178668 140885 178669
rect 140819 178604 140820 178668
rect 140884 178604 140885 178668
rect 140819 178603 140885 178604
rect 137014 174454 141514 174486
rect 137014 174218 137066 174454
rect 137302 174218 137386 174454
rect 137622 174218 137706 174454
rect 137942 174218 138026 174454
rect 138262 174218 138346 174454
rect 138582 174218 138666 174454
rect 138902 174218 138986 174454
rect 139222 174218 139306 174454
rect 139542 174218 139626 174454
rect 139862 174218 139946 174454
rect 140182 174218 140266 174454
rect 140502 174218 140586 174454
rect 140822 174218 140906 174454
rect 141142 174218 141226 174454
rect 141462 174218 141514 174454
rect 137014 174134 141514 174218
rect 137014 173898 137066 174134
rect 137302 173898 137386 174134
rect 137622 173898 137706 174134
rect 137942 173898 138026 174134
rect 138262 173898 138346 174134
rect 138582 173898 138666 174134
rect 138902 173898 138986 174134
rect 139222 173898 139306 174134
rect 139542 173898 139626 174134
rect 139862 173898 139946 174134
rect 140182 173898 140266 174134
rect 140502 173898 140586 174134
rect 140822 173898 140906 174134
rect 141142 173898 141226 174134
rect 141462 173898 141514 174134
rect 137014 173866 141514 173898
rect 142478 172957 142538 180915
rect 142846 178941 142906 184043
rect 144870 182205 144930 190979
rect 146155 188596 146221 188597
rect 146155 188532 146156 188596
rect 146220 188532 146221 188596
rect 146155 188531 146221 188532
rect 144867 182204 144933 182205
rect 144867 182140 144868 182204
rect 144932 182140 144933 182204
rect 144867 182139 144933 182140
rect 145051 181252 145117 181253
rect 145051 181188 145052 181252
rect 145116 181188 145117 181252
rect 145051 181187 145117 181188
rect 142843 178940 142909 178941
rect 142843 178876 142844 178940
rect 142908 178876 142909 178940
rect 142843 178875 142909 178876
rect 145054 177445 145114 181187
rect 145051 177444 145117 177445
rect 145051 177380 145052 177444
rect 145116 177380 145117 177444
rect 145051 177379 145117 177380
rect 142475 172956 142541 172957
rect 142475 172892 142476 172956
rect 142540 172892 142541 172956
rect 142475 172891 142541 172892
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 140000 132914 169398
rect 146158 157997 146218 188531
rect 152595 181252 152661 181253
rect 152595 181188 152596 181252
rect 152660 181188 152661 181252
rect 152595 181187 152661 181188
rect 152598 169557 152658 181187
rect 158667 176492 158733 176493
rect 158667 176428 158668 176492
rect 158732 176428 158733 176492
rect 158667 176427 158733 176428
rect 158670 172957 158730 176427
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 158667 172956 158733 172957
rect 158667 172892 158668 172956
rect 158732 172892 158733 172956
rect 158667 172891 158733 172892
rect 152595 169556 152661 169557
rect 152595 169492 152596 169556
rect 152660 169492 152661 169556
rect 152595 169491 152661 169492
rect 146155 157996 146221 157997
rect 146155 157932 146156 157996
rect 146220 157932 146221 157996
rect 146155 157931 146221 157932
rect 172794 140000 173414 173898
rect 177294 214954 177914 228484
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 140000 177914 142398
rect 181794 219454 182414 228484
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 140000 182414 146898
rect 186294 223954 186914 228484
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 139568 115954 139888 115986
rect 139568 115718 139610 115954
rect 139846 115718 139888 115954
rect 139568 115634 139888 115718
rect 139568 115398 139610 115634
rect 139846 115398 139888 115634
rect 139568 115366 139888 115398
rect 170288 115954 170608 115986
rect 170288 115718 170330 115954
rect 170566 115718 170608 115954
rect 170288 115634 170608 115718
rect 170288 115398 170330 115634
rect 170566 115398 170608 115634
rect 170288 115366 170608 115398
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 153515 78572 153581 78573
rect 144870 78510 145298 78570
rect 144870 78029 144930 78510
rect 145238 78029 145298 78510
rect 153515 78508 153516 78572
rect 153580 78508 153581 78572
rect 153515 78507 153581 78508
rect 164003 78572 164069 78573
rect 164003 78508 164004 78572
rect 164068 78508 164069 78572
rect 164003 78507 164069 78508
rect 165291 78572 165357 78573
rect 165291 78508 165292 78572
rect 165356 78508 165357 78572
rect 165291 78507 165357 78508
rect 173571 78572 173637 78573
rect 173571 78508 173572 78572
rect 173636 78508 173637 78572
rect 173571 78507 173637 78508
rect 145419 78164 145485 78165
rect 145419 78100 145420 78164
rect 145484 78100 145485 78164
rect 145419 78099 145485 78100
rect 130699 78028 130765 78029
rect 130699 77964 130700 78028
rect 130764 78026 130765 78028
rect 131067 78028 131133 78029
rect 131067 78026 131068 78028
rect 130764 77966 131068 78026
rect 130764 77964 130765 77966
rect 130699 77963 130765 77964
rect 131067 77964 131068 77966
rect 131132 77964 131133 78028
rect 131067 77963 131133 77964
rect 144867 78028 144933 78029
rect 144867 77964 144868 78028
rect 144932 77964 144933 78028
rect 144867 77963 144933 77964
rect 145235 78028 145301 78029
rect 145235 77964 145236 78028
rect 145300 77964 145301 78028
rect 145235 77963 145301 77964
rect 126651 77892 126717 77893
rect 126651 77828 126652 77892
rect 126716 77828 126717 77892
rect 126651 77827 126717 77828
rect 128675 77892 128741 77893
rect 128675 77828 128676 77892
rect 128740 77828 128741 77892
rect 128675 77827 128741 77828
rect 129595 77892 129661 77893
rect 129595 77828 129596 77892
rect 129660 77890 129661 77892
rect 130515 77892 130581 77893
rect 129660 77830 130210 77890
rect 129660 77828 129661 77830
rect 129595 77827 129661 77828
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 76000
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 76000
rect 125915 75172 125981 75173
rect 125915 75108 125916 75172
rect 125980 75108 125981 75172
rect 125915 75107 125981 75108
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 125918 3365 125978 75107
rect 126654 71365 126714 77827
rect 127203 76804 127269 76805
rect 127203 76740 127204 76804
rect 127268 76740 127269 76804
rect 127203 76739 127269 76740
rect 126651 71364 126717 71365
rect 126651 71300 126652 71364
rect 126716 71300 126717 71364
rect 126651 71299 126717 71300
rect 127206 6629 127266 76739
rect 128678 76397 128738 77827
rect 129043 76804 129109 76805
rect 129043 76740 129044 76804
rect 129108 76740 129109 76804
rect 129043 76739 129109 76740
rect 127387 76396 127453 76397
rect 127387 76332 127388 76396
rect 127452 76332 127453 76396
rect 127387 76331 127453 76332
rect 128675 76396 128741 76397
rect 128675 76332 128676 76396
rect 128740 76332 128741 76396
rect 128675 76331 128741 76332
rect 127203 6628 127269 6629
rect 127203 6564 127204 6628
rect 127268 6564 127269 6628
rect 127203 6563 127269 6564
rect 127390 6221 127450 76331
rect 128491 76124 128557 76125
rect 128491 76060 128492 76124
rect 128556 76060 128557 76124
rect 128491 76059 128557 76060
rect 127794 57454 128414 76000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127387 6220 127453 6221
rect 127387 6156 127388 6220
rect 127452 6156 127453 6220
rect 127387 6155 127453 6156
rect 125915 3364 125981 3365
rect 125915 3300 125916 3364
rect 125980 3300 125981 3364
rect 125915 3299 125981 3300
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 -4186 128414 20898
rect 128494 6930 128554 76059
rect 128859 75852 128925 75853
rect 128859 75788 128860 75852
rect 128924 75788 128925 75852
rect 128859 75787 128925 75788
rect 128675 75580 128741 75581
rect 128675 75516 128676 75580
rect 128740 75516 128741 75580
rect 128675 75515 128741 75516
rect 128678 9077 128738 75515
rect 128675 9076 128741 9077
rect 128675 9012 128676 9076
rect 128740 9012 128741 9076
rect 128675 9011 128741 9012
rect 128862 8941 128922 75787
rect 129046 71093 129106 76739
rect 129779 76396 129845 76397
rect 129779 76332 129780 76396
rect 129844 76332 129845 76396
rect 129779 76331 129845 76332
rect 129963 76396 130029 76397
rect 129963 76332 129964 76396
rect 130028 76332 130029 76396
rect 129963 76331 130029 76332
rect 129782 72589 129842 76331
rect 129779 72588 129845 72589
rect 129779 72524 129780 72588
rect 129844 72524 129845 72588
rect 129779 72523 129845 72524
rect 129043 71092 129109 71093
rect 129043 71028 129044 71092
rect 129108 71028 129109 71092
rect 129043 71027 129109 71028
rect 129966 9213 130026 76331
rect 129963 9212 130029 9213
rect 129963 9148 129964 9212
rect 130028 9148 130029 9212
rect 129963 9147 130029 9148
rect 128859 8940 128925 8941
rect 128859 8876 128860 8940
rect 128924 8876 128925 8940
rect 128859 8875 128925 8876
rect 130150 7581 130210 77830
rect 130515 77828 130516 77892
rect 130580 77828 130581 77892
rect 130515 77827 130581 77828
rect 131435 77892 131501 77893
rect 131435 77828 131436 77892
rect 131500 77828 131501 77892
rect 131435 77827 131501 77828
rect 131987 77892 132053 77893
rect 131987 77828 131988 77892
rect 132052 77828 132053 77892
rect 131987 77827 132053 77828
rect 132539 77892 132605 77893
rect 132539 77828 132540 77892
rect 132604 77828 132605 77892
rect 132539 77827 132605 77828
rect 132907 77892 132973 77893
rect 132907 77828 132908 77892
rect 132972 77828 132973 77892
rect 132907 77827 132973 77828
rect 134195 77892 134261 77893
rect 134195 77828 134196 77892
rect 134260 77828 134261 77892
rect 134195 77827 134261 77828
rect 136035 77892 136101 77893
rect 136035 77828 136036 77892
rect 136100 77828 136101 77892
rect 136035 77827 136101 77828
rect 136403 77892 136469 77893
rect 136403 77828 136404 77892
rect 136468 77828 136469 77892
rect 136403 77827 136469 77828
rect 144683 77892 144749 77893
rect 144683 77828 144684 77892
rect 144748 77890 144749 77892
rect 145235 77892 145301 77893
rect 145235 77890 145236 77892
rect 144748 77830 145236 77890
rect 144748 77828 144749 77830
rect 144683 77827 144749 77828
rect 145235 77828 145236 77830
rect 145300 77828 145301 77892
rect 145235 77827 145301 77828
rect 130518 75445 130578 77827
rect 130699 77756 130765 77757
rect 130699 77692 130700 77756
rect 130764 77692 130765 77756
rect 130699 77691 130765 77692
rect 130702 75717 130762 77691
rect 131438 77485 131498 77827
rect 131990 77485 132050 77827
rect 131435 77484 131501 77485
rect 131435 77420 131436 77484
rect 131500 77420 131501 77484
rect 131435 77419 131501 77420
rect 131987 77484 132053 77485
rect 131987 77420 131988 77484
rect 132052 77420 132053 77484
rect 131987 77419 132053 77420
rect 132542 77213 132602 77827
rect 132539 77212 132605 77213
rect 132539 77148 132540 77212
rect 132604 77148 132605 77212
rect 132539 77147 132605 77148
rect 132910 76397 132970 77827
rect 133091 77756 133157 77757
rect 133091 77692 133092 77756
rect 133156 77692 133157 77756
rect 133091 77691 133157 77692
rect 132907 76396 132973 76397
rect 132907 76332 132908 76396
rect 132972 76332 132973 76396
rect 132907 76331 132973 76332
rect 133094 76261 133154 77691
rect 133091 76260 133157 76261
rect 133091 76196 133092 76260
rect 133156 76196 133157 76260
rect 133091 76195 133157 76196
rect 130699 75716 130765 75717
rect 130699 75652 130700 75716
rect 130764 75652 130765 75716
rect 130699 75651 130765 75652
rect 130515 75444 130581 75445
rect 130515 75380 130516 75444
rect 130580 75380 130581 75444
rect 130515 75379 130581 75380
rect 131435 74900 131501 74901
rect 131435 74836 131436 74900
rect 131500 74836 131501 74900
rect 131435 74835 131501 74836
rect 131067 74764 131133 74765
rect 131067 74700 131068 74764
rect 131132 74700 131133 74764
rect 131067 74699 131133 74700
rect 130147 7580 130213 7581
rect 130147 7516 130148 7580
rect 130212 7516 130213 7580
rect 130147 7515 130213 7516
rect 128494 6870 128738 6930
rect 128678 6357 128738 6870
rect 131070 6493 131130 74699
rect 131251 74628 131317 74629
rect 131251 74564 131252 74628
rect 131316 74564 131317 74628
rect 131251 74563 131317 74564
rect 131254 11661 131314 74563
rect 131438 71909 131498 74835
rect 131435 71908 131501 71909
rect 131435 71844 131436 71908
rect 131500 71844 131501 71908
rect 131435 71843 131501 71844
rect 132294 61954 132914 76000
rect 133091 75036 133157 75037
rect 133091 74972 133092 75036
rect 133156 74972 133157 75036
rect 133091 74971 133157 74972
rect 134011 75036 134077 75037
rect 134011 74972 134012 75036
rect 134076 74972 134077 75036
rect 134011 74971 134077 74972
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 131251 11660 131317 11661
rect 131251 11596 131252 11660
rect 131316 11596 131317 11660
rect 131251 11595 131317 11596
rect 131067 6492 131133 6493
rect 131067 6428 131068 6492
rect 131132 6428 131133 6492
rect 131067 6427 131133 6428
rect 128675 6356 128741 6357
rect 128675 6292 128676 6356
rect 128740 6292 128741 6356
rect 128675 6291 128741 6292
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 -5146 132914 25398
rect 133094 7717 133154 74971
rect 133275 74492 133341 74493
rect 133275 74428 133276 74492
rect 133340 74428 133341 74492
rect 133275 74427 133341 74428
rect 133278 10301 133338 74427
rect 134014 10437 134074 74971
rect 134198 10573 134258 77827
rect 135299 77756 135365 77757
rect 135299 77692 135300 77756
rect 135364 77692 135365 77756
rect 135299 77691 135365 77692
rect 134379 76396 134445 76397
rect 134379 76332 134380 76396
rect 134444 76332 134445 76396
rect 134379 76331 134445 76332
rect 134195 10572 134261 10573
rect 134195 10508 134196 10572
rect 134260 10508 134261 10572
rect 134195 10507 134261 10508
rect 134011 10436 134077 10437
rect 134011 10372 134012 10436
rect 134076 10372 134077 10436
rect 134011 10371 134077 10372
rect 133275 10300 133341 10301
rect 133275 10236 133276 10300
rect 133340 10236 133341 10300
rect 133275 10235 133341 10236
rect 134382 9349 134442 76331
rect 135302 71773 135362 77691
rect 136038 75037 136098 77827
rect 136406 77485 136466 77827
rect 136955 77756 137021 77757
rect 136955 77692 136956 77756
rect 137020 77692 137021 77756
rect 136955 77691 137021 77692
rect 138611 77756 138677 77757
rect 138611 77692 138612 77756
rect 138676 77692 138677 77756
rect 138611 77691 138677 77692
rect 145051 77756 145117 77757
rect 145051 77692 145052 77756
rect 145116 77692 145117 77756
rect 145051 77691 145117 77692
rect 145235 77756 145301 77757
rect 145235 77692 145236 77756
rect 145300 77692 145301 77756
rect 145235 77691 145301 77692
rect 136403 77484 136469 77485
rect 136403 77420 136404 77484
rect 136468 77420 136469 77484
rect 136403 77419 136469 77420
rect 136958 77310 137018 77691
rect 137691 77484 137757 77485
rect 137691 77420 137692 77484
rect 137756 77420 137757 77484
rect 137691 77419 137757 77420
rect 136590 77250 137018 77310
rect 135667 75036 135733 75037
rect 135667 74972 135668 75036
rect 135732 74972 135733 75036
rect 135667 74971 135733 74972
rect 136035 75036 136101 75037
rect 136035 74972 136036 75036
rect 136100 74972 136101 75036
rect 136035 74971 136101 74972
rect 135299 71772 135365 71773
rect 135299 71708 135300 71772
rect 135364 71708 135365 71772
rect 135299 71707 135365 71708
rect 134379 9348 134445 9349
rect 134379 9284 134380 9348
rect 134444 9284 134445 9348
rect 134379 9283 134445 9284
rect 133091 7716 133157 7717
rect 133091 7652 133092 7716
rect 133156 7652 133157 7716
rect 133091 7651 133157 7652
rect 135670 3365 135730 74971
rect 136403 73812 136469 73813
rect 136403 73748 136404 73812
rect 136468 73748 136469 73812
rect 136403 73747 136469 73748
rect 136406 3365 136466 73747
rect 136590 73405 136650 77250
rect 136587 73404 136653 73405
rect 136587 73340 136588 73404
rect 136652 73340 136653 73404
rect 136587 73339 136653 73340
rect 136794 66454 137414 76000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 135667 3364 135733 3365
rect 135667 3300 135668 3364
rect 135732 3300 135733 3364
rect 135667 3299 135733 3300
rect 136403 3364 136469 3365
rect 136403 3300 136404 3364
rect 136468 3300 136469 3364
rect 136403 3299 136469 3300
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 -6106 137414 29898
rect 137694 16421 137754 77419
rect 137875 75036 137941 75037
rect 137875 74972 137876 75036
rect 137940 74972 137941 75036
rect 137875 74971 137941 74972
rect 137691 16420 137757 16421
rect 137691 16356 137692 16420
rect 137756 16356 137757 16420
rect 137691 16355 137757 16356
rect 137878 4861 137938 74971
rect 138614 73949 138674 77691
rect 140635 77620 140701 77621
rect 140635 77556 140636 77620
rect 140700 77556 140701 77620
rect 140635 77555 140701 77556
rect 144867 77620 144933 77621
rect 144867 77556 144868 77620
rect 144932 77556 144933 77620
rect 144867 77555 144933 77556
rect 138979 76396 139045 76397
rect 138979 76332 138980 76396
rect 139044 76332 139045 76396
rect 138979 76331 139045 76332
rect 139163 76396 139229 76397
rect 139163 76332 139164 76396
rect 139228 76332 139229 76396
rect 139163 76331 139229 76332
rect 138795 75036 138861 75037
rect 138795 74972 138796 75036
rect 138860 74972 138861 75036
rect 138795 74971 138861 74972
rect 138611 73948 138677 73949
rect 138611 73884 138612 73948
rect 138676 73884 138677 73948
rect 138611 73883 138677 73884
rect 138798 65517 138858 74971
rect 138795 65516 138861 65517
rect 138795 65452 138796 65516
rect 138860 65452 138861 65516
rect 138795 65451 138861 65452
rect 138982 63069 139042 76331
rect 138979 63068 139045 63069
rect 138979 63004 138980 63068
rect 139044 63004 139045 63068
rect 138979 63003 139045 63004
rect 139166 33965 139226 76331
rect 140083 75036 140149 75037
rect 140083 74972 140084 75036
rect 140148 74972 140149 75036
rect 140083 74971 140149 74972
rect 140451 75036 140517 75037
rect 140451 74972 140452 75036
rect 140516 74972 140517 75036
rect 140451 74971 140517 74972
rect 140086 62933 140146 74971
rect 140267 74900 140333 74901
rect 140267 74836 140268 74900
rect 140332 74836 140333 74900
rect 140267 74835 140333 74836
rect 140083 62932 140149 62933
rect 140083 62868 140084 62932
rect 140148 62868 140149 62932
rect 140083 62867 140149 62868
rect 140270 57357 140330 74835
rect 140267 57356 140333 57357
rect 140267 57292 140268 57356
rect 140332 57292 140333 57356
rect 140267 57291 140333 57292
rect 139163 33964 139229 33965
rect 139163 33900 139164 33964
rect 139228 33900 139229 33964
rect 139163 33899 139229 33900
rect 140454 27029 140514 74971
rect 140451 27028 140517 27029
rect 140451 26964 140452 27028
rect 140516 26964 140517 27028
rect 140451 26963 140517 26964
rect 140638 18733 140698 77555
rect 144870 77485 144930 77555
rect 144867 77484 144933 77485
rect 144867 77420 144868 77484
rect 144932 77420 144933 77484
rect 144867 77419 144933 77420
rect 145054 77310 145114 77691
rect 144870 77250 145114 77310
rect 141003 74628 141069 74629
rect 141003 74564 141004 74628
rect 141068 74564 141069 74628
rect 141003 74563 141069 74564
rect 140635 18732 140701 18733
rect 140635 18668 140636 18732
rect 140700 18668 140701 18732
rect 140635 18667 140701 18668
rect 141006 12205 141066 74563
rect 141294 70954 141914 76000
rect 144131 75172 144197 75173
rect 144131 75108 144132 75172
rect 144196 75108 144197 75172
rect 144131 75107 144197 75108
rect 142843 74900 142909 74901
rect 142843 74836 142844 74900
rect 142908 74836 142909 74900
rect 142843 74835 142909 74836
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141003 12204 141069 12205
rect 141003 12140 141004 12204
rect 141068 12140 141069 12204
rect 141003 12139 141069 12140
rect 137875 4860 137941 4861
rect 137875 4796 137876 4860
rect 137940 4796 137941 4860
rect 137875 4795 137941 4796
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 -7066 141914 34398
rect 142846 6221 142906 74835
rect 143027 74764 143093 74765
rect 143027 74700 143028 74764
rect 143092 74700 143093 74764
rect 143027 74699 143093 74700
rect 143395 74764 143461 74765
rect 143395 74700 143396 74764
rect 143460 74700 143461 74764
rect 143395 74699 143461 74700
rect 143030 33829 143090 74699
rect 143211 74628 143277 74629
rect 143211 74564 143212 74628
rect 143276 74564 143277 74628
rect 143211 74563 143277 74564
rect 143027 33828 143093 33829
rect 143027 33764 143028 33828
rect 143092 33764 143093 33828
rect 143027 33763 143093 33764
rect 143214 28253 143274 74563
rect 143398 71501 143458 74699
rect 143395 71500 143461 71501
rect 143395 71436 143396 71500
rect 143460 71436 143461 71500
rect 143395 71435 143461 71436
rect 143211 28252 143277 28253
rect 143211 28188 143212 28252
rect 143276 28188 143277 28252
rect 143211 28187 143277 28188
rect 144134 20093 144194 75107
rect 144499 75036 144565 75037
rect 144499 74972 144500 75036
rect 144564 74972 144565 75036
rect 144499 74971 144565 74972
rect 144502 57221 144562 74971
rect 144870 71365 144930 77250
rect 145238 75037 145298 77691
rect 145422 77485 145482 78099
rect 151491 77892 151557 77893
rect 151491 77828 151492 77892
rect 151556 77828 151557 77892
rect 151491 77827 151557 77828
rect 152043 77892 152109 77893
rect 152043 77828 152044 77892
rect 152108 77828 152109 77892
rect 152043 77827 152109 77828
rect 152779 77892 152845 77893
rect 152779 77828 152780 77892
rect 152844 77828 152845 77892
rect 153377 77892 153443 77893
rect 153377 77890 153378 77892
rect 152779 77827 152845 77828
rect 153334 77828 153378 77890
rect 153442 77828 153443 77892
rect 153334 77827 153443 77828
rect 145419 77484 145485 77485
rect 145419 77420 145420 77484
rect 145484 77420 145485 77484
rect 145419 77419 145485 77420
rect 147259 76804 147325 76805
rect 147259 76740 147260 76804
rect 147324 76740 147325 76804
rect 147259 76739 147325 76740
rect 145603 76396 145669 76397
rect 145603 76332 145604 76396
rect 145668 76332 145669 76396
rect 145603 76331 145669 76332
rect 145419 76260 145485 76261
rect 145419 76196 145420 76260
rect 145484 76196 145485 76260
rect 145419 76195 145485 76196
rect 145235 75036 145301 75037
rect 145235 74972 145236 75036
rect 145300 74972 145301 75036
rect 145235 74971 145301 74972
rect 144867 71364 144933 71365
rect 144867 71300 144868 71364
rect 144932 71300 144933 71364
rect 144867 71299 144933 71300
rect 144499 57220 144565 57221
rect 144499 57156 144500 57220
rect 144564 57156 144565 57220
rect 144499 57155 144565 57156
rect 144131 20092 144197 20093
rect 144131 20028 144132 20092
rect 144196 20028 144197 20092
rect 144131 20027 144197 20028
rect 145422 8125 145482 76195
rect 145419 8124 145485 8125
rect 145419 8060 145420 8124
rect 145484 8060 145485 8124
rect 145419 8059 145485 8060
rect 145606 7989 145666 76331
rect 145794 75454 146414 76000
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 147075 73540 147141 73541
rect 147075 73476 147076 73540
rect 147140 73476 147141 73540
rect 147075 73475 147141 73476
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145603 7988 145669 7989
rect 145603 7924 145604 7988
rect 145668 7924 145669 7988
rect 145603 7923 145669 7924
rect 142843 6220 142909 6221
rect 142843 6156 142844 6220
rect 142908 6156 142909 6220
rect 142843 6155 142909 6156
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 3454 146414 38898
rect 147078 9349 147138 73475
rect 147262 35325 147322 76739
rect 149835 76260 149901 76261
rect 149835 76196 149836 76260
rect 149900 76196 149901 76260
rect 149835 76195 149901 76196
rect 148915 75716 148981 75717
rect 148915 75652 148916 75716
rect 148980 75652 148981 75716
rect 148915 75651 148981 75652
rect 149651 75716 149717 75717
rect 149651 75652 149652 75716
rect 149716 75652 149717 75716
rect 149651 75651 149717 75652
rect 148731 75036 148797 75037
rect 148731 74972 148732 75036
rect 148796 74972 148797 75036
rect 148731 74971 148797 74972
rect 148547 74628 148613 74629
rect 148547 74564 148548 74628
rect 148612 74564 148613 74628
rect 148547 74563 148613 74564
rect 147259 35324 147325 35325
rect 147259 35260 147260 35324
rect 147324 35260 147325 35324
rect 147259 35259 147325 35260
rect 148550 19957 148610 74563
rect 148547 19956 148613 19957
rect 148547 19892 148548 19956
rect 148612 19892 148613 19956
rect 148547 19891 148613 19892
rect 147075 9348 147141 9349
rect 147075 9284 147076 9348
rect 147140 9284 147141 9348
rect 147075 9283 147141 9284
rect 148734 9077 148794 74971
rect 148918 9213 148978 75651
rect 149654 25533 149714 75651
rect 149838 35189 149898 76195
rect 150294 43954 150914 76000
rect 151307 75716 151373 75717
rect 151307 75652 151308 75716
rect 151372 75652 151373 75716
rect 151307 75651 151373 75652
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 149835 35188 149901 35189
rect 149835 35124 149836 35188
rect 149900 35124 149901 35188
rect 149835 35123 149901 35124
rect 149651 25532 149717 25533
rect 149651 25468 149652 25532
rect 149716 25468 149717 25532
rect 149651 25467 149717 25468
rect 148915 9212 148981 9213
rect 148915 9148 148916 9212
rect 148980 9148 148981 9212
rect 148915 9147 148981 9148
rect 148731 9076 148797 9077
rect 148731 9012 148732 9076
rect 148796 9012 148797 9076
rect 148731 9011 148797 9012
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 7954 150914 43398
rect 151310 10437 151370 75651
rect 151307 10436 151373 10437
rect 151307 10372 151308 10436
rect 151372 10372 151373 10436
rect 151307 10371 151373 10372
rect 151494 10301 151554 77827
rect 152046 75037 152106 77827
rect 152411 77756 152477 77757
rect 152411 77692 152412 77756
rect 152476 77692 152477 77756
rect 152411 77691 152477 77692
rect 152414 75989 152474 77691
rect 152595 76124 152661 76125
rect 152595 76060 152596 76124
rect 152660 76060 152661 76124
rect 152595 76059 152661 76060
rect 152411 75988 152477 75989
rect 152411 75924 152412 75988
rect 152476 75924 152477 75988
rect 152411 75923 152477 75924
rect 152411 75716 152477 75717
rect 152411 75652 152412 75716
rect 152476 75652 152477 75716
rect 152411 75651 152477 75652
rect 152043 75036 152109 75037
rect 152043 74972 152044 75036
rect 152108 74972 152109 75036
rect 152043 74971 152109 74972
rect 151675 72860 151741 72861
rect 151675 72796 151676 72860
rect 151740 72796 151741 72860
rect 151675 72795 151741 72796
rect 151491 10300 151557 10301
rect 151491 10236 151492 10300
rect 151556 10236 151557 10300
rect 151491 10235 151557 10236
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 151678 7853 151738 72795
rect 152414 12069 152474 75651
rect 152598 17373 152658 76059
rect 152595 17372 152661 17373
rect 152595 17308 152596 17372
rect 152660 17308 152661 17372
rect 152595 17307 152661 17308
rect 152782 14925 152842 77827
rect 153147 77620 153213 77621
rect 153147 77556 153148 77620
rect 153212 77556 153213 77620
rect 153147 77555 153213 77556
rect 153150 71790 153210 77555
rect 153334 76805 153394 77827
rect 153518 77213 153578 78507
rect 162163 78436 162229 78437
rect 162163 78372 162164 78436
rect 162228 78372 162229 78436
rect 162163 78371 162229 78372
rect 155171 78300 155237 78301
rect 155171 78236 155172 78300
rect 155236 78236 155237 78300
rect 155171 78235 155237 78236
rect 155174 78029 155234 78235
rect 155171 78028 155237 78029
rect 155171 77964 155172 78028
rect 155236 77964 155237 78028
rect 155171 77963 155237 77964
rect 162166 77893 162226 78371
rect 164006 78301 164066 78507
rect 163819 78300 163885 78301
rect 163819 78236 163820 78300
rect 163884 78236 163885 78300
rect 163819 78235 163885 78236
rect 164003 78300 164069 78301
rect 164003 78236 164004 78300
rect 164068 78236 164069 78300
rect 164003 78235 164069 78236
rect 153699 77892 153765 77893
rect 153699 77828 153700 77892
rect 153764 77890 153765 77892
rect 154067 77892 154133 77893
rect 153764 77830 153946 77890
rect 153764 77828 153765 77830
rect 153699 77827 153765 77828
rect 153886 77213 153946 77830
rect 154067 77828 154068 77892
rect 154132 77828 154133 77892
rect 154067 77827 154133 77828
rect 154251 77892 154317 77893
rect 154251 77828 154252 77892
rect 154316 77828 154317 77892
rect 154251 77827 154317 77828
rect 154987 77892 155053 77893
rect 154987 77828 154988 77892
rect 155052 77828 155053 77892
rect 154987 77827 155053 77828
rect 156827 77892 156893 77893
rect 156827 77828 156828 77892
rect 156892 77828 156893 77892
rect 156827 77827 156893 77828
rect 158115 77892 158181 77893
rect 158115 77828 158116 77892
rect 158180 77828 158181 77892
rect 158115 77827 158181 77828
rect 158667 77892 158733 77893
rect 158667 77828 158668 77892
rect 158732 77828 158733 77892
rect 158667 77827 158733 77828
rect 162163 77892 162229 77893
rect 162163 77828 162164 77892
rect 162228 77828 162229 77892
rect 162715 77892 162781 77893
rect 162715 77890 162716 77892
rect 162163 77827 162229 77828
rect 162350 77830 162716 77890
rect 153515 77212 153581 77213
rect 153515 77148 153516 77212
rect 153580 77148 153581 77212
rect 153515 77147 153581 77148
rect 153883 77212 153949 77213
rect 153883 77148 153884 77212
rect 153948 77148 153949 77212
rect 153883 77147 153949 77148
rect 153331 76804 153397 76805
rect 153331 76740 153332 76804
rect 153396 76740 153397 76804
rect 153331 76739 153397 76740
rect 153331 76396 153397 76397
rect 153331 76332 153332 76396
rect 153396 76332 153397 76396
rect 153331 76331 153397 76332
rect 153334 75309 153394 76331
rect 154070 76261 154130 77827
rect 154254 77621 154314 77827
rect 154251 77620 154317 77621
rect 154251 77556 154252 77620
rect 154316 77556 154317 77620
rect 154251 77555 154317 77556
rect 154990 77077 155050 77827
rect 156091 77756 156157 77757
rect 156091 77692 156092 77756
rect 156156 77692 156157 77756
rect 156091 77691 156157 77692
rect 156643 77756 156709 77757
rect 156643 77692 156644 77756
rect 156708 77692 156709 77756
rect 156643 77691 156709 77692
rect 156094 77077 156154 77691
rect 156275 77620 156341 77621
rect 156275 77556 156276 77620
rect 156340 77556 156341 77620
rect 156275 77555 156341 77556
rect 154987 77076 155053 77077
rect 154987 77012 154988 77076
rect 155052 77012 155053 77076
rect 154987 77011 155053 77012
rect 156091 77076 156157 77077
rect 156091 77012 156092 77076
rect 156156 77012 156157 77076
rect 156091 77011 156157 77012
rect 154435 76804 154501 76805
rect 154435 76740 154436 76804
rect 154500 76740 154501 76804
rect 154435 76739 154501 76740
rect 155723 76804 155789 76805
rect 155723 76740 155724 76804
rect 155788 76740 155789 76804
rect 155723 76739 155789 76740
rect 154067 76260 154133 76261
rect 154067 76196 154068 76260
rect 154132 76196 154133 76260
rect 154067 76195 154133 76196
rect 153883 75852 153949 75853
rect 153883 75788 153884 75852
rect 153948 75788 153949 75852
rect 153883 75787 153949 75788
rect 153331 75308 153397 75309
rect 153331 75244 153332 75308
rect 153396 75244 153397 75308
rect 153331 75243 153397 75244
rect 152966 71730 153210 71790
rect 152966 66877 153026 71730
rect 152963 66876 153029 66877
rect 152963 66812 152964 66876
rect 153028 66812 153029 66876
rect 152963 66811 153029 66812
rect 152779 14924 152845 14925
rect 152779 14860 152780 14924
rect 152844 14860 152845 14924
rect 152779 14859 152845 14860
rect 152411 12068 152477 12069
rect 152411 12004 152412 12068
rect 152476 12004 152477 12068
rect 152411 12003 152477 12004
rect 153886 11933 153946 75787
rect 154251 75716 154317 75717
rect 154251 75652 154252 75716
rect 154316 75652 154317 75716
rect 154251 75651 154317 75652
rect 154067 75580 154133 75581
rect 154067 75516 154068 75580
rect 154132 75516 154133 75580
rect 154067 75515 154133 75516
rect 154070 16285 154130 75515
rect 154067 16284 154133 16285
rect 154067 16220 154068 16284
rect 154132 16220 154133 16284
rect 154067 16219 154133 16220
rect 154254 13021 154314 75651
rect 154438 68237 154498 76739
rect 154435 68236 154501 68237
rect 154435 68172 154436 68236
rect 154500 68172 154501 68236
rect 154435 68171 154501 68172
rect 154794 48454 155414 76000
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154251 13020 154317 13021
rect 154251 12956 154252 13020
rect 154316 12956 154317 13020
rect 154251 12955 154317 12956
rect 154794 12454 155414 47898
rect 155726 14789 155786 76739
rect 156278 75717 156338 77555
rect 156275 75716 156341 75717
rect 156275 75652 156276 75716
rect 156340 75652 156341 75716
rect 156275 75651 156341 75652
rect 155723 14788 155789 14789
rect 155723 14724 155724 14788
rect 155788 14724 155789 14788
rect 155723 14723 155789 14724
rect 156646 14653 156706 77691
rect 156830 54501 156890 77827
rect 157931 76124 157997 76125
rect 157931 76060 157932 76124
rect 157996 76060 157997 76124
rect 157931 76059 157997 76060
rect 157011 75716 157077 75717
rect 157011 75652 157012 75716
rect 157076 75652 157077 75716
rect 157011 75651 157077 75652
rect 156827 54500 156893 54501
rect 156827 54436 156828 54500
rect 156892 54436 156893 54500
rect 156827 54435 156893 54436
rect 157014 16149 157074 75651
rect 157934 36549 157994 76059
rect 157931 36548 157997 36549
rect 157931 36484 157932 36548
rect 157996 36484 157997 36548
rect 157931 36483 157997 36484
rect 157011 16148 157077 16149
rect 157011 16084 157012 16148
rect 157076 16084 157077 16148
rect 157011 16083 157077 16084
rect 158118 15877 158178 77827
rect 158483 77756 158549 77757
rect 158483 77692 158484 77756
rect 158548 77692 158549 77756
rect 158483 77691 158549 77692
rect 158299 77620 158365 77621
rect 158299 77556 158300 77620
rect 158364 77556 158365 77620
rect 158299 77555 158365 77556
rect 158302 16013 158362 77555
rect 158299 16012 158365 16013
rect 158299 15948 158300 16012
rect 158364 15948 158365 16012
rect 158299 15947 158365 15948
rect 158115 15876 158181 15877
rect 158115 15812 158116 15876
rect 158180 15812 158181 15876
rect 158115 15811 158181 15812
rect 156643 14652 156709 14653
rect 156643 14588 156644 14652
rect 156708 14588 156709 14652
rect 156643 14587 156709 14588
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 153883 11932 153949 11933
rect 153883 11868 153884 11932
rect 153948 11868 153949 11932
rect 153883 11867 153949 11868
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 151675 7852 151741 7853
rect 151675 7788 151676 7852
rect 151740 7788 151741 7852
rect 151675 7787 151741 7788
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 -2266 155414 11898
rect 158486 7717 158546 77691
rect 158670 75717 158730 77827
rect 160323 77756 160389 77757
rect 160323 77692 160324 77756
rect 160388 77692 160389 77756
rect 160691 77756 160757 77757
rect 160691 77754 160692 77756
rect 160323 77691 160389 77692
rect 160510 77694 160692 77754
rect 158667 75716 158733 75717
rect 158667 75652 158668 75716
rect 158732 75652 158733 75716
rect 158667 75651 158733 75652
rect 159035 75172 159101 75173
rect 159035 75108 159036 75172
rect 159100 75108 159101 75172
rect 159035 75107 159101 75108
rect 158851 75036 158917 75037
rect 158851 74972 158852 75036
rect 158916 74972 158917 75036
rect 158851 74971 158917 74972
rect 158854 59941 158914 74971
rect 158851 59940 158917 59941
rect 158851 59876 158852 59940
rect 158916 59876 158917 59940
rect 158851 59875 158917 59876
rect 159038 21453 159098 75107
rect 159294 52954 159914 76000
rect 160326 73133 160386 77691
rect 160510 74493 160570 77694
rect 160691 77692 160692 77694
rect 160756 77692 160757 77756
rect 160691 77691 160757 77692
rect 161243 77756 161309 77757
rect 161243 77692 161244 77756
rect 161308 77692 161309 77756
rect 161243 77691 161309 77692
rect 160691 75988 160757 75989
rect 160691 75924 160692 75988
rect 160756 75924 160757 75988
rect 160691 75923 160757 75924
rect 160507 74492 160573 74493
rect 160507 74428 160508 74492
rect 160572 74428 160573 74492
rect 160507 74427 160573 74428
rect 160323 73132 160389 73133
rect 160323 73068 160324 73132
rect 160388 73068 160389 73132
rect 160323 73067 160389 73068
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159035 21452 159101 21453
rect 159035 21388 159036 21452
rect 159100 21388 159101 21452
rect 159035 21387 159101 21388
rect 159294 16954 159914 52398
rect 160694 30973 160754 75923
rect 160875 75580 160941 75581
rect 160875 75516 160876 75580
rect 160940 75516 160941 75580
rect 160875 75515 160941 75516
rect 161059 75580 161125 75581
rect 161059 75516 161060 75580
rect 161124 75516 161125 75580
rect 161059 75515 161125 75516
rect 160691 30972 160757 30973
rect 160691 30908 160692 30972
rect 160756 30908 160757 30972
rect 160691 30907 160757 30908
rect 160878 18597 160938 75515
rect 160875 18596 160941 18597
rect 160875 18532 160876 18596
rect 160940 18532 160941 18596
rect 160875 18531 160941 18532
rect 161062 17237 161122 75515
rect 161059 17236 161125 17237
rect 161059 17172 161060 17236
rect 161124 17172 161125 17236
rect 161059 17171 161125 17172
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 158483 7716 158549 7717
rect 158483 7652 158484 7716
rect 158548 7652 158549 7716
rect 158483 7651 158549 7652
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 -3226 159914 16398
rect 161246 11797 161306 77691
rect 162350 76394 162410 77830
rect 162715 77828 162716 77830
rect 162780 77828 162781 77892
rect 162715 77827 162781 77828
rect 163083 77892 163149 77893
rect 163083 77828 163084 77892
rect 163148 77828 163149 77892
rect 163083 77827 163149 77828
rect 163267 77892 163333 77893
rect 163267 77828 163268 77892
rect 163332 77828 163333 77892
rect 163267 77827 163333 77828
rect 163635 77892 163701 77893
rect 163635 77828 163636 77892
rect 163700 77828 163701 77892
rect 163635 77827 163701 77828
rect 162715 77756 162781 77757
rect 162715 77692 162716 77756
rect 162780 77692 162781 77756
rect 162715 77691 162781 77692
rect 162166 76334 162410 76394
rect 162531 76396 162597 76397
rect 161243 11796 161309 11797
rect 161243 11732 161244 11796
rect 161308 11732 161309 11796
rect 161243 11731 161309 11732
rect 162166 7581 162226 76334
rect 162531 76332 162532 76396
rect 162596 76332 162597 76396
rect 162531 76331 162597 76332
rect 162347 76260 162413 76261
rect 162347 76196 162348 76260
rect 162412 76196 162413 76260
rect 162347 76195 162413 76196
rect 162350 39269 162410 76195
rect 162347 39268 162413 39269
rect 162347 39204 162348 39268
rect 162412 39204 162413 39268
rect 162347 39203 162413 39204
rect 162534 29613 162594 76331
rect 162718 70005 162778 77691
rect 163086 75989 163146 77827
rect 163083 75988 163149 75989
rect 163083 75924 163084 75988
rect 163148 75924 163149 75988
rect 163083 75923 163149 75924
rect 163270 75581 163330 77827
rect 163451 76260 163517 76261
rect 163451 76196 163452 76260
rect 163516 76196 163517 76260
rect 163451 76195 163517 76196
rect 163267 75580 163333 75581
rect 163267 75516 163268 75580
rect 163332 75516 163333 75580
rect 163267 75515 163333 75516
rect 162715 70004 162781 70005
rect 162715 69940 162716 70004
rect 162780 69940 162781 70004
rect 162715 69939 162781 69940
rect 162531 29612 162597 29613
rect 162531 29548 162532 29612
rect 162596 29548 162597 29612
rect 162531 29547 162597 29548
rect 163454 14517 163514 76195
rect 163451 14516 163517 14517
rect 163451 14452 163452 14516
rect 163516 14452 163517 14516
rect 163451 14451 163517 14452
rect 162163 7580 162229 7581
rect 162163 7516 162164 7580
rect 162228 7516 162229 7580
rect 162163 7515 162229 7516
rect 163638 3501 163698 77827
rect 163822 77757 163882 78235
rect 164371 77892 164437 77893
rect 164371 77828 164372 77892
rect 164436 77828 164437 77892
rect 164923 77892 164989 77893
rect 164923 77890 164924 77892
rect 164371 77827 164437 77828
rect 164742 77830 164924 77890
rect 163819 77756 163885 77757
rect 163819 77692 163820 77756
rect 163884 77692 163885 77756
rect 163819 77691 163885 77692
rect 164374 77485 164434 77827
rect 164555 77620 164621 77621
rect 164555 77556 164556 77620
rect 164620 77556 164621 77620
rect 164555 77555 164621 77556
rect 164371 77484 164437 77485
rect 164371 77420 164372 77484
rect 164436 77420 164437 77484
rect 164371 77419 164437 77420
rect 163794 57454 164414 76000
rect 164558 75309 164618 77555
rect 164555 75308 164621 75309
rect 164555 75244 164556 75308
rect 164620 75244 164621 75308
rect 164555 75243 164621 75244
rect 164742 75173 164802 77830
rect 164923 77828 164924 77830
rect 164988 77828 164989 77892
rect 164923 77827 164989 77828
rect 165107 77892 165173 77893
rect 165107 77828 165108 77892
rect 165172 77828 165173 77892
rect 165107 77827 165173 77828
rect 164923 77076 164989 77077
rect 164923 77012 164924 77076
rect 164988 77012 164989 77076
rect 164923 77011 164989 77012
rect 164739 75172 164805 75173
rect 164739 75108 164740 75172
rect 164804 75108 164805 75172
rect 164739 75107 164805 75108
rect 164926 70413 164986 77011
rect 164923 70412 164989 70413
rect 164923 70348 164924 70412
rect 164988 70348 164989 70412
rect 164923 70347 164989 70348
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163635 3500 163701 3501
rect 163635 3436 163636 3500
rect 163700 3436 163701 3500
rect 163635 3435 163701 3436
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 -4186 164414 20898
rect 165110 8941 165170 77827
rect 165294 77485 165354 78507
rect 171363 78436 171429 78437
rect 171363 78372 171364 78436
rect 171428 78372 171429 78436
rect 171363 78371 171429 78372
rect 171547 78436 171613 78437
rect 171547 78372 171548 78436
rect 171612 78372 171613 78436
rect 171547 78371 171613 78372
rect 169339 78164 169405 78165
rect 169339 78100 169340 78164
rect 169404 78100 169405 78164
rect 169339 78099 169405 78100
rect 167315 78028 167381 78029
rect 167315 77964 167316 78028
rect 167380 77964 167381 78028
rect 167315 77963 167381 77964
rect 167683 78028 167749 78029
rect 167683 77964 167684 78028
rect 167748 77964 167749 78028
rect 167683 77963 167749 77964
rect 165475 77892 165541 77893
rect 165475 77828 165476 77892
rect 165540 77828 165541 77892
rect 165475 77827 165541 77828
rect 165843 77892 165909 77893
rect 165843 77828 165844 77892
rect 165908 77828 165909 77892
rect 165843 77827 165909 77828
rect 166763 77892 166829 77893
rect 166763 77828 166764 77892
rect 166828 77828 166829 77892
rect 166763 77827 166829 77828
rect 165291 77484 165357 77485
rect 165291 77420 165292 77484
rect 165356 77420 165357 77484
rect 165291 77419 165357 77420
rect 165478 73170 165538 77827
rect 165294 73110 165538 73170
rect 165294 21317 165354 73110
rect 165846 70957 165906 77827
rect 166027 77620 166093 77621
rect 166027 77556 166028 77620
rect 166092 77556 166093 77620
rect 166027 77555 166093 77556
rect 166579 77620 166645 77621
rect 166579 77556 166580 77620
rect 166644 77556 166645 77620
rect 166579 77555 166645 77556
rect 166030 73541 166090 77555
rect 166395 77076 166461 77077
rect 166395 77012 166396 77076
rect 166460 77012 166461 77076
rect 166395 77011 166461 77012
rect 166211 76260 166277 76261
rect 166211 76196 166212 76260
rect 166276 76196 166277 76260
rect 166211 76195 166277 76196
rect 166027 73540 166093 73541
rect 166027 73476 166028 73540
rect 166092 73476 166093 73540
rect 166027 73475 166093 73476
rect 165843 70956 165909 70957
rect 165843 70892 165844 70956
rect 165908 70892 165909 70956
rect 165843 70891 165909 70892
rect 166214 62797 166274 76195
rect 166211 62796 166277 62797
rect 166211 62732 166212 62796
rect 166276 62732 166277 62796
rect 166211 62731 166277 62732
rect 166398 32741 166458 77011
rect 166395 32740 166461 32741
rect 166395 32676 166396 32740
rect 166460 32676 166461 32740
rect 166395 32675 166461 32676
rect 166582 22677 166642 77555
rect 166579 22676 166645 22677
rect 166579 22612 166580 22676
rect 166644 22612 166645 22676
rect 166579 22611 166645 22612
rect 165291 21316 165357 21317
rect 165291 21252 165292 21316
rect 165356 21252 165357 21316
rect 165291 21251 165357 21252
rect 165107 8940 165173 8941
rect 165107 8876 165108 8940
rect 165172 8876 165173 8940
rect 165107 8875 165173 8876
rect 166766 4997 166826 77827
rect 167318 74765 167378 77963
rect 167499 77892 167565 77893
rect 167499 77828 167500 77892
rect 167564 77828 167565 77892
rect 167499 77827 167565 77828
rect 167502 76805 167562 77827
rect 167499 76804 167565 76805
rect 167499 76740 167500 76804
rect 167564 76740 167565 76804
rect 167499 76739 167565 76740
rect 167499 76396 167565 76397
rect 167499 76332 167500 76396
rect 167564 76332 167565 76396
rect 167499 76331 167565 76332
rect 167315 74764 167381 74765
rect 167315 74700 167316 74764
rect 167380 74700 167381 74764
rect 167315 74699 167381 74700
rect 167502 32469 167562 76331
rect 167686 32605 167746 77963
rect 168603 77892 168669 77893
rect 168603 77828 168604 77892
rect 168668 77828 168669 77892
rect 168603 77827 168669 77828
rect 168051 76804 168117 76805
rect 168051 76740 168052 76804
rect 168116 76740 168117 76804
rect 168051 76739 168117 76740
rect 167867 75852 167933 75853
rect 167867 75788 167868 75852
rect 167932 75788 167933 75852
rect 167867 75787 167933 75788
rect 167683 32604 167749 32605
rect 167683 32540 167684 32604
rect 167748 32540 167749 32604
rect 167683 32539 167749 32540
rect 167499 32468 167565 32469
rect 167499 32404 167500 32468
rect 167564 32404 167565 32468
rect 167499 32403 167565 32404
rect 167870 24309 167930 75787
rect 167867 24308 167933 24309
rect 167867 24244 167868 24308
rect 167932 24244 167933 24308
rect 167867 24243 167933 24244
rect 166763 4996 166829 4997
rect 166763 4932 166764 4996
rect 166828 4932 166829 4996
rect 166763 4931 166829 4932
rect 168054 4861 168114 76739
rect 168606 76397 168666 77827
rect 169342 77485 169402 78099
rect 170075 77892 170141 77893
rect 170075 77828 170076 77892
rect 170140 77828 170141 77892
rect 170075 77827 170141 77828
rect 170259 77892 170325 77893
rect 170259 77828 170260 77892
rect 170324 77828 170325 77892
rect 170259 77827 170325 77828
rect 170627 77892 170693 77893
rect 170627 77828 170628 77892
rect 170692 77828 170693 77892
rect 170627 77827 170693 77828
rect 170995 77892 171061 77893
rect 170995 77828 170996 77892
rect 171060 77828 171061 77892
rect 170995 77827 171061 77828
rect 169339 77484 169405 77485
rect 169339 77420 169340 77484
rect 169404 77420 169405 77484
rect 169339 77419 169405 77420
rect 168603 76396 168669 76397
rect 168603 76332 168604 76396
rect 168668 76332 168669 76396
rect 168603 76331 168669 76332
rect 169339 76396 169405 76397
rect 169339 76332 169340 76396
rect 169404 76332 169405 76396
rect 169339 76331 169405 76332
rect 168294 61954 168914 76000
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 169342 26893 169402 76331
rect 170078 75717 170138 77827
rect 170075 75716 170141 75717
rect 170075 75652 170076 75716
rect 170140 75652 170141 75716
rect 170075 75651 170141 75652
rect 170262 75037 170322 77827
rect 170259 75036 170325 75037
rect 170259 74972 170260 75036
rect 170324 74972 170325 75036
rect 170259 74971 170325 74972
rect 169339 26892 169405 26893
rect 169339 26828 169340 26892
rect 169404 26828 169405 26892
rect 169339 26827 169405 26828
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168051 4860 168117 4861
rect 168051 4796 168052 4860
rect 168116 4796 168117 4860
rect 168051 4795 168117 4796
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 -5146 168914 25398
rect 170630 11661 170690 77827
rect 170811 77756 170877 77757
rect 170811 77692 170812 77756
rect 170876 77692 170877 77756
rect 170811 77691 170877 77692
rect 170814 24173 170874 77691
rect 170998 77213 171058 77827
rect 170995 77212 171061 77213
rect 170995 77148 170996 77212
rect 171060 77148 171061 77212
rect 170995 77147 171061 77148
rect 171366 76397 171426 78371
rect 171550 77349 171610 78371
rect 171915 77892 171981 77893
rect 171915 77828 171916 77892
rect 171980 77890 171981 77892
rect 172467 77892 172533 77893
rect 171980 77830 172162 77890
rect 171980 77828 171981 77830
rect 171915 77827 171981 77828
rect 172102 77485 172162 77830
rect 172467 77828 172468 77892
rect 172532 77828 172533 77892
rect 172467 77827 172533 77828
rect 173019 77892 173085 77893
rect 173019 77828 173020 77892
rect 173084 77828 173085 77892
rect 173019 77827 173085 77828
rect 172099 77484 172165 77485
rect 172099 77420 172100 77484
rect 172164 77420 172165 77484
rect 172099 77419 172165 77420
rect 171547 77348 171613 77349
rect 171547 77284 171548 77348
rect 171612 77284 171613 77348
rect 171547 77283 171613 77284
rect 171363 76396 171429 76397
rect 171363 76332 171364 76396
rect 171428 76332 171429 76396
rect 171363 76331 171429 76332
rect 172470 76125 172530 77827
rect 173022 76261 173082 77827
rect 173574 77621 173634 78507
rect 173571 77620 173637 77621
rect 173571 77556 173572 77620
rect 173636 77556 173637 77620
rect 173571 77555 173637 77556
rect 173019 76260 173085 76261
rect 173019 76196 173020 76260
rect 173084 76196 173085 76260
rect 173019 76195 173085 76196
rect 172467 76124 172533 76125
rect 172467 76060 172468 76124
rect 172532 76060 172533 76124
rect 172467 76059 172533 76060
rect 170995 75716 171061 75717
rect 170995 75652 170996 75716
rect 171060 75652 171061 75716
rect 170995 75651 171061 75652
rect 170998 71093 171058 75651
rect 171731 74764 171797 74765
rect 171731 74700 171732 74764
rect 171796 74700 171797 74764
rect 171731 74699 171797 74700
rect 170995 71092 171061 71093
rect 170995 71028 170996 71092
rect 171060 71028 171061 71092
rect 170995 71027 171061 71028
rect 170811 24172 170877 24173
rect 170811 24108 170812 24172
rect 170876 24108 170877 24172
rect 170811 24107 170877 24108
rect 170627 11660 170693 11661
rect 170627 11596 170628 11660
rect 170692 11596 170693 11660
rect 170627 11595 170693 11596
rect 171734 3365 171794 74699
rect 171915 73268 171981 73269
rect 171915 73204 171916 73268
rect 171980 73204 171981 73268
rect 171915 73203 171981 73204
rect 171918 50285 171978 73203
rect 172794 66454 173414 76000
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 171915 50284 171981 50285
rect 171915 50220 171916 50284
rect 171980 50220 171981 50284
rect 171915 50219 171981 50220
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 171731 3364 171797 3365
rect 171731 3300 171732 3364
rect 171796 3300 171797 3364
rect 171731 3299 171797 3300
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 70954 177914 76000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 75454 182414 76000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 228453 191414 228484
rect 190794 228217 190826 228453
rect 191062 228217 191146 228453
rect 191382 228217 191414 228453
rect 190794 228133 191414 228217
rect 190794 227897 190826 228133
rect 191062 227897 191146 228133
rect 191382 227897 191414 228133
rect 190794 192454 191414 227897
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 196954 195914 228484
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 201454 200414 228484
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 205954 204914 228484
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 210454 209414 228484
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 214954 213914 228484
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 219454 218414 228484
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 223954 222914 228484
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 228453 227414 228484
rect 226794 228217 226826 228453
rect 227062 228217 227146 228453
rect 227382 228217 227414 228453
rect 226794 228133 227414 228217
rect 226794 227897 226826 228133
rect 227062 227897 227146 228133
rect 227382 227897 227414 228133
rect 226794 192454 227414 227897
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 196954 231914 228484
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 201454 236414 228484
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 205954 240914 228484
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 210454 245414 228484
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 214954 249914 228484
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 219454 254414 228484
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 223954 258914 228484
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 228453 263414 228484
rect 262794 228217 262826 228453
rect 263062 228217 263146 228453
rect 263382 228217 263414 228453
rect 262794 228133 263414 228217
rect 262794 227897 262826 228133
rect 263062 227897 263146 228133
rect 263382 227897 263414 228133
rect 262794 192454 263414 227897
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 196954 267914 228484
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 201454 272414 228484
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 205954 276914 228484
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 210454 281414 228484
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 214954 285914 228484
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 219454 290414 228484
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 223954 294914 228484
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 228453 299414 228484
rect 298794 228217 298826 228453
rect 299062 228217 299146 228453
rect 299382 228217 299414 228453
rect 298794 228133 299414 228217
rect 298794 227897 298826 228133
rect 299062 227897 299146 228133
rect 299382 227897 299414 228133
rect 298794 192454 299414 227897
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 196954 303914 228484
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 201454 308414 228484
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 205954 312914 228484
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 210454 317414 228484
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 214954 321914 228484
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 219454 326414 228484
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 223954 330914 228484
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 228453 335414 228484
rect 334794 228217 334826 228453
rect 335062 228217 335146 228453
rect 335382 228217 335414 228453
rect 334794 228133 335414 228217
rect 334794 227897 334826 228133
rect 335062 227897 335146 228133
rect 335382 227897 335414 228133
rect 334794 192454 335414 227897
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 196954 339914 228484
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 201454 344414 228484
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 205954 348914 228484
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 210454 353414 228484
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 214954 357914 228484
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 219454 362414 228484
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 223954 366914 228484
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 228453 371414 228484
rect 370794 228217 370826 228453
rect 371062 228217 371146 228453
rect 371382 228217 371414 228453
rect 370794 228133 371414 228217
rect 370794 227897 370826 228133
rect 371062 227897 371146 228133
rect 371382 227897 371414 228133
rect 370794 192454 371414 227897
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 196954 375914 228484
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 201454 380414 228484
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 205954 384914 228484
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 210454 389414 228484
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 214954 393914 228484
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 396582 77757 396642 643179
rect 396766 227765 396826 643723
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 248684 398414 254898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 396763 227764 396829 227765
rect 396763 227700 396764 227764
rect 396828 227700 396829 227764
rect 396763 227699 396829 227700
rect 397794 219454 398414 228484
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 396579 77756 396645 77757
rect 396579 77692 396580 77756
rect 396644 77692 396645 77756
rect 396579 77691 396645 77692
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 65342 246067 65578 246303
rect 65662 246067 65898 246303
rect 65982 246067 66218 246303
rect 66302 246067 66538 246303
rect 66622 246067 66858 246303
rect 66942 246067 67178 246303
rect 67262 246067 67498 246303
rect 67582 246067 67818 246303
rect 67902 246067 68138 246303
rect 68222 246067 68458 246303
rect 68542 246067 68778 246303
rect 68862 246067 69098 246303
rect 69182 246067 69418 246303
rect 69502 246067 69738 246303
rect 69822 246067 70058 246303
rect 65462 241717 65698 241953
rect 65782 241717 66018 241953
rect 66102 241717 66338 241953
rect 66422 241717 66658 241953
rect 66742 241717 66978 241953
rect 67062 241717 67298 241953
rect 67382 241717 67618 241953
rect 67702 241717 67938 241953
rect 68022 241717 68258 241953
rect 68342 241717 68578 241953
rect 68662 241717 68898 241953
rect 68982 241717 69218 241953
rect 69302 241717 69538 241953
rect 69622 241717 69858 241953
rect 69942 241717 70178 241953
rect 70262 241717 70498 241953
rect 70582 241717 70818 241953
rect 70902 241717 71138 241953
rect 65462 241397 65698 241633
rect 65782 241397 66018 241633
rect 66102 241397 66338 241633
rect 66422 241397 66658 241633
rect 66742 241397 66978 241633
rect 67062 241397 67298 241633
rect 67382 241397 67618 241633
rect 67702 241397 67938 241633
rect 68022 241397 68258 241633
rect 68342 241397 68578 241633
rect 68662 241397 68898 241633
rect 68982 241397 69218 241633
rect 69302 241397 69538 241633
rect 69622 241397 69858 241633
rect 69942 241397 70178 241633
rect 70262 241397 70498 241633
rect 70582 241397 70818 241633
rect 70902 241397 71138 241633
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 228217 47062 228453
rect 47146 228217 47382 228453
rect 46826 227897 47062 228133
rect 47146 227897 47382 228133
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 228217 83062 228453
rect 83146 228217 83382 228453
rect 82826 227897 83062 228133
rect 83146 227897 83382 228133
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 118826 228217 119062 228453
rect 119146 228217 119382 228453
rect 118826 227897 119062 228133
rect 119146 227897 119382 228133
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 136036 205625 136272 205861
rect 136356 205625 136592 205861
rect 136676 205625 136912 205861
rect 136996 205625 137232 205861
rect 137316 205625 137552 205861
rect 137636 205625 137872 205861
rect 137956 205625 138192 205861
rect 138276 205625 138512 205861
rect 138596 205625 138832 205861
rect 138916 205625 139152 205861
rect 139236 205625 139472 205861
rect 139556 205625 139792 205861
rect 139876 205625 140112 205861
rect 140196 205625 140432 205861
rect 140516 205625 140752 205861
rect 140836 205625 141072 205861
rect 141156 205625 141392 205861
rect 141476 205625 141712 205861
rect 141796 205625 142032 205861
rect 142116 205625 142352 205861
rect 142436 205625 142672 205861
rect 142756 205625 142992 205861
rect 143076 205625 143312 205861
rect 143396 205625 143632 205861
rect 143716 205625 143952 205861
rect 144036 205625 144272 205861
rect 144356 205625 144592 205861
rect 144676 205625 144912 205861
rect 144996 205625 145232 205861
rect 145316 205625 145552 205861
rect 145636 205625 145872 205861
rect 145956 205625 146192 205861
rect 146276 205625 146512 205861
rect 146596 205625 146832 205861
rect 146916 205625 147152 205861
rect 147236 205625 147472 205861
rect 147556 205625 147792 205861
rect 147876 205625 148112 205861
rect 148196 205625 148432 205861
rect 148516 205625 148752 205861
rect 148836 205625 149072 205861
rect 149156 205625 149392 205861
rect 149476 205625 149712 205861
rect 149796 205625 150032 205861
rect 150116 205625 150352 205861
rect 150436 205625 150672 205861
rect 150756 205625 150992 205861
rect 151076 205625 151312 205861
rect 151396 205625 151632 205861
rect 151716 205625 151952 205861
rect 152036 205625 152272 205861
rect 152356 205625 152592 205861
rect 152676 205625 152912 205861
rect 152996 205625 153232 205861
rect 153316 205625 153552 205861
rect 153636 205625 153872 205861
rect 153956 205625 154192 205861
rect 154276 205625 154512 205861
rect 154596 205625 154832 205861
rect 154916 205625 155152 205861
rect 155236 205625 155472 205861
rect 155556 205625 155792 205861
rect 155876 205625 156112 205861
rect 156196 205625 156432 205861
rect 156516 205625 156752 205861
rect 156836 205625 157072 205861
rect 157156 205625 157392 205861
rect 157476 205625 157712 205861
rect 157796 205625 158032 205861
rect 158116 205625 158352 205861
rect 158436 205625 158672 205861
rect 158756 205625 158992 205861
rect 159076 205625 159312 205861
rect 159396 205625 159632 205861
rect 159716 205625 159952 205861
rect 160036 205625 160272 205861
rect 160356 205625 160592 205861
rect 160676 205625 160912 205861
rect 160996 205625 161232 205861
rect 161316 205625 161552 205861
rect 161636 205625 161872 205861
rect 161956 205625 162192 205861
rect 162276 205625 162512 205861
rect 162596 205625 162832 205861
rect 162916 205625 163152 205861
rect 163236 205625 163472 205861
rect 163556 205625 163792 205861
rect 163876 205625 164112 205861
rect 164196 205625 164432 205861
rect 164516 205625 164752 205861
rect 164836 205625 165072 205861
rect 165156 205625 165392 205861
rect 137376 201175 137612 201411
rect 137696 201175 137932 201411
rect 138016 201175 138252 201411
rect 138336 201175 138572 201411
rect 138656 201175 138892 201411
rect 138976 201175 139212 201411
rect 139296 201175 139532 201411
rect 139616 201175 139852 201411
rect 139936 201175 140172 201411
rect 140256 201175 140492 201411
rect 140576 201175 140812 201411
rect 140896 201175 141132 201411
rect 141216 201175 141452 201411
rect 141536 201175 141772 201411
rect 141856 201175 142092 201411
rect 142176 201175 142412 201411
rect 142496 201175 142732 201411
rect 142816 201175 143052 201411
rect 143136 201175 143372 201411
rect 143456 201175 143692 201411
rect 143776 201175 144012 201411
rect 144096 201175 144332 201411
rect 144416 201175 144652 201411
rect 144736 201175 144972 201411
rect 145056 201175 145292 201411
rect 145376 201175 145612 201411
rect 145696 201175 145932 201411
rect 146016 201175 146252 201411
rect 146336 201175 146572 201411
rect 146656 201175 146892 201411
rect 146976 201175 147212 201411
rect 147296 201175 147532 201411
rect 147616 201175 147852 201411
rect 147936 201175 148172 201411
rect 148256 201175 148492 201411
rect 148576 201175 148812 201411
rect 148896 201175 149132 201411
rect 149216 201175 149452 201411
rect 149536 201175 149772 201411
rect 149856 201175 150092 201411
rect 150176 201175 150412 201411
rect 150496 201175 150732 201411
rect 150816 201175 151052 201411
rect 151136 201175 151372 201411
rect 151456 201175 151692 201411
rect 151776 201175 152012 201411
rect 152096 201175 152332 201411
rect 152416 201175 152652 201411
rect 152736 201175 152972 201411
rect 153056 201175 153292 201411
rect 153376 201175 153612 201411
rect 153696 201175 153932 201411
rect 154016 201175 154252 201411
rect 154336 201175 154572 201411
rect 154656 201175 154892 201411
rect 154976 201175 155212 201411
rect 155296 201175 155532 201411
rect 155616 201175 155852 201411
rect 155936 201175 156172 201411
rect 156256 201175 156492 201411
rect 156576 201175 156812 201411
rect 156896 201175 157132 201411
rect 157216 201175 157452 201411
rect 157536 201175 157772 201411
rect 157856 201175 158092 201411
rect 158176 201175 158412 201411
rect 158496 201175 158732 201411
rect 158816 201175 159052 201411
rect 159136 201175 159372 201411
rect 159456 201175 159692 201411
rect 159776 201175 160012 201411
rect 160096 201175 160332 201411
rect 160416 201175 160652 201411
rect 160736 201175 160972 201411
rect 161056 201175 161292 201411
rect 161376 201175 161612 201411
rect 161696 201175 161932 201411
rect 162016 201175 162252 201411
rect 162336 201175 162572 201411
rect 162656 201175 162892 201411
rect 162976 201175 163212 201411
rect 163296 201175 163532 201411
rect 163616 201175 163852 201411
rect 163936 201175 164172 201411
rect 164256 201175 164492 201411
rect 164576 201175 164812 201411
rect 164896 201175 165132 201411
rect 165216 201175 165452 201411
rect 137066 174218 137302 174454
rect 137386 174218 137622 174454
rect 137706 174218 137942 174454
rect 138026 174218 138262 174454
rect 138346 174218 138582 174454
rect 138666 174218 138902 174454
rect 138986 174218 139222 174454
rect 139306 174218 139542 174454
rect 139626 174218 139862 174454
rect 139946 174218 140182 174454
rect 140266 174218 140502 174454
rect 140586 174218 140822 174454
rect 140906 174218 141142 174454
rect 141226 174218 141462 174454
rect 137066 173898 137302 174134
rect 137386 173898 137622 174134
rect 137706 173898 137942 174134
rect 138026 173898 138262 174134
rect 138346 173898 138582 174134
rect 138666 173898 138902 174134
rect 138986 173898 139222 174134
rect 139306 173898 139542 174134
rect 139626 173898 139862 174134
rect 139946 173898 140182 174134
rect 140266 173898 140502 174134
rect 140586 173898 140822 174134
rect 140906 173898 141142 174134
rect 141226 173898 141462 174134
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 139610 115718 139846 115954
rect 139610 115398 139846 115634
rect 170330 115718 170566 115954
rect 170330 115398 170566 115634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 228217 191062 228453
rect 191146 228217 191382 228453
rect 190826 227897 191062 228133
rect 191146 227897 191382 228133
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 228217 227062 228453
rect 227146 228217 227382 228453
rect 226826 227897 227062 228133
rect 227146 227897 227382 228133
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 228217 263062 228453
rect 263146 228217 263382 228453
rect 262826 227897 263062 228133
rect 263146 227897 263382 228133
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 228217 299062 228453
rect 299146 228217 299382 228453
rect 298826 227897 299062 228133
rect 299146 227897 299382 228133
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 228217 335062 228453
rect 335146 228217 335382 228453
rect 334826 227897 335062 228133
rect 335146 227897 335382 228133
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 228217 371062 228453
rect 371146 228217 371382 228453
rect 370826 227897 371062 228133
rect 371146 227897 371382 228133
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246303 424826 246454
rect 29382 246218 65342 246303
rect -8726 246134 65342 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 246067 65342 246134
rect 65578 246067 65662 246303
rect 65898 246067 65982 246303
rect 66218 246067 66302 246303
rect 66538 246067 66622 246303
rect 66858 246067 66942 246303
rect 67178 246067 67262 246303
rect 67498 246067 67582 246303
rect 67818 246067 67902 246303
rect 68138 246067 68222 246303
rect 68458 246067 68542 246303
rect 68778 246067 68862 246303
rect 69098 246067 69182 246303
rect 69418 246067 69502 246303
rect 69738 246067 69822 246303
rect 70058 246218 424826 246303
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect 70058 246134 592650 246218
rect 70058 246067 424826 246134
rect 29382 245898 424826 246067
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241953 420326 241954
rect 24882 241718 65462 241953
rect -8726 241717 65462 241718
rect 65698 241717 65782 241953
rect 66018 241717 66102 241953
rect 66338 241717 66422 241953
rect 66658 241717 66742 241953
rect 66978 241717 67062 241953
rect 67298 241717 67382 241953
rect 67618 241717 67702 241953
rect 67938 241717 68022 241953
rect 68258 241717 68342 241953
rect 68578 241717 68662 241953
rect 68898 241717 68982 241953
rect 69218 241717 69302 241953
rect 69538 241717 69622 241953
rect 69858 241717 69942 241953
rect 70178 241717 70262 241953
rect 70498 241717 70582 241953
rect 70818 241717 70902 241953
rect 71138 241718 420326 241953
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect 71138 241717 592650 241718
rect -8726 241634 592650 241717
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241633 420326 241634
rect 24882 241398 65462 241633
rect -8726 241397 65462 241398
rect 65698 241397 65782 241633
rect 66018 241397 66102 241633
rect 66338 241397 66422 241633
rect 66658 241397 66742 241633
rect 66978 241397 67062 241633
rect 67298 241397 67382 241633
rect 67618 241397 67702 241633
rect 67938 241397 68022 241633
rect 68258 241397 68342 241633
rect 68578 241397 68662 241633
rect 68898 241397 68982 241633
rect 69218 241397 69302 241633
rect 69538 241397 69622 241633
rect 69858 241397 69942 241633
rect 70178 241397 70262 241633
rect 70498 241397 70582 241633
rect 70818 241397 70902 241633
rect 71138 241398 420326 241633
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect 71138 241397 592650 241398
rect -8726 241366 592650 241397
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228453 406826 228454
rect 11382 228218 46826 228453
rect -8726 228217 46826 228218
rect 47062 228217 47146 228453
rect 47382 228217 82826 228453
rect 83062 228217 83146 228453
rect 83382 228217 118826 228453
rect 119062 228217 119146 228453
rect 119382 228217 190826 228453
rect 191062 228217 191146 228453
rect 191382 228217 226826 228453
rect 227062 228217 227146 228453
rect 227382 228217 262826 228453
rect 263062 228217 263146 228453
rect 263382 228217 298826 228453
rect 299062 228217 299146 228453
rect 299382 228217 334826 228453
rect 335062 228217 335146 228453
rect 335382 228217 370826 228453
rect 371062 228217 371146 228453
rect 371382 228218 406826 228453
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect 371382 228217 592650 228218
rect -8726 228134 592650 228217
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 228133 406826 228134
rect 11382 227898 46826 228133
rect -8726 227897 46826 227898
rect 47062 227897 47146 228133
rect 47382 227897 82826 228133
rect 83062 227897 83146 228133
rect 83382 227897 118826 228133
rect 119062 227897 119146 228133
rect 119382 227897 190826 228133
rect 191062 227897 191146 228133
rect 191382 227897 226826 228133
rect 227062 227897 227146 228133
rect 227382 227897 262826 228133
rect 263062 227897 263146 228133
rect 263382 227897 298826 228133
rect 299062 227897 299146 228133
rect 299382 227897 334826 228133
rect 335062 227897 335146 228133
rect 335382 227897 370826 228133
rect 371062 227897 371146 228133
rect 371382 227898 406826 228133
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect 371382 227897 592650 227898
rect -8726 227866 592650 227897
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205861 204326 205954
rect 132882 205718 136036 205861
rect -8726 205634 136036 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205625 136036 205634
rect 136272 205625 136356 205861
rect 136592 205625 136676 205861
rect 136912 205625 136996 205861
rect 137232 205625 137316 205861
rect 137552 205625 137636 205861
rect 137872 205625 137956 205861
rect 138192 205625 138276 205861
rect 138512 205625 138596 205861
rect 138832 205625 138916 205861
rect 139152 205625 139236 205861
rect 139472 205625 139556 205861
rect 139792 205625 139876 205861
rect 140112 205625 140196 205861
rect 140432 205625 140516 205861
rect 140752 205625 140836 205861
rect 141072 205625 141156 205861
rect 141392 205625 141476 205861
rect 141712 205625 141796 205861
rect 142032 205625 142116 205861
rect 142352 205625 142436 205861
rect 142672 205625 142756 205861
rect 142992 205625 143076 205861
rect 143312 205625 143396 205861
rect 143632 205625 143716 205861
rect 143952 205625 144036 205861
rect 144272 205625 144356 205861
rect 144592 205625 144676 205861
rect 144912 205625 144996 205861
rect 145232 205625 145316 205861
rect 145552 205625 145636 205861
rect 145872 205625 145956 205861
rect 146192 205625 146276 205861
rect 146512 205625 146596 205861
rect 146832 205625 146916 205861
rect 147152 205625 147236 205861
rect 147472 205625 147556 205861
rect 147792 205625 147876 205861
rect 148112 205625 148196 205861
rect 148432 205625 148516 205861
rect 148752 205625 148836 205861
rect 149072 205625 149156 205861
rect 149392 205625 149476 205861
rect 149712 205625 149796 205861
rect 150032 205625 150116 205861
rect 150352 205625 150436 205861
rect 150672 205625 150756 205861
rect 150992 205625 151076 205861
rect 151312 205625 151396 205861
rect 151632 205625 151716 205861
rect 151952 205625 152036 205861
rect 152272 205625 152356 205861
rect 152592 205625 152676 205861
rect 152912 205625 152996 205861
rect 153232 205625 153316 205861
rect 153552 205625 153636 205861
rect 153872 205625 153956 205861
rect 154192 205625 154276 205861
rect 154512 205625 154596 205861
rect 154832 205625 154916 205861
rect 155152 205625 155236 205861
rect 155472 205625 155556 205861
rect 155792 205625 155876 205861
rect 156112 205625 156196 205861
rect 156432 205625 156516 205861
rect 156752 205625 156836 205861
rect 157072 205625 157156 205861
rect 157392 205625 157476 205861
rect 157712 205625 157796 205861
rect 158032 205625 158116 205861
rect 158352 205625 158436 205861
rect 158672 205625 158756 205861
rect 158992 205625 159076 205861
rect 159312 205625 159396 205861
rect 159632 205625 159716 205861
rect 159952 205625 160036 205861
rect 160272 205625 160356 205861
rect 160592 205625 160676 205861
rect 160912 205625 160996 205861
rect 161232 205625 161316 205861
rect 161552 205625 161636 205861
rect 161872 205625 161956 205861
rect 162192 205625 162276 205861
rect 162512 205625 162596 205861
rect 162832 205625 162916 205861
rect 163152 205625 163236 205861
rect 163472 205625 163556 205861
rect 163792 205625 163876 205861
rect 164112 205625 164196 205861
rect 164432 205625 164516 205861
rect 164752 205625 164836 205861
rect 165072 205625 165156 205861
rect 165392 205718 204326 205861
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect 165392 205634 592650 205718
rect 165392 205625 204326 205634
rect 132882 205398 204326 205625
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201411 199826 201454
rect 128382 201218 137376 201411
rect -8726 201175 137376 201218
rect 137612 201175 137696 201411
rect 137932 201175 138016 201411
rect 138252 201175 138336 201411
rect 138572 201175 138656 201411
rect 138892 201175 138976 201411
rect 139212 201175 139296 201411
rect 139532 201175 139616 201411
rect 139852 201175 139936 201411
rect 140172 201175 140256 201411
rect 140492 201175 140576 201411
rect 140812 201175 140896 201411
rect 141132 201175 141216 201411
rect 141452 201175 141536 201411
rect 141772 201175 141856 201411
rect 142092 201175 142176 201411
rect 142412 201175 142496 201411
rect 142732 201175 142816 201411
rect 143052 201175 143136 201411
rect 143372 201175 143456 201411
rect 143692 201175 143776 201411
rect 144012 201175 144096 201411
rect 144332 201175 144416 201411
rect 144652 201175 144736 201411
rect 144972 201175 145056 201411
rect 145292 201175 145376 201411
rect 145612 201175 145696 201411
rect 145932 201175 146016 201411
rect 146252 201175 146336 201411
rect 146572 201175 146656 201411
rect 146892 201175 146976 201411
rect 147212 201175 147296 201411
rect 147532 201175 147616 201411
rect 147852 201175 147936 201411
rect 148172 201175 148256 201411
rect 148492 201175 148576 201411
rect 148812 201175 148896 201411
rect 149132 201175 149216 201411
rect 149452 201175 149536 201411
rect 149772 201175 149856 201411
rect 150092 201175 150176 201411
rect 150412 201175 150496 201411
rect 150732 201175 150816 201411
rect 151052 201175 151136 201411
rect 151372 201175 151456 201411
rect 151692 201175 151776 201411
rect 152012 201175 152096 201411
rect 152332 201175 152416 201411
rect 152652 201175 152736 201411
rect 152972 201175 153056 201411
rect 153292 201175 153376 201411
rect 153612 201175 153696 201411
rect 153932 201175 154016 201411
rect 154252 201175 154336 201411
rect 154572 201175 154656 201411
rect 154892 201175 154976 201411
rect 155212 201175 155296 201411
rect 155532 201175 155616 201411
rect 155852 201175 155936 201411
rect 156172 201175 156256 201411
rect 156492 201175 156576 201411
rect 156812 201175 156896 201411
rect 157132 201175 157216 201411
rect 157452 201175 157536 201411
rect 157772 201175 157856 201411
rect 158092 201175 158176 201411
rect 158412 201175 158496 201411
rect 158732 201175 158816 201411
rect 159052 201175 159136 201411
rect 159372 201175 159456 201411
rect 159692 201175 159776 201411
rect 160012 201175 160096 201411
rect 160332 201175 160416 201411
rect 160652 201175 160736 201411
rect 160972 201175 161056 201411
rect 161292 201175 161376 201411
rect 161612 201175 161696 201411
rect 161932 201175 162016 201411
rect 162252 201175 162336 201411
rect 162572 201175 162656 201411
rect 162892 201175 162976 201411
rect 163212 201175 163296 201411
rect 163532 201175 163616 201411
rect 163852 201175 163936 201411
rect 164172 201175 164256 201411
rect 164492 201175 164576 201411
rect 164812 201175 164896 201411
rect 165132 201175 165216 201411
rect 165452 201218 199826 201411
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect 165452 201175 592650 201218
rect -8726 201134 592650 201175
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 137066 174454
rect 137302 174218 137386 174454
rect 137622 174218 137706 174454
rect 137942 174218 138026 174454
rect 138262 174218 138346 174454
rect 138582 174218 138666 174454
rect 138902 174218 138986 174454
rect 139222 174218 139306 174454
rect 139542 174218 139626 174454
rect 139862 174218 139946 174454
rect 140182 174218 140266 174454
rect 140502 174218 140586 174454
rect 140822 174218 140906 174454
rect 141142 174218 141226 174454
rect 141462 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 137066 174134
rect 137302 173898 137386 174134
rect 137622 173898 137706 174134
rect 137942 173898 138026 174134
rect 138262 173898 138346 174134
rect 138582 173898 138666 174134
rect 138902 173898 138986 174134
rect 139222 173898 139306 174134
rect 139542 173898 139626 174134
rect 139862 173898 139946 174134
rect 140182 173898 140266 174134
rect 140502 173898 140586 174134
rect 140822 173898 140906 174134
rect 141142 173898 141226 174134
rect 141462 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 139610 115954
rect 139846 115718 170330 115954
rect 170566 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 139610 115634
rect 139846 115398 170330 115634
rect 170566 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 154970 111454
rect 155206 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 154970 111134
rect 155206 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use PD_M1_M2  PD_M1_M2_macro0
timestamp 0
transform 1 0 16000 0 1 232484
box 30000 -2000 380500 14200
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 120000 0 1 78000
box 0 0 60000 60000
use SystemLevel  sl_macro0
timestamp 0
transform 1 0 148914 0 1 188300
box -13000 -15200 17500 18000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 248684 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 248684 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 248684 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 76000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 140000 182414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 248684 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 248684 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 248684 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 248684 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 248684 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 248684 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 228484 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 248684 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 248684 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 248684 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 140000 119414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 248684 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 76000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 248684 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 248684 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 248684 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 248684 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 248684 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 248684 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 228484 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 248684 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 248684 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 248684 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 140000 128414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 248684 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 76000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 248684 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 248684 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 248684 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 248684 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 248684 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 248684 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 228484 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 248684 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 248684 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 248684 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 248684 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 76000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 140000 173414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 248684 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 248684 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 248684 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 248684 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 248684 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 248684 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 228484 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 248684 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 248684 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 248684 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 140000 132914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 248684 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 76000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 248684 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 248684 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 248684 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 248684 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 248684 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 248684 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 228484 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 248684 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 248684 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 248684 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 248684 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 76000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 140000 177914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 248684 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 248684 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 248684 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 248684 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 248684 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 248684 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 228484 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 248684 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 248684 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 248684 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 76000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 248684 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 248684 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 248684 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 248684 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 248684 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 248684 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 228484 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 248684 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 248684 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 248684 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 140000 123914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 248684 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 76000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 248684 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 248684 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 248684 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 248684 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 248684 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 248684 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 228484 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 248684 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
